module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    compressor_CLA256_16 compressor_CLA256_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
        src12 <= 256'h0;
        src13 <= 256'h0;
        src14 <= 256'h0;
        src15 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA256_16(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    input [255:0]src12,
    input [255:0]src13,
    input [255:0]src14,
    input [255:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [0:0] comp_out23;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      input wire [255:0] src12,
      input wire [255:0] src13,
      input wire [255:0] src14,
      input wire [255:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [0:0] dst23);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [255:0] stage0_12;
   wire [255:0] stage0_13;
   wire [255:0] stage0_14;
   wire [255:0] stage0_15;
   wire [48:0] stage1_0;
   wire [97:0] stage1_1;
   wire [97:0] stage1_2;
   wire [113:0] stage1_3;
   wire [126:0] stage1_4;
   wire [104:0] stage1_5;
   wire [103:0] stage1_6;
   wire [114:0] stage1_7;
   wire [105:0] stage1_8;
   wire [115:0] stage1_9;
   wire [113:0] stage1_10;
   wire [114:0] stage1_11;
   wire [101:0] stage1_12;
   wire [132:0] stage1_13;
   wire [156:0] stage1_14;
   wire [75:0] stage1_15;
   wire [67:0] stage1_16;
   wire [41:0] stage1_17;
   wire [8:0] stage2_0;
   wire [25:0] stage2_1;
   wire [45:0] stage2_2;
   wire [33:0] stage2_3;
   wire [49:0] stage2_4;
   wire [54:0] stage2_5;
   wire [39:0] stage2_6;
   wire [58:0] stage2_7;
   wire [49:0] stage2_8;
   wire [47:0] stage2_9;
   wire [35:0] stage2_10;
   wire [47:0] stage2_11;
   wire [60:0] stage2_12;
   wire [44:0] stage2_13;
   wire [50:0] stage2_14;
   wire [50:0] stage2_15;
   wire [47:0] stage2_16;
   wire [33:0] stage2_17;
   wire [13:0] stage2_18;
   wire [4:0] stage2_19;
   wire [6:0] stage3_0;
   wire [5:0] stage3_1;
   wire [13:0] stage3_2;
   wire [13:0] stage3_3;
   wire [13:0] stage3_4;
   wire [19:0] stage3_5;
   wire [24:0] stage3_6;
   wire [22:0] stage3_7;
   wire [16:0] stage3_8;
   wire [20:0] stage3_9;
   wire [22:0] stage3_10;
   wire [16:0] stage3_11;
   wire [22:0] stage3_12;
   wire [20:0] stage3_13;
   wire [21:0] stage3_14;
   wire [24:0] stage3_15;
   wire [24:0] stage3_16;
   wire [18:0] stage3_17;
   wire [13:0] stage3_18;
   wire [11:0] stage3_19;
   wire [1:0] stage3_20;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [9:0] stage4_2;
   wire [5:0] stage4_3;
   wire [5:0] stage4_4;
   wire [5:0] stage4_5;
   wire [7:0] stage4_6;
   wire [16:0] stage4_7;
   wire [7:0] stage4_8;
   wire [8:0] stage4_9;
   wire [9:0] stage4_10;
   wire [9:0] stage4_11;
   wire [6:0] stage4_12;
   wire [7:0] stage4_13;
   wire [10:0] stage4_14;
   wire [8:0] stage4_15;
   wire [8:0] stage4_16;
   wire [9:0] stage4_17;
   wire [8:0] stage4_18;
   wire [9:0] stage4_19;
   wire [3:0] stage4_20;
   wire [1:0] stage4_21;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [5:0] stage5_2;
   wire [1:0] stage5_3;
   wire [6:0] stage5_4;
   wire [0:0] stage5_5;
   wire [4:0] stage5_6;
   wire [3:0] stage5_7;
   wire [3:0] stage5_8;
   wire [3:0] stage5_9;
   wire [5:0] stage5_10;
   wire [4:0] stage5_11;
   wire [2:0] stage5_12;
   wire [3:0] stage5_13;
   wire [3:0] stage5_14;
   wire [5:0] stage5_15;
   wire [4:0] stage5_16;
   wire [2:0] stage5_17;
   wire [3:0] stage5_18;
   wire [5:0] stage5_19;
   wire [5:0] stage5_20;
   wire [1:0] stage5_21;
   wire [0:0] stage5_22;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;
   wire [0:0] stage6_23;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[30], stage0_1[31], stage0_1[32]},
      {stage0_2[10]},
      {stage0_3[20], stage0_3[21]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc2135_5 gpc11 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[11]},
      {stage0_3[22], stage0_3[23]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc2135_5 gpc12 (
      {stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[36], stage0_1[37], stage0_1[38]},
      {stage0_2[12]},
      {stage0_3[24], stage0_3[25]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc2135_5 gpc13 (
      {stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[13]},
      {stage0_3[26], stage0_3[27]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc2135_5 gpc14 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_1[42], stage0_1[43], stage0_1[44]},
      {stage0_2[14]},
      {stage0_3[28], stage0_3[29]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc2135_5 gpc15 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[15]},
      {stage0_3[30], stage0_3[31]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc2135_5 gpc16 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_1[48], stage0_1[49], stage0_1[50]},
      {stage0_2[16]},
      {stage0_3[32], stage0_3[33]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc117_4 gpc17 (
      {stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_1[51]},
      {stage0_2[17]},
      {stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc117_4 gpc18 (
      {stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_1[52]},
      {stage0_2[18]},
      {stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc117_4 gpc19 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[53]},
      {stage0_2[19]},
      {stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[20]},
      {stage0_3[34]},
      {stage1_4[17],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[21]},
      {stage0_3[35]},
      {stage1_4[18],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[22]},
      {stage0_3[36]},
      {stage1_4[19],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[23]},
      {stage0_3[37]},
      {stage1_4[20],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[24]},
      {stage0_3[38]},
      {stage1_4[21],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[25]},
      {stage0_3[39]},
      {stage1_4[22],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[26]},
      {stage0_3[40]},
      {stage1_4[23],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[27]},
      {stage0_3[41]},
      {stage1_4[24],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33]},
      {stage1_4[25],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39]},
      {stage1_4[26],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45]},
      {stage1_4[27],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51]},
      {stage1_4[28],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57]},
      {stage1_4[29],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163], stage0_0[164], stage0_0[165]},
      {stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63]},
      {stage1_4[30],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169], stage0_0[170], stage0_0[171]},
      {stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69]},
      {stage1_4[31],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175], stage0_0[176], stage0_0[177]},
      {stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75]},
      {stage1_4[32],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181], stage0_0[182], stage0_0[183]},
      {stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81]},
      {stage1_4[33],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187], stage0_0[188], stage0_0[189]},
      {stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87]},
      {stage1_4[34],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195]},
      {stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93]},
      {stage1_4[35],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201]},
      {stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99]},
      {stage1_4[36],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207]},
      {stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105]},
      {stage1_4[37],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213]},
      {stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111]},
      {stage1_4[38],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[214], stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219]},
      {stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117]},
      {stage1_4[39],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[220], stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225]},
      {stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123]},
      {stage1_4[40],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[226], stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231]},
      {stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129]},
      {stage1_4[41],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[232], stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237]},
      {stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135]},
      {stage1_4[42],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[238], stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243]},
      {stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141]},
      {stage1_4[43],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[244], stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249]},
      {stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147]},
      {stage1_4[44],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[250], stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255]},
      {stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153]},
      {stage1_4[45],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage1_5[0],stage1_4[46],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53]},
      {stage1_5[1],stage1_4[47],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59]},
      {stage1_5[2],stage1_4[48],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65]},
      {stage1_5[3],stage1_4[49],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71]},
      {stage1_5[4],stage1_4[50],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77]},
      {stage1_5[5],stage1_4[51],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83]},
      {stage1_5[6],stage1_4[52],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89]},
      {stage1_5[7],stage1_4[53],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95]},
      {stage1_5[8],stage1_4[54],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage1_5[9],stage1_4[55],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107]},
      {stage1_5[10],stage1_4[56],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113]},
      {stage1_5[11],stage1_4[57],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119]},
      {stage1_5[12],stage1_4[58],stage1_3[61],stage1_2[61],stage1_1[61]}
   );
   gpc606_5 gpc62 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125]},
      {stage1_5[13],stage1_4[59],stage1_3[62],stage1_2[62],stage1_1[62]}
   );
   gpc606_5 gpc63 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[126], stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131]},
      {stage1_5[14],stage1_4[60],stage1_3[63],stage1_2[63],stage1_1[63]}
   );
   gpc606_5 gpc64 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[132], stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137]},
      {stage1_5[15],stage1_4[61],stage1_3[64],stage1_2[64],stage1_1[64]}
   );
   gpc606_5 gpc65 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[138], stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143]},
      {stage1_5[16],stage1_4[62],stage1_3[65],stage1_2[65],stage1_1[65]}
   );
   gpc606_5 gpc66 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[144], stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149]},
      {stage1_5[17],stage1_4[63],stage1_3[66],stage1_2[66],stage1_1[66]}
   );
   gpc606_5 gpc67 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155]},
      {stage1_5[18],stage1_4[64],stage1_3[67],stage1_2[67],stage1_1[67]}
   );
   gpc606_5 gpc68 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161]},
      {stage1_5[19],stage1_4[65],stage1_3[68],stage1_2[68],stage1_1[68]}
   );
   gpc606_5 gpc69 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[162], stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166], stage0_3[167]},
      {stage1_5[20],stage1_4[66],stage1_3[69],stage1_2[69],stage1_1[69]}
   );
   gpc606_5 gpc70 (
      {stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158], stage0_2[159]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[21],stage1_4[67],stage1_3[70],stage1_2[70]}
   );
   gpc606_5 gpc71 (
      {stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164], stage0_2[165]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[22],stage1_4[68],stage1_3[71],stage1_2[71]}
   );
   gpc615_5 gpc72 (
      {stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage0_3[168]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[23],stage1_4[69],stage1_3[72],stage1_2[72]}
   );
   gpc615_5 gpc73 (
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175]},
      {stage0_3[169]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[24],stage1_4[70],stage1_3[73],stage1_2[73]}
   );
   gpc615_5 gpc74 (
      {stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage0_3[170]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[25],stage1_4[71],stage1_3[74],stage1_2[74]}
   );
   gpc615_5 gpc75 (
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185]},
      {stage0_3[171]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[26],stage1_4[72],stage1_3[75],stage1_2[75]}
   );
   gpc615_5 gpc76 (
      {stage0_2[186], stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190]},
      {stage0_3[172]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[27],stage1_4[73],stage1_3[76],stage1_2[76]}
   );
   gpc615_5 gpc77 (
      {stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194], stage0_2[195]},
      {stage0_3[173]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[28],stage1_4[74],stage1_3[77],stage1_2[77]}
   );
   gpc615_5 gpc78 (
      {stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage0_3[174]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[29],stage1_4[75],stage1_3[78],stage1_2[78]}
   );
   gpc615_5 gpc79 (
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205]},
      {stage0_3[175]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[30],stage1_4[76],stage1_3[79],stage1_2[79]}
   );
   gpc615_5 gpc80 (
      {stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage0_3[176]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[31],stage1_4[77],stage1_3[80],stage1_2[80]}
   );
   gpc615_5 gpc81 (
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215]},
      {stage0_3[177]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[32],stage1_4[78],stage1_3[81],stage1_2[81]}
   );
   gpc615_5 gpc82 (
      {stage0_2[216], stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220]},
      {stage0_3[178]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[33],stage1_4[79],stage1_3[82],stage1_2[82]}
   );
   gpc615_5 gpc83 (
      {stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224], stage0_2[225]},
      {stage0_3[179]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[34],stage1_4[80],stage1_3[83],stage1_2[83]}
   );
   gpc615_5 gpc84 (
      {stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage0_3[180]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[35],stage1_4[81],stage1_3[84],stage1_2[84]}
   );
   gpc615_5 gpc85 (
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235]},
      {stage0_3[181]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[36],stage1_4[82],stage1_3[85],stage1_2[85]}
   );
   gpc615_5 gpc86 (
      {stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240]},
      {stage0_3[182]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[37],stage1_4[83],stage1_3[86],stage1_2[86]}
   );
   gpc615_5 gpc87 (
      {stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244], stage0_2[245]},
      {stage0_3[183]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[38],stage1_4[84],stage1_3[87],stage1_2[87]}
   );
   gpc1343_5 gpc88 (
      {stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111]},
      {stage0_5[0], stage0_5[1], stage0_5[2]},
      {stage0_6[0]},
      {stage1_7[0],stage1_6[18],stage1_5[39],stage1_4[85],stage1_3[88]}
   );
   gpc615_5 gpc89 (
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191]},
      {stage0_4[112]},
      {stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage1_7[1],stage1_6[19],stage1_5[40],stage1_4[86],stage1_3[89]}
   );
   gpc615_5 gpc90 (
      {stage0_3[192], stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196]},
      {stage0_4[113]},
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage1_7[2],stage1_6[20],stage1_5[41],stage1_4[87],stage1_3[90]}
   );
   gpc615_5 gpc91 (
      {stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200], stage0_3[201]},
      {stage0_4[114]},
      {stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20]},
      {stage1_7[3],stage1_6[21],stage1_5[42],stage1_4[88],stage1_3[91]}
   );
   gpc615_5 gpc92 (
      {stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage0_4[115]},
      {stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26]},
      {stage1_7[4],stage1_6[22],stage1_5[43],stage1_4[89],stage1_3[92]}
   );
   gpc615_5 gpc93 (
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211]},
      {stage0_4[116]},
      {stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31], stage0_5[32]},
      {stage1_7[5],stage1_6[23],stage1_5[44],stage1_4[90],stage1_3[93]}
   );
   gpc615_5 gpc94 (
      {stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage0_4[117]},
      {stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37], stage0_5[38]},
      {stage1_7[6],stage1_6[24],stage1_5[45],stage1_4[91],stage1_3[94]}
   );
   gpc615_5 gpc95 (
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221]},
      {stage0_4[118]},
      {stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43], stage0_5[44]},
      {stage1_7[7],stage1_6[25],stage1_5[46],stage1_4[92],stage1_3[95]}
   );
   gpc615_5 gpc96 (
      {stage0_3[222], stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226]},
      {stage0_4[119]},
      {stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49], stage0_5[50]},
      {stage1_7[8],stage1_6[26],stage1_5[47],stage1_4[93],stage1_3[96]}
   );
   gpc615_5 gpc97 (
      {stage0_3[227], stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231]},
      {stage0_4[120]},
      {stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55], stage0_5[56]},
      {stage1_7[9],stage1_6[27],stage1_5[48],stage1_4[94],stage1_3[97]}
   );
   gpc615_5 gpc98 (
      {stage0_3[232], stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236]},
      {stage0_4[121]},
      {stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61], stage0_5[62]},
      {stage1_7[10],stage1_6[28],stage1_5[49],stage1_4[95],stage1_3[98]}
   );
   gpc615_5 gpc99 (
      {stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241]},
      {stage0_4[122]},
      {stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66], stage0_5[67], stage0_5[68]},
      {stage1_7[11],stage1_6[29],stage1_5[50],stage1_4[96],stage1_3[99]}
   );
   gpc606_5 gpc100 (
      {stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128]},
      {stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6]},
      {stage1_8[0],stage1_7[12],stage1_6[30],stage1_5[51],stage1_4[97]}
   );
   gpc606_5 gpc101 (
      {stage0_4[129], stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134]},
      {stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11], stage0_6[12]},
      {stage1_8[1],stage1_7[13],stage1_6[31],stage1_5[52],stage1_4[98]}
   );
   gpc606_5 gpc102 (
      {stage0_4[135], stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140]},
      {stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17], stage0_6[18]},
      {stage1_8[2],stage1_7[14],stage1_6[32],stage1_5[53],stage1_4[99]}
   );
   gpc606_5 gpc103 (
      {stage0_4[141], stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146]},
      {stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23], stage0_6[24]},
      {stage1_8[3],stage1_7[15],stage1_6[33],stage1_5[54],stage1_4[100]}
   );
   gpc606_5 gpc104 (
      {stage0_4[147], stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152]},
      {stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29], stage0_6[30]},
      {stage1_8[4],stage1_7[16],stage1_6[34],stage1_5[55],stage1_4[101]}
   );
   gpc606_5 gpc105 (
      {stage0_4[153], stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158]},
      {stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35], stage0_6[36]},
      {stage1_8[5],stage1_7[17],stage1_6[35],stage1_5[56],stage1_4[102]}
   );
   gpc606_5 gpc106 (
      {stage0_4[159], stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164]},
      {stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41], stage0_6[42]},
      {stage1_8[6],stage1_7[18],stage1_6[36],stage1_5[57],stage1_4[103]}
   );
   gpc606_5 gpc107 (
      {stage0_4[165], stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170]},
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47], stage0_6[48]},
      {stage1_8[7],stage1_7[19],stage1_6[37],stage1_5[58],stage1_4[104]}
   );
   gpc606_5 gpc108 (
      {stage0_4[171], stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176]},
      {stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53], stage0_6[54]},
      {stage1_8[8],stage1_7[20],stage1_6[38],stage1_5[59],stage1_4[105]}
   );
   gpc606_5 gpc109 (
      {stage0_4[177], stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182]},
      {stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59], stage0_6[60]},
      {stage1_8[9],stage1_7[21],stage1_6[39],stage1_5[60],stage1_4[106]}
   );
   gpc606_5 gpc110 (
      {stage0_4[183], stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188]},
      {stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65], stage0_6[66]},
      {stage1_8[10],stage1_7[22],stage1_6[40],stage1_5[61],stage1_4[107]}
   );
   gpc615_5 gpc111 (
      {stage0_4[189], stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193]},
      {stage0_5[69]},
      {stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71], stage0_6[72]},
      {stage1_8[11],stage1_7[23],stage1_6[41],stage1_5[62],stage1_4[108]}
   );
   gpc615_5 gpc112 (
      {stage0_4[194], stage0_4[195], stage0_4[196], stage0_4[197], stage0_4[198]},
      {stage0_5[70]},
      {stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77], stage0_6[78]},
      {stage1_8[12],stage1_7[24],stage1_6[42],stage1_5[63],stage1_4[109]}
   );
   gpc615_5 gpc113 (
      {stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202], stage0_4[203]},
      {stage0_5[71]},
      {stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83], stage0_6[84]},
      {stage1_8[13],stage1_7[25],stage1_6[43],stage1_5[64],stage1_4[110]}
   );
   gpc615_5 gpc114 (
      {stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208]},
      {stage0_5[72]},
      {stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89], stage0_6[90]},
      {stage1_8[14],stage1_7[26],stage1_6[44],stage1_5[65],stage1_4[111]}
   );
   gpc615_5 gpc115 (
      {stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213]},
      {stage0_5[73]},
      {stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95], stage0_6[96]},
      {stage1_8[15],stage1_7[27],stage1_6[45],stage1_5[66],stage1_4[112]}
   );
   gpc615_5 gpc116 (
      {stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218]},
      {stage0_5[74]},
      {stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101], stage0_6[102]},
      {stage1_8[16],stage1_7[28],stage1_6[46],stage1_5[67],stage1_4[113]}
   );
   gpc615_5 gpc117 (
      {stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223]},
      {stage0_5[75]},
      {stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107], stage0_6[108]},
      {stage1_8[17],stage1_7[29],stage1_6[47],stage1_5[68],stage1_4[114]}
   );
   gpc615_5 gpc118 (
      {stage0_4[224], stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228]},
      {stage0_5[76]},
      {stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113], stage0_6[114]},
      {stage1_8[18],stage1_7[30],stage1_6[48],stage1_5[69],stage1_4[115]}
   );
   gpc615_5 gpc119 (
      {stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232], stage0_4[233]},
      {stage0_5[77]},
      {stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119], stage0_6[120]},
      {stage1_8[19],stage1_7[31],stage1_6[49],stage1_5[70],stage1_4[116]}
   );
   gpc615_5 gpc120 (
      {stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238]},
      {stage0_5[78]},
      {stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125], stage0_6[126]},
      {stage1_8[20],stage1_7[32],stage1_6[50],stage1_5[71],stage1_4[117]}
   );
   gpc615_5 gpc121 (
      {stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243]},
      {stage0_5[79]},
      {stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131], stage0_6[132]},
      {stage1_8[21],stage1_7[33],stage1_6[51],stage1_5[72],stage1_4[118]}
   );
   gpc615_5 gpc122 (
      {stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248]},
      {stage0_5[80]},
      {stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137], stage0_6[138]},
      {stage1_8[22],stage1_7[34],stage1_6[52],stage1_5[73],stage1_4[119]}
   );
   gpc606_5 gpc123 (
      {stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84], stage0_5[85], stage0_5[86]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[23],stage1_7[35],stage1_6[53],stage1_5[74]}
   );
   gpc606_5 gpc124 (
      {stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90], stage0_5[91], stage0_5[92]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[24],stage1_7[36],stage1_6[54],stage1_5[75]}
   );
   gpc606_5 gpc125 (
      {stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96], stage0_5[97], stage0_5[98]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[25],stage1_7[37],stage1_6[55],stage1_5[76]}
   );
   gpc606_5 gpc126 (
      {stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102], stage0_5[103], stage0_5[104]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[26],stage1_7[38],stage1_6[56],stage1_5[77]}
   );
   gpc606_5 gpc127 (
      {stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108], stage0_5[109], stage0_5[110]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[27],stage1_7[39],stage1_6[57],stage1_5[78]}
   );
   gpc606_5 gpc128 (
      {stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[28],stage1_7[40],stage1_6[58],stage1_5[79]}
   );
   gpc606_5 gpc129 (
      {stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120], stage0_5[121], stage0_5[122]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[29],stage1_7[41],stage1_6[59],stage1_5[80]}
   );
   gpc606_5 gpc130 (
      {stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126], stage0_5[127], stage0_5[128]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[30],stage1_7[42],stage1_6[60],stage1_5[81]}
   );
   gpc606_5 gpc131 (
      {stage0_5[129], stage0_5[130], stage0_5[131], stage0_5[132], stage0_5[133], stage0_5[134]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[31],stage1_7[43],stage1_6[61],stage1_5[82]}
   );
   gpc606_5 gpc132 (
      {stage0_5[135], stage0_5[136], stage0_5[137], stage0_5[138], stage0_5[139], stage0_5[140]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[32],stage1_7[44],stage1_6[62],stage1_5[83]}
   );
   gpc606_5 gpc133 (
      {stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144], stage0_5[145], stage0_5[146]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[33],stage1_7[45],stage1_6[63],stage1_5[84]}
   );
   gpc606_5 gpc134 (
      {stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150], stage0_5[151], stage0_5[152]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[34],stage1_7[46],stage1_6[64],stage1_5[85]}
   );
   gpc606_5 gpc135 (
      {stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156], stage0_5[157], stage0_5[158]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[35],stage1_7[47],stage1_6[65],stage1_5[86]}
   );
   gpc606_5 gpc136 (
      {stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162], stage0_5[163], stage0_5[164]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[36],stage1_7[48],stage1_6[66],stage1_5[87]}
   );
   gpc606_5 gpc137 (
      {stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168], stage0_5[169], stage0_5[170]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[37],stage1_7[49],stage1_6[67],stage1_5[88]}
   );
   gpc606_5 gpc138 (
      {stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174], stage0_5[175], stage0_5[176]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[38],stage1_7[50],stage1_6[68],stage1_5[89]}
   );
   gpc606_5 gpc139 (
      {stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180], stage0_5[181], stage0_5[182]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[39],stage1_7[51],stage1_6[69],stage1_5[90]}
   );
   gpc606_5 gpc140 (
      {stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186], stage0_5[187], stage0_5[188]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[40],stage1_7[52],stage1_6[70],stage1_5[91]}
   );
   gpc606_5 gpc141 (
      {stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192], stage0_5[193], stage0_5[194]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[41],stage1_7[53],stage1_6[71],stage1_5[92]}
   );
   gpc606_5 gpc142 (
      {stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198], stage0_5[199], stage0_5[200]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[42],stage1_7[54],stage1_6[72],stage1_5[93]}
   );
   gpc606_5 gpc143 (
      {stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204], stage0_5[205], stage0_5[206]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[43],stage1_7[55],stage1_6[73],stage1_5[94]}
   );
   gpc606_5 gpc144 (
      {stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210], stage0_5[211], stage0_5[212]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[44],stage1_7[56],stage1_6[74],stage1_5[95]}
   );
   gpc606_5 gpc145 (
      {stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216], stage0_5[217], stage0_5[218]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[45],stage1_7[57],stage1_6[75],stage1_5[96]}
   );
   gpc606_5 gpc146 (
      {stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222], stage0_5[223], stage0_5[224]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[46],stage1_7[58],stage1_6[76],stage1_5[97]}
   );
   gpc606_5 gpc147 (
      {stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228], stage0_5[229], stage0_5[230]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[47],stage1_7[59],stage1_6[77],stage1_5[98]}
   );
   gpc606_5 gpc148 (
      {stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234], stage0_5[235], stage0_5[236]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[48],stage1_7[60],stage1_6[78],stage1_5[99]}
   );
   gpc606_5 gpc149 (
      {stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240], stage0_5[241], stage0_5[242]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[49],stage1_7[61],stage1_6[79],stage1_5[100]}
   );
   gpc606_5 gpc150 (
      {stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246], stage0_5[247], stage0_5[248]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[50],stage1_7[62],stage1_6[80],stage1_5[101]}
   );
   gpc615_5 gpc151 (
      {stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252], stage0_5[253]},
      {stage0_6[139]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[51],stage1_7[63],stage1_6[81],stage1_5[102]}
   );
   gpc606_5 gpc152 (
      {stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143], stage0_6[144], stage0_6[145]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[29],stage1_8[52],stage1_7[64],stage1_6[82]}
   );
   gpc606_5 gpc153 (
      {stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149], stage0_6[150], stage0_6[151]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[30],stage1_8[53],stage1_7[65],stage1_6[83]}
   );
   gpc606_5 gpc154 (
      {stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155], stage0_6[156], stage0_6[157]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[31],stage1_8[54],stage1_7[66],stage1_6[84]}
   );
   gpc606_5 gpc155 (
      {stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161], stage0_6[162], stage0_6[163]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[32],stage1_8[55],stage1_7[67],stage1_6[85]}
   );
   gpc606_5 gpc156 (
      {stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167], stage0_6[168], stage0_6[169]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[33],stage1_8[56],stage1_7[68],stage1_6[86]}
   );
   gpc606_5 gpc157 (
      {stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173], stage0_6[174], stage0_6[175]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[34],stage1_8[57],stage1_7[69],stage1_6[87]}
   );
   gpc606_5 gpc158 (
      {stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179], stage0_6[180], stage0_6[181]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[35],stage1_8[58],stage1_7[70],stage1_6[88]}
   );
   gpc606_5 gpc159 (
      {stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185], stage0_6[186], stage0_6[187]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[36],stage1_8[59],stage1_7[71],stage1_6[89]}
   );
   gpc606_5 gpc160 (
      {stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191], stage0_6[192], stage0_6[193]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[37],stage1_8[60],stage1_7[72],stage1_6[90]}
   );
   gpc606_5 gpc161 (
      {stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197], stage0_6[198], stage0_6[199]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[38],stage1_8[61],stage1_7[73],stage1_6[91]}
   );
   gpc615_5 gpc162 (
      {stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203], stage0_6[204]},
      {stage0_7[174]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[39],stage1_8[62],stage1_7[74],stage1_6[92]}
   );
   gpc615_5 gpc163 (
      {stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage0_7[175]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[40],stage1_8[63],stage1_7[75],stage1_6[93]}
   );
   gpc615_5 gpc164 (
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214]},
      {stage0_7[176]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[41],stage1_8[64],stage1_7[76],stage1_6[94]}
   );
   gpc615_5 gpc165 (
      {stage0_6[215], stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219]},
      {stage0_7[177]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[42],stage1_8[65],stage1_7[77],stage1_6[95]}
   );
   gpc615_5 gpc166 (
      {stage0_6[220], stage0_6[221], stage0_6[222], stage0_6[223], stage0_6[224]},
      {stage0_7[178]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[43],stage1_8[66],stage1_7[78],stage1_6[96]}
   );
   gpc615_5 gpc167 (
      {stage0_6[225], stage0_6[226], stage0_6[227], stage0_6[228], stage0_6[229]},
      {stage0_7[179]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[44],stage1_8[67],stage1_7[79],stage1_6[97]}
   );
   gpc615_5 gpc168 (
      {stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233], stage0_6[234]},
      {stage0_7[180]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[45],stage1_8[68],stage1_7[80],stage1_6[98]}
   );
   gpc615_5 gpc169 (
      {stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage0_7[181]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[46],stage1_8[69],stage1_7[81],stage1_6[99]}
   );
   gpc615_5 gpc170 (
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244]},
      {stage0_7[182]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[47],stage1_8[70],stage1_7[82],stage1_6[100]}
   );
   gpc615_5 gpc171 (
      {stage0_6[245], stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249]},
      {stage0_7[183]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[48],stage1_8[71],stage1_7[83],stage1_6[101]}
   );
   gpc615_5 gpc172 (
      {stage0_6[250], stage0_6[251], stage0_6[252], stage0_6[253], stage0_6[254]},
      {stage0_7[184]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[49],stage1_8[72],stage1_7[84],stage1_6[102]}
   );
   gpc606_5 gpc173 (
      {stage0_7[185], stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[21],stage1_9[50],stage1_8[73],stage1_7[85]}
   );
   gpc615_5 gpc174 (
      {stage0_7[191], stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195]},
      {stage0_8[126]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[22],stage1_9[51],stage1_8[74],stage1_7[86]}
   );
   gpc615_5 gpc175 (
      {stage0_7[196], stage0_7[197], stage0_7[198], stage0_7[199], stage0_7[200]},
      {stage0_8[127]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[23],stage1_9[52],stage1_8[75],stage1_7[87]}
   );
   gpc615_5 gpc176 (
      {stage0_7[201], stage0_7[202], stage0_7[203], stage0_7[204], stage0_7[205]},
      {stage0_8[128]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[24],stage1_9[53],stage1_8[76],stage1_7[88]}
   );
   gpc615_5 gpc177 (
      {stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209], stage0_7[210]},
      {stage0_8[129]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[25],stage1_9[54],stage1_8[77],stage1_7[89]}
   );
   gpc615_5 gpc178 (
      {stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage0_8[130]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[26],stage1_9[55],stage1_8[78],stage1_7[90]}
   );
   gpc615_5 gpc179 (
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220]},
      {stage0_8[131]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[27],stage1_9[56],stage1_8[79],stage1_7[91]}
   );
   gpc615_5 gpc180 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[132]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[28],stage1_9[57],stage1_8[80],stage1_7[92]}
   );
   gpc615_5 gpc181 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[133]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[29],stage1_9[58],stage1_8[81],stage1_7[93]}
   );
   gpc615_5 gpc182 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[134]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[30],stage1_9[59],stage1_8[82],stage1_7[94]}
   );
   gpc606_5 gpc183 (
      {stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[10],stage1_10[31],stage1_9[60],stage1_8[83]}
   );
   gpc606_5 gpc184 (
      {stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[11],stage1_10[32],stage1_9[61],stage1_8[84]}
   );
   gpc606_5 gpc185 (
      {stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151], stage0_8[152]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[12],stage1_10[33],stage1_9[62],stage1_8[85]}
   );
   gpc606_5 gpc186 (
      {stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157], stage0_8[158]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[13],stage1_10[34],stage1_9[63],stage1_8[86]}
   );
   gpc606_5 gpc187 (
      {stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162], stage0_8[163], stage0_8[164]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[14],stage1_10[35],stage1_9[64],stage1_8[87]}
   );
   gpc606_5 gpc188 (
      {stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168], stage0_8[169], stage0_8[170]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[15],stage1_10[36],stage1_9[65],stage1_8[88]}
   );
   gpc606_5 gpc189 (
      {stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174], stage0_8[175], stage0_8[176]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[16],stage1_10[37],stage1_9[66],stage1_8[89]}
   );
   gpc606_5 gpc190 (
      {stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181], stage0_8[182]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[17],stage1_10[38],stage1_9[67],stage1_8[90]}
   );
   gpc606_5 gpc191 (
      {stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187], stage0_8[188]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[18],stage1_10[39],stage1_9[68],stage1_8[91]}
   );
   gpc606_5 gpc192 (
      {stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192], stage0_8[193], stage0_8[194]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[19],stage1_10[40],stage1_9[69],stage1_8[92]}
   );
   gpc615_5 gpc193 (
      {stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198], stage0_8[199]},
      {stage0_9[60]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[20],stage1_10[41],stage1_9[70],stage1_8[93]}
   );
   gpc615_5 gpc194 (
      {stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_9[61]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[21],stage1_10[42],stage1_9[71],stage1_8[94]}
   );
   gpc615_5 gpc195 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage0_9[62]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[22],stage1_10[43],stage1_9[72],stage1_8[95]}
   );
   gpc615_5 gpc196 (
      {stage0_8[210], stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214]},
      {stage0_9[63]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[23],stage1_10[44],stage1_9[73],stage1_8[96]}
   );
   gpc615_5 gpc197 (
      {stage0_8[215], stage0_8[216], stage0_8[217], stage0_8[218], stage0_8[219]},
      {stage0_9[64]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[24],stage1_10[45],stage1_9[74],stage1_8[97]}
   );
   gpc615_5 gpc198 (
      {stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223], stage0_8[224]},
      {stage0_9[65]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[25],stage1_10[46],stage1_9[75],stage1_8[98]}
   );
   gpc615_5 gpc199 (
      {stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229]},
      {stage0_9[66]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[26],stage1_10[47],stage1_9[76],stage1_8[99]}
   );
   gpc615_5 gpc200 (
      {stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234]},
      {stage0_9[67]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[27],stage1_10[48],stage1_9[77],stage1_8[100]}
   );
   gpc615_5 gpc201 (
      {stage0_8[235], stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239]},
      {stage0_9[68]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[28],stage1_10[49],stage1_9[78],stage1_8[101]}
   );
   gpc615_5 gpc202 (
      {stage0_8[240], stage0_8[241], stage0_8[242], stage0_8[243], stage0_8[244]},
      {stage0_9[69]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[29],stage1_10[50],stage1_9[79],stage1_8[102]}
   );
   gpc615_5 gpc203 (
      {stage0_8[245], stage0_8[246], stage0_8[247], stage0_8[248], stage0_8[249]},
      {stage0_9[70]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[30],stage1_10[51],stage1_9[80],stage1_8[103]}
   );
   gpc615_5 gpc204 (
      {stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253], stage0_8[254]},
      {stage0_9[71]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[31],stage1_10[52],stage1_9[81],stage1_8[104]}
   );
   gpc606_5 gpc205 (
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[22],stage1_11[32],stage1_10[53],stage1_9[82]}
   );
   gpc606_5 gpc206 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[23],stage1_11[33],stage1_10[54],stage1_9[83]}
   );
   gpc606_5 gpc207 (
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[24],stage1_11[34],stage1_10[55],stage1_9[84]}
   );
   gpc606_5 gpc208 (
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[25],stage1_11[35],stage1_10[56],stage1_9[85]}
   );
   gpc606_5 gpc209 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[26],stage1_11[36],stage1_10[57],stage1_9[86]}
   );
   gpc606_5 gpc210 (
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[27],stage1_11[37],stage1_10[58],stage1_9[87]}
   );
   gpc606_5 gpc211 (
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[28],stage1_11[38],stage1_10[59],stage1_9[88]}
   );
   gpc606_5 gpc212 (
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[29],stage1_11[39],stage1_10[60],stage1_9[89]}
   );
   gpc606_5 gpc213 (
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[30],stage1_11[40],stage1_10[61],stage1_9[90]}
   );
   gpc606_5 gpc214 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[31],stage1_11[41],stage1_10[62],stage1_9[91]}
   );
   gpc606_5 gpc215 (
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[32],stage1_11[42],stage1_10[63],stage1_9[92]}
   );
   gpc606_5 gpc216 (
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[33],stage1_11[43],stage1_10[64],stage1_9[93]}
   );
   gpc606_5 gpc217 (
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[34],stage1_11[44],stage1_10[65],stage1_9[94]}
   );
   gpc606_5 gpc218 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[35],stage1_11[45],stage1_10[66],stage1_9[95]}
   );
   gpc615_5 gpc219 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_10[132]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[36],stage1_11[46],stage1_10[67],stage1_9[96]}
   );
   gpc615_5 gpc220 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165]},
      {stage0_10[133]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[37],stage1_11[47],stage1_10[68],stage1_9[97]}
   );
   gpc615_5 gpc221 (
      {stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_10[134]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[38],stage1_11[48],stage1_10[69],stage1_9[98]}
   );
   gpc615_5 gpc222 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175]},
      {stage0_10[135]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[39],stage1_11[49],stage1_10[70],stage1_9[99]}
   );
   gpc615_5 gpc223 (
      {stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_10[136]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[40],stage1_11[50],stage1_10[71],stage1_9[100]}
   );
   gpc615_5 gpc224 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_10[137]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[41],stage1_11[51],stage1_10[72],stage1_9[101]}
   );
   gpc615_5 gpc225 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190]},
      {stage0_10[138]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[42],stage1_11[52],stage1_10[73],stage1_9[102]}
   );
   gpc615_5 gpc226 (
      {stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_10[139]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[43],stage1_11[53],stage1_10[74],stage1_9[103]}
   );
   gpc615_5 gpc227 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_10[140]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[44],stage1_11[54],stage1_10[75],stage1_9[104]}
   );
   gpc615_5 gpc228 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205]},
      {stage0_10[141]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[45],stage1_11[55],stage1_10[76],stage1_9[105]}
   );
   gpc615_5 gpc229 (
      {stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_10[142]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[46],stage1_11[56],stage1_10[77],stage1_9[106]}
   );
   gpc615_5 gpc230 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_10[143]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[47],stage1_11[57],stage1_10[78],stage1_9[107]}
   );
   gpc615_5 gpc231 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220]},
      {stage0_10[144]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[48],stage1_11[58],stage1_10[79],stage1_9[108]}
   );
   gpc615_5 gpc232 (
      {stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_10[145]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[49],stage1_11[59],stage1_10[80],stage1_9[109]}
   );
   gpc615_5 gpc233 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_10[146]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[50],stage1_11[60],stage1_10[81],stage1_9[110]}
   );
   gpc615_5 gpc234 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235]},
      {stage0_10[147]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[51],stage1_11[61],stage1_10[82],stage1_9[111]}
   );
   gpc615_5 gpc235 (
      {stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_10[148]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[52],stage1_11[62],stage1_10[83],stage1_9[112]}
   );
   gpc615_5 gpc236 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_10[149]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[53],stage1_11[63],stage1_10[84],stage1_9[113]}
   );
   gpc615_5 gpc237 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250]},
      {stage0_10[150]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[54],stage1_11[64],stage1_10[85],stage1_9[114]}
   );
   gpc615_5 gpc238 (
      {stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_10[151]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[55],stage1_11[65],stage1_10[86],stage1_9[115]}
   );
   gpc606_5 gpc239 (
      {stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155], stage0_10[156], stage0_10[157]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[34],stage1_12[56],stage1_11[66],stage1_10[87]}
   );
   gpc606_5 gpc240 (
      {stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161], stage0_10[162], stage0_10[163]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[35],stage1_12[57],stage1_11[67],stage1_10[88]}
   );
   gpc606_5 gpc241 (
      {stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167], stage0_10[168], stage0_10[169]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[36],stage1_12[58],stage1_11[68],stage1_10[89]}
   );
   gpc606_5 gpc242 (
      {stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173], stage0_10[174], stage0_10[175]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[37],stage1_12[59],stage1_11[69],stage1_10[90]}
   );
   gpc606_5 gpc243 (
      {stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179], stage0_10[180], stage0_10[181]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[38],stage1_12[60],stage1_11[70],stage1_10[91]}
   );
   gpc606_5 gpc244 (
      {stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185], stage0_10[186], stage0_10[187]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[39],stage1_12[61],stage1_11[71],stage1_10[92]}
   );
   gpc606_5 gpc245 (
      {stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191], stage0_10[192], stage0_10[193]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[40],stage1_12[62],stage1_11[72],stage1_10[93]}
   );
   gpc606_5 gpc246 (
      {stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197], stage0_10[198], stage0_10[199]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[41],stage1_12[63],stage1_11[73],stage1_10[94]}
   );
   gpc606_5 gpc247 (
      {stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203], stage0_10[204], stage0_10[205]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[42],stage1_12[64],stage1_11[74],stage1_10[95]}
   );
   gpc606_5 gpc248 (
      {stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209], stage0_10[210], stage0_10[211]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[43],stage1_12[65],stage1_11[75],stage1_10[96]}
   );
   gpc606_5 gpc249 (
      {stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215], stage0_10[216], stage0_10[217]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[44],stage1_12[66],stage1_11[76],stage1_10[97]}
   );
   gpc606_5 gpc250 (
      {stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221], stage0_10[222], stage0_10[223]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[45],stage1_12[67],stage1_11[77],stage1_10[98]}
   );
   gpc606_5 gpc251 (
      {stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227], stage0_10[228], stage0_10[229]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[46],stage1_12[68],stage1_11[78],stage1_10[99]}
   );
   gpc615_5 gpc252 (
      {stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233], stage0_10[234]},
      {stage0_11[204]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[47],stage1_12[69],stage1_11[79],stage1_10[100]}
   );
   gpc615_5 gpc253 (
      {stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage0_11[205]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[48],stage1_12[70],stage1_11[80],stage1_10[101]}
   );
   gpc615_5 gpc254 (
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244]},
      {stage0_11[206]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[49],stage1_12[71],stage1_11[81],stage1_10[102]}
   );
   gpc615_5 gpc255 (
      {stage0_11[207], stage0_11[208], stage0_11[209], stage0_11[210], stage0_11[211]},
      {stage0_12[96]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[16],stage1_13[50],stage1_12[72],stage1_11[82]}
   );
   gpc615_5 gpc256 (
      {stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215], stage0_11[216]},
      {stage0_12[97]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[17],stage1_13[51],stage1_12[73],stage1_11[83]}
   );
   gpc615_5 gpc257 (
      {stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage0_12[98]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[18],stage1_13[52],stage1_12[74],stage1_11[84]}
   );
   gpc615_5 gpc258 (
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226]},
      {stage0_12[99]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[19],stage1_13[53],stage1_12[75],stage1_11[85]}
   );
   gpc606_5 gpc259 (
      {stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[4],stage1_14[20],stage1_13[54],stage1_12[76]}
   );
   gpc606_5 gpc260 (
      {stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[5],stage1_14[21],stage1_13[55],stage1_12[77]}
   );
   gpc606_5 gpc261 (
      {stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[6],stage1_14[22],stage1_13[56],stage1_12[78]}
   );
   gpc606_5 gpc262 (
      {stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[7],stage1_14[23],stage1_13[57],stage1_12[79]}
   );
   gpc606_5 gpc263 (
      {stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[8],stage1_14[24],stage1_13[58],stage1_12[80]}
   );
   gpc606_5 gpc264 (
      {stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[9],stage1_14[25],stage1_13[59],stage1_12[81]}
   );
   gpc606_5 gpc265 (
      {stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[10],stage1_14[26],stage1_13[60],stage1_12[82]}
   );
   gpc606_5 gpc266 (
      {stage0_12[142], stage0_12[143], stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[11],stage1_14[27],stage1_13[61],stage1_12[83]}
   );
   gpc606_5 gpc267 (
      {stage0_12[148], stage0_12[149], stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[12],stage1_14[28],stage1_13[62],stage1_12[84]}
   );
   gpc606_5 gpc268 (
      {stage0_12[154], stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[13],stage1_14[29],stage1_13[63],stage1_12[85]}
   );
   gpc606_5 gpc269 (
      {stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[14],stage1_14[30],stage1_13[64],stage1_12[86]}
   );
   gpc606_5 gpc270 (
      {stage0_12[166], stage0_12[167], stage0_12[168], stage0_12[169], stage0_12[170], stage0_12[171]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[15],stage1_14[31],stage1_13[65],stage1_12[87]}
   );
   gpc606_5 gpc271 (
      {stage0_12[172], stage0_12[173], stage0_12[174], stage0_12[175], stage0_12[176], stage0_12[177]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[16],stage1_14[32],stage1_13[66],stage1_12[88]}
   );
   gpc606_5 gpc272 (
      {stage0_12[178], stage0_12[179], stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[17],stage1_14[33],stage1_13[67],stage1_12[89]}
   );
   gpc606_5 gpc273 (
      {stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[18],stage1_14[34],stage1_13[68],stage1_12[90]}
   );
   gpc606_5 gpc274 (
      {stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193], stage0_12[194], stage0_12[195]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[19],stage1_14[35],stage1_13[69],stage1_12[91]}
   );
   gpc606_5 gpc275 (
      {stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199], stage0_12[200], stage0_12[201]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[20],stage1_14[36],stage1_13[70],stage1_12[92]}
   );
   gpc606_5 gpc276 (
      {stage0_12[202], stage0_12[203], stage0_12[204], stage0_12[205], stage0_12[206], stage0_12[207]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[21],stage1_14[37],stage1_13[71],stage1_12[93]}
   );
   gpc606_5 gpc277 (
      {stage0_12[208], stage0_12[209], stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[22],stage1_14[38],stage1_13[72],stage1_12[94]}
   );
   gpc606_5 gpc278 (
      {stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[23],stage1_14[39],stage1_13[73],stage1_12[95]}
   );
   gpc606_5 gpc279 (
      {stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223], stage0_12[224], stage0_12[225]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[24],stage1_14[40],stage1_13[74],stage1_12[96]}
   );
   gpc606_5 gpc280 (
      {stage0_12[226], stage0_12[227], stage0_12[228], stage0_12[229], stage0_12[230], stage0_12[231]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[25],stage1_14[41],stage1_13[75],stage1_12[97]}
   );
   gpc606_5 gpc281 (
      {stage0_12[232], stage0_12[233], stage0_12[234], stage0_12[235], stage0_12[236], stage0_12[237]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[26],stage1_14[42],stage1_13[76],stage1_12[98]}
   );
   gpc606_5 gpc282 (
      {stage0_12[238], stage0_12[239], stage0_12[240], stage0_12[241], stage0_12[242], stage0_12[243]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[27],stage1_14[43],stage1_13[77],stage1_12[99]}
   );
   gpc606_5 gpc283 (
      {stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247], stage0_12[248], stage0_12[249]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[28],stage1_14[44],stage1_13[78],stage1_12[100]}
   );
   gpc606_5 gpc284 (
      {stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253], stage0_12[254], stage0_12[255]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[29],stage1_14[45],stage1_13[79],stage1_12[101]}
   );
   gpc606_5 gpc285 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[26],stage1_15[30],stage1_14[46],stage1_13[80]}
   );
   gpc606_5 gpc286 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[27],stage1_15[31],stage1_14[47],stage1_13[81]}
   );
   gpc606_5 gpc287 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[28],stage1_15[32],stage1_14[48],stage1_13[82]}
   );
   gpc606_5 gpc288 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[29],stage1_15[33],stage1_14[49],stage1_13[83]}
   );
   gpc606_5 gpc289 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[30],stage1_15[34],stage1_14[50],stage1_13[84]}
   );
   gpc606_5 gpc290 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[31],stage1_15[35],stage1_14[51],stage1_13[85]}
   );
   gpc606_5 gpc291 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[32],stage1_15[36],stage1_14[52],stage1_13[86]}
   );
   gpc606_5 gpc292 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[33],stage1_15[37],stage1_14[53],stage1_13[87]}
   );
   gpc606_5 gpc293 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[34],stage1_15[38],stage1_14[54],stage1_13[88]}
   );
   gpc606_5 gpc294 (
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[35],stage1_15[39],stage1_14[55],stage1_13[89]}
   );
   gpc606_5 gpc295 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[36],stage1_15[40],stage1_14[56],stage1_13[90]}
   );
   gpc615_5 gpc296 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94]},
      {stage0_14[156]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[37],stage1_15[41],stage1_14[57],stage1_13[91]}
   );
   gpc615_5 gpc297 (
      {stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99]},
      {stage0_14[157]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[38],stage1_15[42],stage1_14[58],stage1_13[92]}
   );
   gpc615_5 gpc298 (
      {stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103], stage0_13[104]},
      {stage0_14[158]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[39],stage1_15[43],stage1_14[59],stage1_13[93]}
   );
   gpc615_5 gpc299 (
      {stage0_13[105], stage0_13[106], stage0_13[107], stage0_13[108], stage0_13[109]},
      {stage0_14[159]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[40],stage1_15[44],stage1_14[60],stage1_13[94]}
   );
   gpc615_5 gpc300 (
      {stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113], stage0_13[114]},
      {stage0_14[160]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[41],stage1_15[45],stage1_14[61],stage1_13[95]}
   );
   gpc615_5 gpc301 (
      {stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_14[161]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[42],stage1_15[46],stage1_14[62],stage1_13[96]}
   );
   gpc615_5 gpc302 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124]},
      {stage0_14[162]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[43],stage1_15[47],stage1_14[63],stage1_13[97]}
   );
   gpc615_5 gpc303 (
      {stage0_13[125], stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129]},
      {stage0_14[163]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[44],stage1_15[48],stage1_14[64],stage1_13[98]}
   );
   gpc615_5 gpc304 (
      {stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133], stage0_13[134]},
      {stage0_14[164]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[45],stage1_15[49],stage1_14[65],stage1_13[99]}
   );
   gpc615_5 gpc305 (
      {stage0_13[135], stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139]},
      {stage0_14[165]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[46],stage1_15[50],stage1_14[66],stage1_13[100]}
   );
   gpc615_5 gpc306 (
      {stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143], stage0_13[144]},
      {stage0_14[166]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[47],stage1_15[51],stage1_14[67],stage1_13[101]}
   );
   gpc615_5 gpc307 (
      {stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_14[167]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[48],stage1_15[52],stage1_14[68],stage1_13[102]}
   );
   gpc615_5 gpc308 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154]},
      {stage0_14[168]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[49],stage1_15[53],stage1_14[69],stage1_13[103]}
   );
   gpc615_5 gpc309 (
      {stage0_13[155], stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159]},
      {stage0_14[169]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[50],stage1_15[54],stage1_14[70],stage1_13[104]}
   );
   gpc615_5 gpc310 (
      {stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163], stage0_13[164]},
      {stage0_14[170]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[51],stage1_15[55],stage1_14[71],stage1_13[105]}
   );
   gpc615_5 gpc311 (
      {stage0_13[165], stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169]},
      {stage0_14[171]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[52],stage1_15[56],stage1_14[72],stage1_13[106]}
   );
   gpc615_5 gpc312 (
      {stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174]},
      {stage0_14[172]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[53],stage1_15[57],stage1_14[73],stage1_13[107]}
   );
   gpc615_5 gpc313 (
      {stage0_13[175], stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179]},
      {stage0_14[173]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[54],stage1_15[58],stage1_14[74],stage1_13[108]}
   );
   gpc615_5 gpc314 (
      {stage0_13[180], stage0_13[181], stage0_13[182], stage0_13[183], stage0_13[184]},
      {stage0_14[174]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[55],stage1_15[59],stage1_14[75],stage1_13[109]}
   );
   gpc615_5 gpc315 (
      {stage0_13[185], stage0_13[186], stage0_13[187], stage0_13[188], stage0_13[189]},
      {stage0_14[175]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[56],stage1_15[60],stage1_14[76],stage1_13[110]}
   );
   gpc615_5 gpc316 (
      {stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193], stage0_13[194]},
      {stage0_14[176]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[57],stage1_15[61],stage1_14[77],stage1_13[111]}
   );
   gpc615_5 gpc317 (
      {stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199]},
      {stage0_14[177]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[58],stage1_15[62],stage1_14[78],stage1_13[112]}
   );
   gpc615_5 gpc318 (
      {stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204]},
      {stage0_14[178]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[59],stage1_15[63],stage1_14[79],stage1_13[113]}
   );
   gpc615_5 gpc319 (
      {stage0_13[205], stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209]},
      {stage0_14[179]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[60],stage1_15[64],stage1_14[80],stage1_13[114]}
   );
   gpc615_5 gpc320 (
      {stage0_13[210], stage0_13[211], stage0_13[212], stage0_13[213], stage0_13[214]},
      {stage0_14[180]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[61],stage1_15[65],stage1_14[81],stage1_13[115]}
   );
   gpc615_5 gpc321 (
      {stage0_13[215], stage0_13[216], stage0_13[217], stage0_13[218], stage0_13[219]},
      {stage0_14[181]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[62],stage1_15[66],stage1_14[82],stage1_13[116]}
   );
   gpc615_5 gpc322 (
      {stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223], stage0_13[224]},
      {stage0_14[182]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[63],stage1_15[67],stage1_14[83],stage1_13[117]}
   );
   gpc615_5 gpc323 (
      {stage0_13[225], stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229]},
      {stage0_14[183]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[64],stage1_15[68],stage1_14[84],stage1_13[118]}
   );
   gpc615_5 gpc324 (
      {stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234]},
      {stage0_14[184]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[65],stage1_15[69],stage1_14[85],stage1_13[119]}
   );
   gpc615_5 gpc325 (
      {stage0_13[235], stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239]},
      {stage0_14[185]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[66],stage1_15[70],stage1_14[86],stage1_13[120]}
   );
   gpc615_5 gpc326 (
      {stage0_13[240], stage0_13[241], stage0_13[242], stage0_13[243], stage0_13[244]},
      {stage0_14[186]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[67],stage1_15[71],stage1_14[87],stage1_13[121]}
   );
   gpc1_1 gpc327 (
      {stage0_1[228]},
      {stage1_1[70]}
   );
   gpc1_1 gpc328 (
      {stage0_1[229]},
      {stage1_1[71]}
   );
   gpc1_1 gpc329 (
      {stage0_1[230]},
      {stage1_1[72]}
   );
   gpc1_1 gpc330 (
      {stage0_1[231]},
      {stage1_1[73]}
   );
   gpc1_1 gpc331 (
      {stage0_1[232]},
      {stage1_1[74]}
   );
   gpc1_1 gpc332 (
      {stage0_1[233]},
      {stage1_1[75]}
   );
   gpc1_1 gpc333 (
      {stage0_1[234]},
      {stage1_1[76]}
   );
   gpc1_1 gpc334 (
      {stage0_1[235]},
      {stage1_1[77]}
   );
   gpc1_1 gpc335 (
      {stage0_1[236]},
      {stage1_1[78]}
   );
   gpc1_1 gpc336 (
      {stage0_1[237]},
      {stage1_1[79]}
   );
   gpc1_1 gpc337 (
      {stage0_1[238]},
      {stage1_1[80]}
   );
   gpc1_1 gpc338 (
      {stage0_1[239]},
      {stage1_1[81]}
   );
   gpc1_1 gpc339 (
      {stage0_1[240]},
      {stage1_1[82]}
   );
   gpc1_1 gpc340 (
      {stage0_1[241]},
      {stage1_1[83]}
   );
   gpc1_1 gpc341 (
      {stage0_1[242]},
      {stage1_1[84]}
   );
   gpc1_1 gpc342 (
      {stage0_1[243]},
      {stage1_1[85]}
   );
   gpc1_1 gpc343 (
      {stage0_1[244]},
      {stage1_1[86]}
   );
   gpc1_1 gpc344 (
      {stage0_1[245]},
      {stage1_1[87]}
   );
   gpc1_1 gpc345 (
      {stage0_1[246]},
      {stage1_1[88]}
   );
   gpc1_1 gpc346 (
      {stage0_1[247]},
      {stage1_1[89]}
   );
   gpc1_1 gpc347 (
      {stage0_1[248]},
      {stage1_1[90]}
   );
   gpc1_1 gpc348 (
      {stage0_1[249]},
      {stage1_1[91]}
   );
   gpc1_1 gpc349 (
      {stage0_1[250]},
      {stage1_1[92]}
   );
   gpc1_1 gpc350 (
      {stage0_1[251]},
      {stage1_1[93]}
   );
   gpc1_1 gpc351 (
      {stage0_1[252]},
      {stage1_1[94]}
   );
   gpc1_1 gpc352 (
      {stage0_1[253]},
      {stage1_1[95]}
   );
   gpc1_1 gpc353 (
      {stage0_1[254]},
      {stage1_1[96]}
   );
   gpc1_1 gpc354 (
      {stage0_1[255]},
      {stage1_1[97]}
   );
   gpc1_1 gpc355 (
      {stage0_2[246]},
      {stage1_2[88]}
   );
   gpc1_1 gpc356 (
      {stage0_2[247]},
      {stage1_2[89]}
   );
   gpc1_1 gpc357 (
      {stage0_2[248]},
      {stage1_2[90]}
   );
   gpc1_1 gpc358 (
      {stage0_2[249]},
      {stage1_2[91]}
   );
   gpc1_1 gpc359 (
      {stage0_2[250]},
      {stage1_2[92]}
   );
   gpc1_1 gpc360 (
      {stage0_2[251]},
      {stage1_2[93]}
   );
   gpc1_1 gpc361 (
      {stage0_2[252]},
      {stage1_2[94]}
   );
   gpc1_1 gpc362 (
      {stage0_2[253]},
      {stage1_2[95]}
   );
   gpc1_1 gpc363 (
      {stage0_2[254]},
      {stage1_2[96]}
   );
   gpc1_1 gpc364 (
      {stage0_2[255]},
      {stage1_2[97]}
   );
   gpc1_1 gpc365 (
      {stage0_3[242]},
      {stage1_3[100]}
   );
   gpc1_1 gpc366 (
      {stage0_3[243]},
      {stage1_3[101]}
   );
   gpc1_1 gpc367 (
      {stage0_3[244]},
      {stage1_3[102]}
   );
   gpc1_1 gpc368 (
      {stage0_3[245]},
      {stage1_3[103]}
   );
   gpc1_1 gpc369 (
      {stage0_3[246]},
      {stage1_3[104]}
   );
   gpc1_1 gpc370 (
      {stage0_3[247]},
      {stage1_3[105]}
   );
   gpc1_1 gpc371 (
      {stage0_3[248]},
      {stage1_3[106]}
   );
   gpc1_1 gpc372 (
      {stage0_3[249]},
      {stage1_3[107]}
   );
   gpc1_1 gpc373 (
      {stage0_3[250]},
      {stage1_3[108]}
   );
   gpc1_1 gpc374 (
      {stage0_3[251]},
      {stage1_3[109]}
   );
   gpc1_1 gpc375 (
      {stage0_3[252]},
      {stage1_3[110]}
   );
   gpc1_1 gpc376 (
      {stage0_3[253]},
      {stage1_3[111]}
   );
   gpc1_1 gpc377 (
      {stage0_3[254]},
      {stage1_3[112]}
   );
   gpc1_1 gpc378 (
      {stage0_3[255]},
      {stage1_3[113]}
   );
   gpc1_1 gpc379 (
      {stage0_4[249]},
      {stage1_4[120]}
   );
   gpc1_1 gpc380 (
      {stage0_4[250]},
      {stage1_4[121]}
   );
   gpc1_1 gpc381 (
      {stage0_4[251]},
      {stage1_4[122]}
   );
   gpc1_1 gpc382 (
      {stage0_4[252]},
      {stage1_4[123]}
   );
   gpc1_1 gpc383 (
      {stage0_4[253]},
      {stage1_4[124]}
   );
   gpc1_1 gpc384 (
      {stage0_4[254]},
      {stage1_4[125]}
   );
   gpc1_1 gpc385 (
      {stage0_4[255]},
      {stage1_4[126]}
   );
   gpc1_1 gpc386 (
      {stage0_5[254]},
      {stage1_5[103]}
   );
   gpc1_1 gpc387 (
      {stage0_5[255]},
      {stage1_5[104]}
   );
   gpc1_1 gpc388 (
      {stage0_6[255]},
      {stage1_6[103]}
   );
   gpc1_1 gpc389 (
      {stage0_7[236]},
      {stage1_7[95]}
   );
   gpc1_1 gpc390 (
      {stage0_7[237]},
      {stage1_7[96]}
   );
   gpc1_1 gpc391 (
      {stage0_7[238]},
      {stage1_7[97]}
   );
   gpc1_1 gpc392 (
      {stage0_7[239]},
      {stage1_7[98]}
   );
   gpc1_1 gpc393 (
      {stage0_7[240]},
      {stage1_7[99]}
   );
   gpc1_1 gpc394 (
      {stage0_7[241]},
      {stage1_7[100]}
   );
   gpc1_1 gpc395 (
      {stage0_7[242]},
      {stage1_7[101]}
   );
   gpc1_1 gpc396 (
      {stage0_7[243]},
      {stage1_7[102]}
   );
   gpc1_1 gpc397 (
      {stage0_7[244]},
      {stage1_7[103]}
   );
   gpc1_1 gpc398 (
      {stage0_7[245]},
      {stage1_7[104]}
   );
   gpc1_1 gpc399 (
      {stage0_7[246]},
      {stage1_7[105]}
   );
   gpc1_1 gpc400 (
      {stage0_7[247]},
      {stage1_7[106]}
   );
   gpc1_1 gpc401 (
      {stage0_7[248]},
      {stage1_7[107]}
   );
   gpc1_1 gpc402 (
      {stage0_7[249]},
      {stage1_7[108]}
   );
   gpc1_1 gpc403 (
      {stage0_7[250]},
      {stage1_7[109]}
   );
   gpc1_1 gpc404 (
      {stage0_7[251]},
      {stage1_7[110]}
   );
   gpc1_1 gpc405 (
      {stage0_7[252]},
      {stage1_7[111]}
   );
   gpc1_1 gpc406 (
      {stage0_7[253]},
      {stage1_7[112]}
   );
   gpc1_1 gpc407 (
      {stage0_7[254]},
      {stage1_7[113]}
   );
   gpc1_1 gpc408 (
      {stage0_7[255]},
      {stage1_7[114]}
   );
   gpc1_1 gpc409 (
      {stage0_8[255]},
      {stage1_8[105]}
   );
   gpc1_1 gpc410 (
      {stage0_10[245]},
      {stage1_10[103]}
   );
   gpc1_1 gpc411 (
      {stage0_10[246]},
      {stage1_10[104]}
   );
   gpc1_1 gpc412 (
      {stage0_10[247]},
      {stage1_10[105]}
   );
   gpc1_1 gpc413 (
      {stage0_10[248]},
      {stage1_10[106]}
   );
   gpc1_1 gpc414 (
      {stage0_10[249]},
      {stage1_10[107]}
   );
   gpc1_1 gpc415 (
      {stage0_10[250]},
      {stage1_10[108]}
   );
   gpc1_1 gpc416 (
      {stage0_10[251]},
      {stage1_10[109]}
   );
   gpc1_1 gpc417 (
      {stage0_10[252]},
      {stage1_10[110]}
   );
   gpc1_1 gpc418 (
      {stage0_10[253]},
      {stage1_10[111]}
   );
   gpc1_1 gpc419 (
      {stage0_10[254]},
      {stage1_10[112]}
   );
   gpc1_1 gpc420 (
      {stage0_10[255]},
      {stage1_10[113]}
   );
   gpc1_1 gpc421 (
      {stage0_11[227]},
      {stage1_11[86]}
   );
   gpc1_1 gpc422 (
      {stage0_11[228]},
      {stage1_11[87]}
   );
   gpc1_1 gpc423 (
      {stage0_11[229]},
      {stage1_11[88]}
   );
   gpc1_1 gpc424 (
      {stage0_11[230]},
      {stage1_11[89]}
   );
   gpc1_1 gpc425 (
      {stage0_11[231]},
      {stage1_11[90]}
   );
   gpc1_1 gpc426 (
      {stage0_11[232]},
      {stage1_11[91]}
   );
   gpc1_1 gpc427 (
      {stage0_11[233]},
      {stage1_11[92]}
   );
   gpc1_1 gpc428 (
      {stage0_11[234]},
      {stage1_11[93]}
   );
   gpc1_1 gpc429 (
      {stage0_11[235]},
      {stage1_11[94]}
   );
   gpc1_1 gpc430 (
      {stage0_11[236]},
      {stage1_11[95]}
   );
   gpc1_1 gpc431 (
      {stage0_11[237]},
      {stage1_11[96]}
   );
   gpc1_1 gpc432 (
      {stage0_11[238]},
      {stage1_11[97]}
   );
   gpc1_1 gpc433 (
      {stage0_11[239]},
      {stage1_11[98]}
   );
   gpc1_1 gpc434 (
      {stage0_11[240]},
      {stage1_11[99]}
   );
   gpc1_1 gpc435 (
      {stage0_11[241]},
      {stage1_11[100]}
   );
   gpc1_1 gpc436 (
      {stage0_11[242]},
      {stage1_11[101]}
   );
   gpc1_1 gpc437 (
      {stage0_11[243]},
      {stage1_11[102]}
   );
   gpc1_1 gpc438 (
      {stage0_11[244]},
      {stage1_11[103]}
   );
   gpc1_1 gpc439 (
      {stage0_11[245]},
      {stage1_11[104]}
   );
   gpc1_1 gpc440 (
      {stage0_11[246]},
      {stage1_11[105]}
   );
   gpc1_1 gpc441 (
      {stage0_11[247]},
      {stage1_11[106]}
   );
   gpc1_1 gpc442 (
      {stage0_11[248]},
      {stage1_11[107]}
   );
   gpc1_1 gpc443 (
      {stage0_11[249]},
      {stage1_11[108]}
   );
   gpc1_1 gpc444 (
      {stage0_11[250]},
      {stage1_11[109]}
   );
   gpc1_1 gpc445 (
      {stage0_11[251]},
      {stage1_11[110]}
   );
   gpc1_1 gpc446 (
      {stage0_11[252]},
      {stage1_11[111]}
   );
   gpc1_1 gpc447 (
      {stage0_11[253]},
      {stage1_11[112]}
   );
   gpc1_1 gpc448 (
      {stage0_11[254]},
      {stage1_11[113]}
   );
   gpc1_1 gpc449 (
      {stage0_11[255]},
      {stage1_11[114]}
   );
   gpc1_1 gpc450 (
      {stage0_13[245]},
      {stage1_13[122]}
   );
   gpc1_1 gpc451 (
      {stage0_13[246]},
      {stage1_13[123]}
   );
   gpc1_1 gpc452 (
      {stage0_13[247]},
      {stage1_13[124]}
   );
   gpc1_1 gpc453 (
      {stage0_13[248]},
      {stage1_13[125]}
   );
   gpc1_1 gpc454 (
      {stage0_13[249]},
      {stage1_13[126]}
   );
   gpc1_1 gpc455 (
      {stage0_13[250]},
      {stage1_13[127]}
   );
   gpc1_1 gpc456 (
      {stage0_13[251]},
      {stage1_13[128]}
   );
   gpc1_1 gpc457 (
      {stage0_13[252]},
      {stage1_13[129]}
   );
   gpc1_1 gpc458 (
      {stage0_13[253]},
      {stage1_13[130]}
   );
   gpc1_1 gpc459 (
      {stage0_13[254]},
      {stage1_13[131]}
   );
   gpc1_1 gpc460 (
      {stage0_13[255]},
      {stage1_13[132]}
   );
   gpc1_1 gpc461 (
      {stage0_14[187]},
      {stage1_14[88]}
   );
   gpc1_1 gpc462 (
      {stage0_14[188]},
      {stage1_14[89]}
   );
   gpc1_1 gpc463 (
      {stage0_14[189]},
      {stage1_14[90]}
   );
   gpc1_1 gpc464 (
      {stage0_14[190]},
      {stage1_14[91]}
   );
   gpc1_1 gpc465 (
      {stage0_14[191]},
      {stage1_14[92]}
   );
   gpc1_1 gpc466 (
      {stage0_14[192]},
      {stage1_14[93]}
   );
   gpc1_1 gpc467 (
      {stage0_14[193]},
      {stage1_14[94]}
   );
   gpc1_1 gpc468 (
      {stage0_14[194]},
      {stage1_14[95]}
   );
   gpc1_1 gpc469 (
      {stage0_14[195]},
      {stage1_14[96]}
   );
   gpc1_1 gpc470 (
      {stage0_14[196]},
      {stage1_14[97]}
   );
   gpc1_1 gpc471 (
      {stage0_14[197]},
      {stage1_14[98]}
   );
   gpc1_1 gpc472 (
      {stage0_14[198]},
      {stage1_14[99]}
   );
   gpc1_1 gpc473 (
      {stage0_14[199]},
      {stage1_14[100]}
   );
   gpc1_1 gpc474 (
      {stage0_14[200]},
      {stage1_14[101]}
   );
   gpc1_1 gpc475 (
      {stage0_14[201]},
      {stage1_14[102]}
   );
   gpc1_1 gpc476 (
      {stage0_14[202]},
      {stage1_14[103]}
   );
   gpc1_1 gpc477 (
      {stage0_14[203]},
      {stage1_14[104]}
   );
   gpc1_1 gpc478 (
      {stage0_14[204]},
      {stage1_14[105]}
   );
   gpc1_1 gpc479 (
      {stage0_14[205]},
      {stage1_14[106]}
   );
   gpc1_1 gpc480 (
      {stage0_14[206]},
      {stage1_14[107]}
   );
   gpc1_1 gpc481 (
      {stage0_14[207]},
      {stage1_14[108]}
   );
   gpc1_1 gpc482 (
      {stage0_14[208]},
      {stage1_14[109]}
   );
   gpc1_1 gpc483 (
      {stage0_14[209]},
      {stage1_14[110]}
   );
   gpc1_1 gpc484 (
      {stage0_14[210]},
      {stage1_14[111]}
   );
   gpc1_1 gpc485 (
      {stage0_14[211]},
      {stage1_14[112]}
   );
   gpc1_1 gpc486 (
      {stage0_14[212]},
      {stage1_14[113]}
   );
   gpc1_1 gpc487 (
      {stage0_14[213]},
      {stage1_14[114]}
   );
   gpc1_1 gpc488 (
      {stage0_14[214]},
      {stage1_14[115]}
   );
   gpc1_1 gpc489 (
      {stage0_14[215]},
      {stage1_14[116]}
   );
   gpc1_1 gpc490 (
      {stage0_14[216]},
      {stage1_14[117]}
   );
   gpc1_1 gpc491 (
      {stage0_14[217]},
      {stage1_14[118]}
   );
   gpc1_1 gpc492 (
      {stage0_14[218]},
      {stage1_14[119]}
   );
   gpc1_1 gpc493 (
      {stage0_14[219]},
      {stage1_14[120]}
   );
   gpc1_1 gpc494 (
      {stage0_14[220]},
      {stage1_14[121]}
   );
   gpc1_1 gpc495 (
      {stage0_14[221]},
      {stage1_14[122]}
   );
   gpc1_1 gpc496 (
      {stage0_14[222]},
      {stage1_14[123]}
   );
   gpc1_1 gpc497 (
      {stage0_14[223]},
      {stage1_14[124]}
   );
   gpc1_1 gpc498 (
      {stage0_14[224]},
      {stage1_14[125]}
   );
   gpc1_1 gpc499 (
      {stage0_14[225]},
      {stage1_14[126]}
   );
   gpc1_1 gpc500 (
      {stage0_14[226]},
      {stage1_14[127]}
   );
   gpc1_1 gpc501 (
      {stage0_14[227]},
      {stage1_14[128]}
   );
   gpc1_1 gpc502 (
      {stage0_14[228]},
      {stage1_14[129]}
   );
   gpc1_1 gpc503 (
      {stage0_14[229]},
      {stage1_14[130]}
   );
   gpc1_1 gpc504 (
      {stage0_14[230]},
      {stage1_14[131]}
   );
   gpc1_1 gpc505 (
      {stage0_14[231]},
      {stage1_14[132]}
   );
   gpc1_1 gpc506 (
      {stage0_14[232]},
      {stage1_14[133]}
   );
   gpc1_1 gpc507 (
      {stage0_14[233]},
      {stage1_14[134]}
   );
   gpc1_1 gpc508 (
      {stage0_14[234]},
      {stage1_14[135]}
   );
   gpc1_1 gpc509 (
      {stage0_14[235]},
      {stage1_14[136]}
   );
   gpc1_1 gpc510 (
      {stage0_14[236]},
      {stage1_14[137]}
   );
   gpc1_1 gpc511 (
      {stage0_14[237]},
      {stage1_14[138]}
   );
   gpc1_1 gpc512 (
      {stage0_14[238]},
      {stage1_14[139]}
   );
   gpc1_1 gpc513 (
      {stage0_14[239]},
      {stage1_14[140]}
   );
   gpc1_1 gpc514 (
      {stage0_14[240]},
      {stage1_14[141]}
   );
   gpc1_1 gpc515 (
      {stage0_14[241]},
      {stage1_14[142]}
   );
   gpc1_1 gpc516 (
      {stage0_14[242]},
      {stage1_14[143]}
   );
   gpc1_1 gpc517 (
      {stage0_14[243]},
      {stage1_14[144]}
   );
   gpc1_1 gpc518 (
      {stage0_14[244]},
      {stage1_14[145]}
   );
   gpc1_1 gpc519 (
      {stage0_14[245]},
      {stage1_14[146]}
   );
   gpc1_1 gpc520 (
      {stage0_14[246]},
      {stage1_14[147]}
   );
   gpc1_1 gpc521 (
      {stage0_14[247]},
      {stage1_14[148]}
   );
   gpc1_1 gpc522 (
      {stage0_14[248]},
      {stage1_14[149]}
   );
   gpc1_1 gpc523 (
      {stage0_14[249]},
      {stage1_14[150]}
   );
   gpc1_1 gpc524 (
      {stage0_14[250]},
      {stage1_14[151]}
   );
   gpc1_1 gpc525 (
      {stage0_14[251]},
      {stage1_14[152]}
   );
   gpc1_1 gpc526 (
      {stage0_14[252]},
      {stage1_14[153]}
   );
   gpc1_1 gpc527 (
      {stage0_14[253]},
      {stage1_14[154]}
   );
   gpc1_1 gpc528 (
      {stage0_14[254]},
      {stage1_14[155]}
   );
   gpc1_1 gpc529 (
      {stage0_14[255]},
      {stage1_14[156]}
   );
   gpc1_1 gpc530 (
      {stage0_15[252]},
      {stage1_15[72]}
   );
   gpc1_1 gpc531 (
      {stage0_15[253]},
      {stage1_15[73]}
   );
   gpc1_1 gpc532 (
      {stage0_15[254]},
      {stage1_15[74]}
   );
   gpc1_1 gpc533 (
      {stage0_15[255]},
      {stage1_15[75]}
   );
   gpc606_5 gpc534 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc535 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc536 (
      {stage1_0[12], stage1_0[13], stage1_0[14], stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc537 (
      {stage1_0[18], stage1_0[19], stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc538 (
      {stage1_0[24], stage1_0[25], stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc539 (
      {stage1_0[30], stage1_0[31], stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc540 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc541 (
      {stage1_0[42], stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc542 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc606_5 gpc543 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9]}
   );
   gpc606_5 gpc544 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10]}
   );
   gpc606_5 gpc545 (
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11]}
   );
   gpc606_5 gpc546 (
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29]},
      {stage2_5[4],stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12]}
   );
   gpc606_5 gpc547 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage2_5[5],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc548 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage2_5[6],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc549 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage2_5[7],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc606_5 gpc550 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage2_5[8],stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16]}
   );
   gpc606_5 gpc551 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59]},
      {stage2_5[9],stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17]}
   );
   gpc606_5 gpc552 (
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage2_5[10],stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18]}
   );
   gpc606_5 gpc553 (
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage2_5[11],stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19]}
   );
   gpc606_5 gpc554 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77]},
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77]},
      {stage2_5[12],stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20]}
   );
   gpc606_5 gpc555 (
      {stage1_1[78], stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83]},
      {stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage2_5[13],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc606_5 gpc556 (
      {stage1_1[84], stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89]},
      {stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89]},
      {stage2_5[14],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc606_5 gpc557 (
      {stage1_1[90], stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95]},
      {stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage2_5[15],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc558 (
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[16],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc606_5 gpc559 (
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[17],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc606_5 gpc560 (
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[18],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc606_5 gpc561 (
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[19],stage2_4[27],stage2_3[27],stage2_2[27]}
   );
   gpc615_5 gpc562 (
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76]},
      {stage1_3[96]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[20],stage2_4[28],stage2_3[28],stage2_2[28]}
   );
   gpc615_5 gpc563 (
      {stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81]},
      {stage1_3[97]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[21],stage2_4[29],stage2_3[29],stage2_2[29]}
   );
   gpc615_5 gpc564 (
      {stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101], stage1_3[102]},
      {stage1_4[36]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[6],stage2_5[22],stage2_4[30],stage2_3[30]}
   );
   gpc615_5 gpc565 (
      {stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage1_4[37]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[7],stage2_5[23],stage2_4[31],stage2_3[31]}
   );
   gpc615_5 gpc566 (
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112]},
      {stage1_4[38]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[8],stage2_5[24],stage2_4[32],stage2_3[32]}
   );
   gpc606_5 gpc567 (
      {stage1_4[39], stage1_4[40], stage1_4[41], stage1_4[42], stage1_4[43], stage1_4[44]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[3],stage2_6[9],stage2_5[25],stage2_4[33]}
   );
   gpc606_5 gpc568 (
      {stage1_4[45], stage1_4[46], stage1_4[47], stage1_4[48], stage1_4[49], stage1_4[50]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[4],stage2_6[10],stage2_5[26],stage2_4[34]}
   );
   gpc606_5 gpc569 (
      {stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[5],stage2_6[11],stage2_5[27],stage2_4[35]}
   );
   gpc615_5 gpc570 (
      {stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61]},
      {stage1_5[18]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[6],stage2_6[12],stage2_5[28],stage2_4[36]}
   );
   gpc615_5 gpc571 (
      {stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65], stage1_4[66]},
      {stage1_5[19]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[7],stage2_6[13],stage2_5[29],stage2_4[37]}
   );
   gpc615_5 gpc572 (
      {stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage1_5[20]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[8],stage2_6[14],stage2_5[30],stage2_4[38]}
   );
   gpc615_5 gpc573 (
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76]},
      {stage1_5[21]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[9],stage2_6[15],stage2_5[31],stage2_4[39]}
   );
   gpc615_5 gpc574 (
      {stage1_4[77], stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81]},
      {stage1_5[22]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[10],stage2_6[16],stage2_5[32],stage2_4[40]}
   );
   gpc615_5 gpc575 (
      {stage1_4[82], stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86]},
      {stage1_5[23]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[11],stage2_6[17],stage2_5[33],stage2_4[41]}
   );
   gpc615_5 gpc576 (
      {stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_5[24]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[12],stage2_6[18],stage2_5[34],stage2_4[42]}
   );
   gpc615_5 gpc577 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96]},
      {stage1_5[25]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[13],stage2_6[19],stage2_5[35],stage2_4[43]}
   );
   gpc615_5 gpc578 (
      {stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage1_5[26]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[14],stage2_6[20],stage2_5[36],stage2_4[44]}
   );
   gpc615_5 gpc579 (
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106]},
      {stage1_5[27]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[15],stage2_6[21],stage2_5[37],stage2_4[45]}
   );
   gpc615_5 gpc580 (
      {stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111]},
      {stage1_5[28]},
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage2_8[13],stage2_7[16],stage2_6[22],stage2_5[38],stage2_4[46]}
   );
   gpc615_5 gpc581 (
      {stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116]},
      {stage1_5[29]},
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage2_8[14],stage2_7[17],stage2_6[23],stage2_5[39],stage2_4[47]}
   );
   gpc615_5 gpc582 (
      {stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_5[30]},
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage2_8[15],stage2_7[18],stage2_6[24],stage2_5[40],stage2_4[48]}
   );
   gpc615_5 gpc583 (
      {stage1_4[122], stage1_4[123], stage1_4[124], stage1_4[125], stage1_4[126]},
      {stage1_5[31]},
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage2_8[16],stage2_7[19],stage2_6[25],stage2_5[41],stage2_4[49]}
   );
   gpc606_5 gpc584 (
      {stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36], stage1_5[37]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[17],stage2_7[20],stage2_6[26],stage2_5[42]}
   );
   gpc606_5 gpc585 (
      {stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41], stage1_5[42], stage1_5[43]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[18],stage2_7[21],stage2_6[27],stage2_5[43]}
   );
   gpc606_5 gpc586 (
      {stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47], stage1_5[48], stage1_5[49]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[19],stage2_7[22],stage2_6[28],stage2_5[44]}
   );
   gpc606_5 gpc587 (
      {stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53], stage1_5[54], stage1_5[55]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[20],stage2_7[23],stage2_6[29],stage2_5[45]}
   );
   gpc606_5 gpc588 (
      {stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59], stage1_5[60], stage1_5[61]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[21],stage2_7[24],stage2_6[30],stage2_5[46]}
   );
   gpc606_5 gpc589 (
      {stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66], stage1_5[67]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[22],stage2_7[25],stage2_6[31],stage2_5[47]}
   );
   gpc606_5 gpc590 (
      {stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71], stage1_5[72], stage1_5[73]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[23],stage2_7[26],stage2_6[32],stage2_5[48]}
   );
   gpc606_5 gpc591 (
      {stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77], stage1_5[78], stage1_5[79]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[24],stage2_7[27],stage2_6[33],stage2_5[49]}
   );
   gpc606_5 gpc592 (
      {stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83], stage1_5[84], stage1_5[85]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[25],stage2_7[28],stage2_6[34],stage2_5[50]}
   );
   gpc606_5 gpc593 (
      {stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89], stage1_5[90], stage1_5[91]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[26],stage2_7[29],stage2_6[35],stage2_5[51]}
   );
   gpc606_5 gpc594 (
      {stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95], stage1_5[96], stage1_5[97]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[27],stage2_7[30],stage2_6[36],stage2_5[52]}
   );
   gpc606_5 gpc595 (
      {stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101], stage1_5[102], stage1_5[103]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[28],stage2_7[31],stage2_6[37],stage2_5[53]}
   );
   gpc615_5 gpc596 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[0]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[12],stage2_8[29],stage2_7[32]}
   );
   gpc615_5 gpc597 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[1]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[1],stage2_9[13],stage2_8[30],stage2_7[33]}
   );
   gpc615_5 gpc598 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[2]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[2],stage2_9[14],stage2_8[31],stage2_7[34]}
   );
   gpc615_5 gpc599 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], stage1_7[91]},
      {stage1_8[3]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[3],stage2_9[15],stage2_8[32],stage2_7[35]}
   );
   gpc606_5 gpc600 (
      {stage1_8[4], stage1_8[5], stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[4],stage2_10[4],stage2_9[16],stage2_8[33]}
   );
   gpc606_5 gpc601 (
      {stage1_8[10], stage1_8[11], stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[5],stage2_10[5],stage2_9[17],stage2_8[34]}
   );
   gpc606_5 gpc602 (
      {stage1_8[16], stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[6],stage2_10[6],stage2_9[18],stage2_8[35]}
   );
   gpc606_5 gpc603 (
      {stage1_8[22], stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[7],stage2_10[7],stage2_9[19],stage2_8[36]}
   );
   gpc606_5 gpc604 (
      {stage1_8[28], stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[8],stage2_10[8],stage2_9[20],stage2_8[37]}
   );
   gpc606_5 gpc605 (
      {stage1_8[34], stage1_8[35], stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[9],stage2_10[9],stage2_9[21],stage2_8[38]}
   );
   gpc606_5 gpc606 (
      {stage1_8[40], stage1_8[41], stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[10],stage2_10[10],stage2_9[22],stage2_8[39]}
   );
   gpc606_5 gpc607 (
      {stage1_8[46], stage1_8[47], stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[11],stage2_10[11],stage2_9[23],stage2_8[40]}
   );
   gpc606_5 gpc608 (
      {stage1_8[52], stage1_8[53], stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[12],stage2_10[12],stage2_9[24],stage2_8[41]}
   );
   gpc606_5 gpc609 (
      {stage1_8[58], stage1_8[59], stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[13],stage2_10[13],stage2_9[25],stage2_8[42]}
   );
   gpc606_5 gpc610 (
      {stage1_8[64], stage1_8[65], stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[14],stage2_10[14],stage2_9[26],stage2_8[43]}
   );
   gpc606_5 gpc611 (
      {stage1_8[70], stage1_8[71], stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[15],stage2_10[15],stage2_9[27],stage2_8[44]}
   );
   gpc606_5 gpc612 (
      {stage1_8[76], stage1_8[77], stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[16],stage2_10[16],stage2_9[28],stage2_8[45]}
   );
   gpc606_5 gpc613 (
      {stage1_8[82], stage1_8[83], stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[17],stage2_10[17],stage2_9[29],stage2_8[46]}
   );
   gpc606_5 gpc614 (
      {stage1_8[88], stage1_8[89], stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[18],stage2_10[18],stage2_9[30],stage2_8[47]}
   );
   gpc606_5 gpc615 (
      {stage1_8[94], stage1_8[95], stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[19],stage2_10[19],stage2_9[31],stage2_8[48]}
   );
   gpc606_5 gpc616 (
      {stage1_8[100], stage1_8[101], stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[20],stage2_10[20],stage2_9[32],stage2_8[49]}
   );
   gpc117_4 gpc617 (
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30]},
      {stage1_10[102]},
      {stage1_11[0]},
      {stage2_12[17],stage2_11[21],stage2_10[21],stage2_9[33]}
   );
   gpc117_4 gpc618 (
      {stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35], stage1_9[36], stage1_9[37]},
      {stage1_10[103]},
      {stage1_11[1]},
      {stage2_12[18],stage2_11[22],stage2_10[22],stage2_9[34]}
   );
   gpc117_4 gpc619 (
      {stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41], stage1_9[42], stage1_9[43], stage1_9[44]},
      {stage1_10[104]},
      {stage1_11[2]},
      {stage2_12[19],stage2_11[23],stage2_10[23],stage2_9[35]}
   );
   gpc117_4 gpc620 (
      {stage1_9[45], stage1_9[46], stage1_9[47], stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51]},
      {stage1_10[105]},
      {stage1_11[3]},
      {stage2_12[20],stage2_11[24],stage2_10[24],stage2_9[36]}
   );
   gpc117_4 gpc621 (
      {stage1_9[52], stage1_9[53], stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58]},
      {stage1_10[106]},
      {stage1_11[4]},
      {stage2_12[21],stage2_11[25],stage2_10[25],stage2_9[37]}
   );
   gpc117_4 gpc622 (
      {stage1_9[59], stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_10[107]},
      {stage1_11[5]},
      {stage2_12[22],stage2_11[26],stage2_10[26],stage2_9[38]}
   );
   gpc117_4 gpc623 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71], stage1_9[72]},
      {stage1_10[108]},
      {stage1_11[6]},
      {stage2_12[23],stage2_11[27],stage2_10[27],stage2_9[39]}
   );
   gpc606_5 gpc624 (
      {stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77], stage1_9[78]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[0],stage2_12[24],stage2_11[28],stage2_10[28],stage2_9[40]}
   );
   gpc606_5 gpc625 (
      {stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83], stage1_9[84]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[1],stage2_12[25],stage2_11[29],stage2_10[29],stage2_9[41]}
   );
   gpc606_5 gpc626 (
      {stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89], stage1_9[90]},
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage2_13[2],stage2_12[26],stage2_11[30],stage2_10[30],stage2_9[42]}
   );
   gpc606_5 gpc627 (
      {stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95], stage1_9[96]},
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29], stage1_11[30]},
      {stage2_13[3],stage2_12[27],stage2_11[31],stage2_10[31],stage2_9[43]}
   );
   gpc606_5 gpc628 (
      {stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101], stage1_9[102]},
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage2_13[4],stage2_12[28],stage2_11[32],stage2_10[32],stage2_9[44]}
   );
   gpc606_5 gpc629 (
      {stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107], stage1_9[108]},
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage2_13[5],stage2_12[29],stage2_11[33],stage2_10[33],stage2_9[45]}
   );
   gpc606_5 gpc630 (
      {stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113], stage1_9[114]},
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage2_13[6],stage2_12[30],stage2_11[34],stage2_10[34],stage2_9[46]}
   );
   gpc615_5 gpc631 (
      {stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage1_11[49]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[7],stage2_12[31],stage2_11[35],stage2_10[35]}
   );
   gpc606_5 gpc632 (
      {stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54], stage1_11[55]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[1],stage2_13[8],stage2_12[32],stage2_11[36]}
   );
   gpc606_5 gpc633 (
      {stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59], stage1_11[60], stage1_11[61]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[2],stage2_13[9],stage2_12[33],stage2_11[37]}
   );
   gpc606_5 gpc634 (
      {stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65], stage1_11[66], stage1_11[67]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[3],stage2_13[10],stage2_12[34],stage2_11[38]}
   );
   gpc606_5 gpc635 (
      {stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72], stage1_11[73]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[4],stage2_13[11],stage2_12[35],stage2_11[39]}
   );
   gpc606_5 gpc636 (
      {stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77], stage1_11[78], stage1_11[79]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[5],stage2_13[12],stage2_12[36],stage2_11[40]}
   );
   gpc615_5 gpc637 (
      {stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83], stage1_11[84]},
      {stage1_12[6]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[6],stage2_13[13],stage2_12[37],stage2_11[41]}
   );
   gpc615_5 gpc638 (
      {stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage1_12[7]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[7],stage2_13[14],stage2_12[38],stage2_11[42]}
   );
   gpc615_5 gpc639 (
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94]},
      {stage1_12[8]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[8],stage2_13[15],stage2_12[39],stage2_11[43]}
   );
   gpc615_5 gpc640 (
      {stage1_11[95], stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99]},
      {stage1_12[9]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[9],stage2_13[16],stage2_12[40],stage2_11[44]}
   );
   gpc615_5 gpc641 (
      {stage1_11[100], stage1_11[101], stage1_11[102], stage1_11[103], stage1_11[104]},
      {stage1_12[10]},
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage2_15[9],stage2_14[10],stage2_13[17],stage2_12[41],stage2_11[45]}
   );
   gpc615_5 gpc642 (
      {stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108], stage1_11[109]},
      {stage1_12[11]},
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage2_15[10],stage2_14[11],stage2_13[18],stage2_12[42],stage2_11[46]}
   );
   gpc615_5 gpc643 (
      {stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[12]},
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage2_15[11],stage2_14[12],stage2_13[19],stage2_12[43],stage2_11[47]}
   );
   gpc606_5 gpc644 (
      {stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[12],stage2_14[13],stage2_13[20],stage2_12[44]}
   );
   gpc606_5 gpc645 (
      {stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[13],stage2_14[14],stage2_13[21],stage2_12[45]}
   );
   gpc606_5 gpc646 (
      {stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[14],stage2_14[15],stage2_13[22],stage2_12[46]}
   );
   gpc606_5 gpc647 (
      {stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35], stage1_12[36]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[15],stage2_14[16],stage2_13[23],stage2_12[47]}
   );
   gpc615_5 gpc648 (
      {stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[72]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[16],stage2_14[17],stage2_13[24],stage2_12[48]}
   );
   gpc615_5 gpc649 (
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46]},
      {stage1_13[73]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[17],stage2_14[18],stage2_13[25],stage2_12[49]}
   );
   gpc615_5 gpc650 (
      {stage1_12[47], stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51]},
      {stage1_13[74]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[18],stage2_14[19],stage2_13[26],stage2_12[50]}
   );
   gpc615_5 gpc651 (
      {stage1_12[52], stage1_12[53], stage1_12[54], stage1_12[55], stage1_12[56]},
      {stage1_13[75]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[19],stage2_14[20],stage2_13[27],stage2_12[51]}
   );
   gpc615_5 gpc652 (
      {stage1_12[57], stage1_12[58], stage1_12[59], stage1_12[60], stage1_12[61]},
      {stage1_13[76]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[20],stage2_14[21],stage2_13[28],stage2_12[52]}
   );
   gpc615_5 gpc653 (
      {stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65], stage1_12[66]},
      {stage1_13[77]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[21],stage2_14[22],stage2_13[29],stage2_12[53]}
   );
   gpc615_5 gpc654 (
      {stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage1_13[78]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[22],stage2_14[23],stage2_13[30],stage2_12[54]}
   );
   gpc615_5 gpc655 (
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76]},
      {stage1_13[79]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[23],stage2_14[24],stage2_13[31],stage2_12[55]}
   );
   gpc615_5 gpc656 (
      {stage1_12[77], stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81]},
      {stage1_13[80]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[24],stage2_14[25],stage2_13[32],stage2_12[56]}
   );
   gpc615_5 gpc657 (
      {stage1_12[82], stage1_12[83], stage1_12[84], stage1_12[85], stage1_12[86]},
      {stage1_13[81]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[25],stage2_14[26],stage2_13[33],stage2_12[57]}
   );
   gpc615_5 gpc658 (
      {stage1_12[87], stage1_12[88], stage1_12[89], stage1_12[90], stage1_12[91]},
      {stage1_13[82]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[26],stage2_14[27],stage2_13[34],stage2_12[58]}
   );
   gpc615_5 gpc659 (
      {stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95], stage1_12[96]},
      {stage1_13[83]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[27],stage2_14[28],stage2_13[35],stage2_12[59]}
   );
   gpc615_5 gpc660 (
      {stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage1_13[84]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[28],stage2_14[29],stage2_13[36],stage2_12[60]}
   );
   gpc606_5 gpc661 (
      {stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89], stage1_13[90]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[17],stage2_15[29],stage2_14[30],stage2_13[37]}
   );
   gpc606_5 gpc662 (
      {stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95], stage1_13[96]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[18],stage2_15[30],stage2_14[31],stage2_13[38]}
   );
   gpc606_5 gpc663 (
      {stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101], stage1_13[102]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[19],stage2_15[31],stage2_14[32],stage2_13[39]}
   );
   gpc606_5 gpc664 (
      {stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107], stage1_13[108]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[20],stage2_15[32],stage2_14[33],stage2_13[40]}
   );
   gpc606_5 gpc665 (
      {stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113], stage1_13[114]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[21],stage2_15[33],stage2_14[34],stage2_13[41]}
   );
   gpc606_5 gpc666 (
      {stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119], stage1_13[120]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[22],stage2_15[34],stage2_14[35],stage2_13[42]}
   );
   gpc606_5 gpc667 (
      {stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125], stage1_13[126]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[23],stage2_15[35],stage2_14[36],stage2_13[43]}
   );
   gpc606_5 gpc668 (
      {stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131], stage1_13[132]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[24],stage2_15[36],stage2_14[37],stage2_13[44]}
   );
   gpc606_5 gpc669 (
      {stage1_14[102], stage1_14[103], stage1_14[104], stage1_14[105], stage1_14[106], stage1_14[107]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[8],stage2_16[25],stage2_15[37],stage2_14[38]}
   );
   gpc606_5 gpc670 (
      {stage1_14[108], stage1_14[109], stage1_14[110], stage1_14[111], stage1_14[112], stage1_14[113]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[9],stage2_16[26],stage2_15[38],stage2_14[39]}
   );
   gpc606_5 gpc671 (
      {stage1_14[114], stage1_14[115], stage1_14[116], stage1_14[117], stage1_14[118], stage1_14[119]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[10],stage2_16[27],stage2_15[39],stage2_14[40]}
   );
   gpc606_5 gpc672 (
      {stage1_14[120], stage1_14[121], stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[11],stage2_16[28],stage2_15[40],stage2_14[41]}
   );
   gpc606_5 gpc673 (
      {stage1_14[126], stage1_14[127], stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[12],stage2_16[29],stage2_15[41],stage2_14[42]}
   );
   gpc606_5 gpc674 (
      {stage1_14[132], stage1_14[133], stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[13],stage2_16[30],stage2_15[42],stage2_14[43]}
   );
   gpc615_5 gpc675 (
      {stage1_14[138], stage1_14[139], stage1_14[140], stage1_14[141], stage1_14[142]},
      {stage1_15[48]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[14],stage2_16[31],stage2_15[43],stage2_14[44]}
   );
   gpc615_5 gpc676 (
      {stage1_14[143], stage1_14[144], stage1_14[145], stage1_14[146], stage1_14[147]},
      {stage1_15[49]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[15],stage2_16[32],stage2_15[44],stage2_14[45]}
   );
   gpc615_5 gpc677 (
      {stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151], stage1_14[152]},
      {stage1_15[50]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[16],stage2_16[33],stage2_15[45],stage2_14[46]}
   );
   gpc615_5 gpc678 (
      {stage1_15[51], stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55]},
      {stage1_16[54]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[9],stage2_17[17],stage2_16[34],stage2_15[46]}
   );
   gpc615_5 gpc679 (
      {stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60]},
      {stage1_16[55]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[10],stage2_17[18],stage2_16[35],stage2_15[47]}
   );
   gpc615_5 gpc680 (
      {stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage1_16[56]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[11],stage2_17[19],stage2_16[36],stage2_15[48]}
   );
   gpc615_5 gpc681 (
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70]},
      {stage1_16[57]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[12],stage2_17[20],stage2_16[37],stage2_15[49]}
   );
   gpc615_5 gpc682 (
      {stage1_15[71], stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75]},
      {stage1_16[58]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[13],stage2_17[21],stage2_16[38],stage2_15[50]}
   );
   gpc1_1 gpc683 (
      {stage1_0[48]},
      {stage2_0[8]}
   );
   gpc1_1 gpc684 (
      {stage1_1[96]},
      {stage2_1[24]}
   );
   gpc1_1 gpc685 (
      {stage1_1[97]},
      {stage2_1[25]}
   );
   gpc1_1 gpc686 (
      {stage1_2[82]},
      {stage2_2[30]}
   );
   gpc1_1 gpc687 (
      {stage1_2[83]},
      {stage2_2[31]}
   );
   gpc1_1 gpc688 (
      {stage1_2[84]},
      {stage2_2[32]}
   );
   gpc1_1 gpc689 (
      {stage1_2[85]},
      {stage2_2[33]}
   );
   gpc1_1 gpc690 (
      {stage1_2[86]},
      {stage2_2[34]}
   );
   gpc1_1 gpc691 (
      {stage1_2[87]},
      {stage2_2[35]}
   );
   gpc1_1 gpc692 (
      {stage1_2[88]},
      {stage2_2[36]}
   );
   gpc1_1 gpc693 (
      {stage1_2[89]},
      {stage2_2[37]}
   );
   gpc1_1 gpc694 (
      {stage1_2[90]},
      {stage2_2[38]}
   );
   gpc1_1 gpc695 (
      {stage1_2[91]},
      {stage2_2[39]}
   );
   gpc1_1 gpc696 (
      {stage1_2[92]},
      {stage2_2[40]}
   );
   gpc1_1 gpc697 (
      {stage1_2[93]},
      {stage2_2[41]}
   );
   gpc1_1 gpc698 (
      {stage1_2[94]},
      {stage2_2[42]}
   );
   gpc1_1 gpc699 (
      {stage1_2[95]},
      {stage2_2[43]}
   );
   gpc1_1 gpc700 (
      {stage1_2[96]},
      {stage2_2[44]}
   );
   gpc1_1 gpc701 (
      {stage1_2[97]},
      {stage2_2[45]}
   );
   gpc1_1 gpc702 (
      {stage1_3[113]},
      {stage2_3[33]}
   );
   gpc1_1 gpc703 (
      {stage1_5[104]},
      {stage2_5[54]}
   );
   gpc1_1 gpc704 (
      {stage1_6[102]},
      {stage2_6[38]}
   );
   gpc1_1 gpc705 (
      {stage1_6[103]},
      {stage2_6[39]}
   );
   gpc1_1 gpc706 (
      {stage1_7[92]},
      {stage2_7[36]}
   );
   gpc1_1 gpc707 (
      {stage1_7[93]},
      {stage2_7[37]}
   );
   gpc1_1 gpc708 (
      {stage1_7[94]},
      {stage2_7[38]}
   );
   gpc1_1 gpc709 (
      {stage1_7[95]},
      {stage2_7[39]}
   );
   gpc1_1 gpc710 (
      {stage1_7[96]},
      {stage2_7[40]}
   );
   gpc1_1 gpc711 (
      {stage1_7[97]},
      {stage2_7[41]}
   );
   gpc1_1 gpc712 (
      {stage1_7[98]},
      {stage2_7[42]}
   );
   gpc1_1 gpc713 (
      {stage1_7[99]},
      {stage2_7[43]}
   );
   gpc1_1 gpc714 (
      {stage1_7[100]},
      {stage2_7[44]}
   );
   gpc1_1 gpc715 (
      {stage1_7[101]},
      {stage2_7[45]}
   );
   gpc1_1 gpc716 (
      {stage1_7[102]},
      {stage2_7[46]}
   );
   gpc1_1 gpc717 (
      {stage1_7[103]},
      {stage2_7[47]}
   );
   gpc1_1 gpc718 (
      {stage1_7[104]},
      {stage2_7[48]}
   );
   gpc1_1 gpc719 (
      {stage1_7[105]},
      {stage2_7[49]}
   );
   gpc1_1 gpc720 (
      {stage1_7[106]},
      {stage2_7[50]}
   );
   gpc1_1 gpc721 (
      {stage1_7[107]},
      {stage2_7[51]}
   );
   gpc1_1 gpc722 (
      {stage1_7[108]},
      {stage2_7[52]}
   );
   gpc1_1 gpc723 (
      {stage1_7[109]},
      {stage2_7[53]}
   );
   gpc1_1 gpc724 (
      {stage1_7[110]},
      {stage2_7[54]}
   );
   gpc1_1 gpc725 (
      {stage1_7[111]},
      {stage2_7[55]}
   );
   gpc1_1 gpc726 (
      {stage1_7[112]},
      {stage2_7[56]}
   );
   gpc1_1 gpc727 (
      {stage1_7[113]},
      {stage2_7[57]}
   );
   gpc1_1 gpc728 (
      {stage1_7[114]},
      {stage2_7[58]}
   );
   gpc1_1 gpc729 (
      {stage1_9[115]},
      {stage2_9[47]}
   );
   gpc1_1 gpc730 (
      {stage1_14[153]},
      {stage2_14[47]}
   );
   gpc1_1 gpc731 (
      {stage1_14[154]},
      {stage2_14[48]}
   );
   gpc1_1 gpc732 (
      {stage1_14[155]},
      {stage2_14[49]}
   );
   gpc1_1 gpc733 (
      {stage1_14[156]},
      {stage2_14[50]}
   );
   gpc1_1 gpc734 (
      {stage1_16[59]},
      {stage2_16[39]}
   );
   gpc1_1 gpc735 (
      {stage1_16[60]},
      {stage2_16[40]}
   );
   gpc1_1 gpc736 (
      {stage1_16[61]},
      {stage2_16[41]}
   );
   gpc1_1 gpc737 (
      {stage1_16[62]},
      {stage2_16[42]}
   );
   gpc1_1 gpc738 (
      {stage1_16[63]},
      {stage2_16[43]}
   );
   gpc1_1 gpc739 (
      {stage1_16[64]},
      {stage2_16[44]}
   );
   gpc1_1 gpc740 (
      {stage1_16[65]},
      {stage2_16[45]}
   );
   gpc1_1 gpc741 (
      {stage1_16[66]},
      {stage2_16[46]}
   );
   gpc1_1 gpc742 (
      {stage1_16[67]},
      {stage2_16[47]}
   );
   gpc1_1 gpc743 (
      {stage1_17[30]},
      {stage2_17[22]}
   );
   gpc1_1 gpc744 (
      {stage1_17[31]},
      {stage2_17[23]}
   );
   gpc1_1 gpc745 (
      {stage1_17[32]},
      {stage2_17[24]}
   );
   gpc1_1 gpc746 (
      {stage1_17[33]},
      {stage2_17[25]}
   );
   gpc1_1 gpc747 (
      {stage1_17[34]},
      {stage2_17[26]}
   );
   gpc1_1 gpc748 (
      {stage1_17[35]},
      {stage2_17[27]}
   );
   gpc1_1 gpc749 (
      {stage1_17[36]},
      {stage2_17[28]}
   );
   gpc1_1 gpc750 (
      {stage1_17[37]},
      {stage2_17[29]}
   );
   gpc1_1 gpc751 (
      {stage1_17[38]},
      {stage2_17[30]}
   );
   gpc1_1 gpc752 (
      {stage1_17[39]},
      {stage2_17[31]}
   );
   gpc1_1 gpc753 (
      {stage1_17[40]},
      {stage2_17[32]}
   );
   gpc1_1 gpc754 (
      {stage1_17[41]},
      {stage2_17[33]}
   );
   gpc1163_5 gpc755 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc756 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6]},
      {stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc606_5 gpc757 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12]},
      {stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc758 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage3_5[2],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc759 (
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[3],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc606_5 gpc760 (
      {stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11], stage2_2[12]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[4],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc606_5 gpc761 (
      {stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17], stage2_2[18]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[5],stage3_4[6],stage3_3[6],stage3_2[6]}
   );
   gpc615_5 gpc762 (
      {stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage2_3[19]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[6],stage3_4[7],stage3_3[7],stage3_2[7]}
   );
   gpc615_5 gpc763 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[20]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[7],stage3_4[8],stage3_3[8],stage3_2[8]}
   );
   gpc615_5 gpc764 (
      {stage2_2[29], stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33]},
      {stage2_3[21]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[8],stage3_4[9],stage3_3[9],stage3_2[9]}
   );
   gpc615_5 gpc765 (
      {stage2_2[34], stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38]},
      {stage2_3[22]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[9],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc615_5 gpc766 (
      {stage2_2[39], stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43]},
      {stage2_3[23]},
      {stage2_4[42], stage2_4[43], stage2_4[44], stage2_4[45], stage2_4[46], stage2_4[47]},
      {stage3_6[7],stage3_5[10],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc767 (
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28]},
      {stage2_4[48]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[8],stage3_5[11],stage3_4[12],stage3_3[12]}
   );
   gpc615_5 gpc768 (
      {stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage2_4[49]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[9],stage3_5[12],stage3_4[13],stage3_3[13]}
   );
   gpc7_3 gpc769 (
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17], stage2_5[18]},
      {stage3_7[2],stage3_6[10],stage3_5[13]}
   );
   gpc207_4 gpc770 (
      {stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23], stage2_5[24], stage2_5[25]},
      {stage2_7[0], stage2_7[1]},
      {stage3_8[0],stage3_7[3],stage3_6[11],stage3_5[14]}
   );
   gpc606_5 gpc771 (
      {stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29], stage2_5[30], stage2_5[31]},
      {stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6], stage2_7[7]},
      {stage3_9[0],stage3_8[1],stage3_7[4],stage3_6[12],stage3_5[15]}
   );
   gpc606_5 gpc772 (
      {stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35], stage2_5[36], stage2_5[37]},
      {stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11], stage2_7[12], stage2_7[13]},
      {stage3_9[1],stage3_8[2],stage3_7[5],stage3_6[13],stage3_5[16]}
   );
   gpc606_5 gpc773 (
      {stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41], stage2_5[42], stage2_5[43]},
      {stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18], stage2_7[19]},
      {stage3_9[2],stage3_8[3],stage3_7[6],stage3_6[14],stage3_5[17]}
   );
   gpc606_5 gpc774 (
      {stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47], stage2_5[48], stage2_5[49]},
      {stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25]},
      {stage3_9[3],stage3_8[4],stage3_7[7],stage3_6[15],stage3_5[18]}
   );
   gpc606_5 gpc775 (
      {stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53], stage2_5[54], 1'b0},
      {stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage3_9[4],stage3_8[5],stage3_7[8],stage3_6[16],stage3_5[19]}
   );
   gpc615_5 gpc776 (
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4]},
      {stage2_7[32]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[5],stage3_8[6],stage3_7[9],stage3_6[17]}
   );
   gpc615_5 gpc777 (
      {stage2_6[5], stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9]},
      {stage2_7[33]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[6],stage3_8[7],stage3_7[10],stage3_6[18]}
   );
   gpc615_5 gpc778 (
      {stage2_6[10], stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14]},
      {stage2_7[34]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[7],stage3_8[8],stage3_7[11],stage3_6[19]}
   );
   gpc615_5 gpc779 (
      {stage2_6[15], stage2_6[16], stage2_6[17], stage2_6[18], stage2_6[19]},
      {stage2_7[35]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[8],stage3_8[9],stage3_7[12],stage3_6[20]}
   );
   gpc615_5 gpc780 (
      {stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24]},
      {stage2_7[36]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[9],stage3_8[10],stage3_7[13],stage3_6[21]}
   );
   gpc615_5 gpc781 (
      {stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage2_7[37]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[10],stage3_8[11],stage3_7[14],stage3_6[22]}
   );
   gpc615_5 gpc782 (
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34]},
      {stage2_7[38]},
      {stage2_8[36], stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41]},
      {stage3_10[6],stage3_9[11],stage3_8[12],stage3_7[15],stage3_6[23]}
   );
   gpc615_5 gpc783 (
      {stage2_6[35], stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39]},
      {stage2_7[39]},
      {stage2_8[42], stage2_8[43], stage2_8[44], stage2_8[45], stage2_8[46], stage2_8[47]},
      {stage3_10[7],stage3_9[12],stage3_8[13],stage3_7[16],stage3_6[24]}
   );
   gpc606_5 gpc784 (
      {stage2_7[40], stage2_7[41], stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[8],stage3_9[13],stage3_8[14],stage3_7[17]}
   );
   gpc615_5 gpc785 (
      {stage2_7[46], stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50]},
      {stage2_8[48]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[9],stage3_9[14],stage3_8[15],stage3_7[18]}
   );
   gpc615_5 gpc786 (
      {stage2_7[51], stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55]},
      {stage2_8[49]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[10],stage3_9[15],stage3_8[16],stage3_7[19]}
   );
   gpc606_5 gpc787 (
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[0],stage3_11[3],stage3_10[11],stage3_9[16]}
   );
   gpc606_5 gpc788 (
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[1],stage3_11[4],stage3_10[12],stage3_9[17]}
   );
   gpc606_5 gpc789 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[2],stage3_11[5],stage3_10[13],stage3_9[18]}
   );
   gpc606_5 gpc790 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[3],stage3_11[6],stage3_10[14],stage3_9[19]}
   );
   gpc606_5 gpc791 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], stage2_11[29]},
      {stage3_13[4],stage3_12[4],stage3_11[7],stage3_10[15],stage3_9[20]}
   );
   gpc606_5 gpc792 (
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[5],stage3_12[5],stage3_11[8],stage3_10[16]}
   );
   gpc615_5 gpc793 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10]},
      {stage2_11[30]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[6],stage3_12[6],stage3_11[9],stage3_10[17]}
   );
   gpc615_5 gpc794 (
      {stage2_10[11], stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15]},
      {stage2_11[31]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[7],stage3_12[7],stage3_11[10],stage3_10[18]}
   );
   gpc615_5 gpc795 (
      {stage2_10[16], stage2_10[17], stage2_10[18], stage2_10[19], stage2_10[20]},
      {stage2_11[32]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[8],stage3_12[8],stage3_11[11],stage3_10[19]}
   );
   gpc615_5 gpc796 (
      {stage2_10[21], stage2_10[22], stage2_10[23], stage2_10[24], stage2_10[25]},
      {stage2_11[33]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[9],stage3_12[9],stage3_11[12],stage3_10[20]}
   );
   gpc615_5 gpc797 (
      {stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29], stage2_10[30]},
      {stage2_11[34]},
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage3_14[5],stage3_13[10],stage3_12[10],stage3_11[13],stage3_10[21]}
   );
   gpc615_5 gpc798 (
      {stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage2_11[35]},
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage3_14[6],stage3_13[11],stage3_12[11],stage3_11[14],stage3_10[22]}
   );
   gpc606_5 gpc799 (
      {stage2_11[36], stage2_11[37], stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[7],stage3_13[12],stage3_12[12],stage3_11[15]}
   );
   gpc606_5 gpc800 (
      {stage2_11[42], stage2_11[43], stage2_11[44], stage2_11[45], stage2_11[46], stage2_11[47]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[8],stage3_13[13],stage3_12[13],stage3_11[16]}
   );
   gpc606_5 gpc801 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[2],stage3_14[9],stage3_13[14],stage3_12[14]}
   );
   gpc606_5 gpc802 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[3],stage3_14[10],stage3_13[15],stage3_12[15]}
   );
   gpc117_4 gpc803 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17], stage2_13[18]},
      {stage2_14[12]},
      {stage2_15[0]},
      {stage3_16[2],stage3_15[4],stage3_14[11],stage3_13[16]}
   );
   gpc117_4 gpc804 (
      {stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23], stage2_13[24], stage2_13[25]},
      {stage2_14[13]},
      {stage2_15[1]},
      {stage3_16[3],stage3_15[5],stage3_14[12],stage3_13[17]}
   );
   gpc117_4 gpc805 (
      {stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29], stage2_13[30], stage2_13[31], stage2_13[32]},
      {stage2_14[14]},
      {stage2_15[2]},
      {stage3_16[4],stage3_15[6],stage3_14[13],stage3_13[18]}
   );
   gpc606_5 gpc806 (
      {stage2_13[33], stage2_13[34], stage2_13[35], stage2_13[36], stage2_13[37], stage2_13[38]},
      {stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8]},
      {stage3_17[0],stage3_16[5],stage3_15[7],stage3_14[14],stage3_13[19]}
   );
   gpc606_5 gpc807 (
      {stage2_13[39], stage2_13[40], stage2_13[41], stage2_13[42], stage2_13[43], stage2_13[44]},
      {stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage3_17[1],stage3_16[6],stage3_15[8],stage3_14[15],stage3_13[20]}
   );
   gpc117_4 gpc808 (
      {stage2_14[15], stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21]},
      {stage2_15[15]},
      {stage2_16[0]},
      {stage3_17[2],stage3_16[7],stage3_15[9],stage3_14[16]}
   );
   gpc606_5 gpc809 (
      {stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27]},
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage3_18[0],stage3_17[3],stage3_16[8],stage3_15[10],stage3_14[17]}
   );
   gpc606_5 gpc810 (
      {stage2_14[28], stage2_14[29], stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33]},
      {stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11], stage2_16[12]},
      {stage3_18[1],stage3_17[4],stage3_16[9],stage3_15[11],stage3_14[18]}
   );
   gpc606_5 gpc811 (
      {stage2_14[34], stage2_14[35], stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39]},
      {stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17], stage2_16[18]},
      {stage3_18[2],stage3_17[5],stage3_16[10],stage3_15[12],stage3_14[19]}
   );
   gpc606_5 gpc812 (
      {stage2_14[40], stage2_14[41], stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45]},
      {stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23], stage2_16[24]},
      {stage3_18[3],stage3_17[6],stage3_16[11],stage3_15[13],stage3_14[20]}
   );
   gpc606_5 gpc813 (
      {stage2_14[46], stage2_14[47], stage2_14[48], stage2_14[49], stage2_14[50], 1'b0},
      {stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29], stage2_16[30]},
      {stage3_18[4],stage3_17[7],stage3_16[12],stage3_15[14],stage3_14[21]}
   );
   gpc606_5 gpc814 (
      {stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[5],stage3_17[8],stage3_16[13],stage3_15[15]}
   );
   gpc606_5 gpc815 (
      {stage2_15[22], stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[6],stage3_17[9],stage3_16[14],stage3_15[16]}
   );
   gpc606_5 gpc816 (
      {stage2_15[28], stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[7],stage3_17[10],stage3_16[15],stage3_15[17]}
   );
   gpc606_5 gpc817 (
      {stage2_15[34], stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[8],stage3_17[11],stage3_16[16],stage3_15[18]}
   );
   gpc606_5 gpc818 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44], stage2_15[45]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[9],stage3_17[12],stage3_16[17],stage3_15[19]}
   );
   gpc606_5 gpc819 (
      {stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35], stage2_16[36]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[5],stage3_18[10],stage3_17[13],stage3_16[18]}
   );
   gpc606_5 gpc820 (
      {stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41], stage2_16[42]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[6],stage3_18[11],stage3_17[14],stage3_16[19]}
   );
   gpc1_1 gpc821 (
      {stage2_0[3]},
      {stage3_0[1]}
   );
   gpc1_1 gpc822 (
      {stage2_0[4]},
      {stage3_0[2]}
   );
   gpc1_1 gpc823 (
      {stage2_0[5]},
      {stage3_0[3]}
   );
   gpc1_1 gpc824 (
      {stage2_0[6]},
      {stage3_0[4]}
   );
   gpc1_1 gpc825 (
      {stage2_0[7]},
      {stage3_0[5]}
   );
   gpc1_1 gpc826 (
      {stage2_0[8]},
      {stage3_0[6]}
   );
   gpc1_1 gpc827 (
      {stage2_1[24]},
      {stage3_1[4]}
   );
   gpc1_1 gpc828 (
      {stage2_1[25]},
      {stage3_1[5]}
   );
   gpc1_1 gpc829 (
      {stage2_2[44]},
      {stage3_2[12]}
   );
   gpc1_1 gpc830 (
      {stage2_2[45]},
      {stage3_2[13]}
   );
   gpc1_1 gpc831 (
      {stage2_7[56]},
      {stage3_7[20]}
   );
   gpc1_1 gpc832 (
      {stage2_7[57]},
      {stage3_7[21]}
   );
   gpc1_1 gpc833 (
      {stage2_7[58]},
      {stage3_7[22]}
   );
   gpc1_1 gpc834 (
      {stage2_12[54]},
      {stage3_12[16]}
   );
   gpc1_1 gpc835 (
      {stage2_12[55]},
      {stage3_12[17]}
   );
   gpc1_1 gpc836 (
      {stage2_12[56]},
      {stage3_12[18]}
   );
   gpc1_1 gpc837 (
      {stage2_12[57]},
      {stage3_12[19]}
   );
   gpc1_1 gpc838 (
      {stage2_12[58]},
      {stage3_12[20]}
   );
   gpc1_1 gpc839 (
      {stage2_12[59]},
      {stage3_12[21]}
   );
   gpc1_1 gpc840 (
      {stage2_12[60]},
      {stage3_12[22]}
   );
   gpc1_1 gpc841 (
      {stage2_15[46]},
      {stage3_15[20]}
   );
   gpc1_1 gpc842 (
      {stage2_15[47]},
      {stage3_15[21]}
   );
   gpc1_1 gpc843 (
      {stage2_15[48]},
      {stage3_15[22]}
   );
   gpc1_1 gpc844 (
      {stage2_15[49]},
      {stage3_15[23]}
   );
   gpc1_1 gpc845 (
      {stage2_15[50]},
      {stage3_15[24]}
   );
   gpc1_1 gpc846 (
      {stage2_16[43]},
      {stage3_16[20]}
   );
   gpc1_1 gpc847 (
      {stage2_16[44]},
      {stage3_16[21]}
   );
   gpc1_1 gpc848 (
      {stage2_16[45]},
      {stage3_16[22]}
   );
   gpc1_1 gpc849 (
      {stage2_16[46]},
      {stage3_16[23]}
   );
   gpc1_1 gpc850 (
      {stage2_16[47]},
      {stage3_16[24]}
   );
   gpc1_1 gpc851 (
      {stage2_17[30]},
      {stage3_17[15]}
   );
   gpc1_1 gpc852 (
      {stage2_17[31]},
      {stage3_17[16]}
   );
   gpc1_1 gpc853 (
      {stage2_17[32]},
      {stage3_17[17]}
   );
   gpc1_1 gpc854 (
      {stage2_17[33]},
      {stage3_17[18]}
   );
   gpc1_1 gpc855 (
      {stage2_18[12]},
      {stage3_18[12]}
   );
   gpc1_1 gpc856 (
      {stage2_18[13]},
      {stage3_18[13]}
   );
   gpc1_1 gpc857 (
      {stage2_19[0]},
      {stage3_19[7]}
   );
   gpc1_1 gpc858 (
      {stage2_19[1]},
      {stage3_19[8]}
   );
   gpc1_1 gpc859 (
      {stage2_19[2]},
      {stage3_19[9]}
   );
   gpc1_1 gpc860 (
      {stage2_19[3]},
      {stage3_19[10]}
   );
   gpc1_1 gpc861 (
      {stage2_19[4]},
      {stage3_19[11]}
   );
   gpc606_5 gpc862 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc606_5 gpc863 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc864 (
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10]},
      {stage3_4[0]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc606_5 gpc865 (
      {stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5], stage3_4[6]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[1],stage4_6[1],stage4_5[2],stage4_4[3]}
   );
   gpc606_5 gpc866 (
      {stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11], stage3_4[12]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[2],stage4_6[2],stage4_5[3],stage4_4[4]}
   );
   gpc7_3 gpc867 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11], stage3_5[12]},
      {stage4_7[3],stage4_6[3],stage4_5[4]}
   );
   gpc7_3 gpc868 (
      {stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17], stage3_5[18], stage3_5[19]},
      {stage4_7[4],stage4_6[4],stage4_5[5]}
   );
   gpc207_4 gpc869 (
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17], stage3_6[18]},
      {stage3_8[0], stage3_8[1]},
      {stage4_9[0],stage4_8[2],stage4_7[5],stage4_6[5]}
   );
   gpc615_5 gpc870 (
      {stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_7[0]},
      {stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5], stage3_8[6], stage3_8[7]},
      {stage4_10[0],stage4_9[1],stage4_8[3],stage4_7[6],stage4_6[6]}
   );
   gpc615_5 gpc871 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[8]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[2],stage4_8[4],stage4_7[7]}
   );
   gpc615_5 gpc872 (
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10]},
      {stage3_8[9]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[3],stage4_8[5],stage4_7[8]}
   );
   gpc615_5 gpc873 (
      {stage3_7[11], stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15]},
      {stage3_8[10]},
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage4_11[2],stage4_10[3],stage4_9[4],stage4_8[6],stage4_7[9]}
   );
   gpc606_5 gpc874 (
      {stage3_8[11], stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[3],stage4_10[4],stage4_9[5],stage4_8[7]}
   );
   gpc615_5 gpc875 (
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10]},
      {stage3_11[0]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[0],stage4_12[1],stage4_11[4],stage4_10[5]}
   );
   gpc615_5 gpc876 (
      {stage3_10[11], stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15]},
      {stage3_11[1]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[1],stage4_12[2],stage4_11[5],stage4_10[6]}
   );
   gpc615_5 gpc877 (
      {stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19], stage3_10[20]},
      {stage3_11[2]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[2],stage4_12[3],stage4_11[6],stage4_10[7]}
   );
   gpc207_4 gpc878 (
      {stage3_11[3], stage3_11[4], stage3_11[5], stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[3],stage4_13[3],stage4_12[4],stage4_11[7]}
   );
   gpc606_5 gpc879 (
      {stage3_11[10], stage3_11[11], stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15]},
      {stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7]},
      {stage4_15[0],stage4_14[4],stage4_13[4],stage4_12[5],stage4_11[8]}
   );
   gpc615_5 gpc880 (
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22]},
      {stage3_13[8]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[5],stage4_13[5],stage4_12[6]}
   );
   gpc606_5 gpc881 (
      {stage3_13[9], stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[6],stage4_13[6]}
   );
   gpc606_5 gpc882 (
      {stage3_13[15], stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[2],stage4_15[3],stage4_14[7],stage4_13[7]}
   );
   gpc606_5 gpc883 (
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[2],stage4_16[3],stage4_15[4],stage4_14[8]}
   );
   gpc615_5 gpc884 (
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[12]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[3],stage4_16[4],stage4_15[5],stage4_14[9]}
   );
   gpc615_5 gpc885 (
      {stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21]},
      {stage3_15[13]},
      {stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15], stage3_16[16], stage3_16[17]},
      {stage4_18[2],stage4_17[4],stage4_16[5],stage4_15[6],stage4_14[10]}
   );
   gpc606_5 gpc886 (
      {stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[3],stage4_17[5],stage4_16[6],stage4_15[7]}
   );
   gpc615_5 gpc887 (
      {stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24]},
      {stage3_16[18]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[4],stage4_17[6],stage4_16[7],stage4_15[8]}
   );
   gpc606_5 gpc888 (
      {stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22], stage3_16[23], stage3_16[24]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[2],stage4_18[5],stage4_17[7],stage4_16[8]}
   );
   gpc606_5 gpc889 (
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[1],stage4_19[3],stage4_18[6],stage4_17[8]}
   );
   gpc117_4 gpc890 (
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11], stage3_18[12]},
      {stage3_19[6]},
      {stage3_20[0]},
      {stage4_21[1],stage4_20[2],stage4_19[4],stage4_18[7]}
   );
   gpc1_1 gpc891 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc892 (
      {stage3_2[6]},
      {stage4_2[2]}
   );
   gpc1_1 gpc893 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc894 (
      {stage3_2[8]},
      {stage4_2[4]}
   );
   gpc1_1 gpc895 (
      {stage3_2[9]},
      {stage4_2[5]}
   );
   gpc1_1 gpc896 (
      {stage3_2[10]},
      {stage4_2[6]}
   );
   gpc1_1 gpc897 (
      {stage3_2[11]},
      {stage4_2[7]}
   );
   gpc1_1 gpc898 (
      {stage3_2[12]},
      {stage4_2[8]}
   );
   gpc1_1 gpc899 (
      {stage3_2[13]},
      {stage4_2[9]}
   );
   gpc1_1 gpc900 (
      {stage3_3[11]},
      {stage4_3[3]}
   );
   gpc1_1 gpc901 (
      {stage3_3[12]},
      {stage4_3[4]}
   );
   gpc1_1 gpc902 (
      {stage3_3[13]},
      {stage4_3[5]}
   );
   gpc1_1 gpc903 (
      {stage3_4[13]},
      {stage4_4[5]}
   );
   gpc1_1 gpc904 (
      {stage3_6[24]},
      {stage4_6[7]}
   );
   gpc1_1 gpc905 (
      {stage3_7[16]},
      {stage4_7[10]}
   );
   gpc1_1 gpc906 (
      {stage3_7[17]},
      {stage4_7[11]}
   );
   gpc1_1 gpc907 (
      {stage3_7[18]},
      {stage4_7[12]}
   );
   gpc1_1 gpc908 (
      {stage3_7[19]},
      {stage4_7[13]}
   );
   gpc1_1 gpc909 (
      {stage3_7[20]},
      {stage4_7[14]}
   );
   gpc1_1 gpc910 (
      {stage3_7[21]},
      {stage4_7[15]}
   );
   gpc1_1 gpc911 (
      {stage3_7[22]},
      {stage4_7[16]}
   );
   gpc1_1 gpc912 (
      {stage3_9[18]},
      {stage4_9[6]}
   );
   gpc1_1 gpc913 (
      {stage3_9[19]},
      {stage4_9[7]}
   );
   gpc1_1 gpc914 (
      {stage3_9[20]},
      {stage4_9[8]}
   );
   gpc1_1 gpc915 (
      {stage3_10[21]},
      {stage4_10[8]}
   );
   gpc1_1 gpc916 (
      {stage3_10[22]},
      {stage4_10[9]}
   );
   gpc1_1 gpc917 (
      {stage3_11[16]},
      {stage4_11[9]}
   );
   gpc1_1 gpc918 (
      {stage3_17[18]},
      {stage4_17[9]}
   );
   gpc1_1 gpc919 (
      {stage3_18[13]},
      {stage4_18[8]}
   );
   gpc1_1 gpc920 (
      {stage3_19[7]},
      {stage4_19[5]}
   );
   gpc1_1 gpc921 (
      {stage3_19[8]},
      {stage4_19[6]}
   );
   gpc1_1 gpc922 (
      {stage3_19[9]},
      {stage4_19[7]}
   );
   gpc1_1 gpc923 (
      {stage3_19[10]},
      {stage4_19[8]}
   );
   gpc1_1 gpc924 (
      {stage3_19[11]},
      {stage4_19[9]}
   );
   gpc1_1 gpc925 (
      {stage3_20[1]},
      {stage4_20[3]}
   );
   gpc15_3 gpc926 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[0]},
      {stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc615_5 gpc927 (
      {stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage4_4[0]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[1],stage5_3[1]}
   );
   gpc1163_5 gpc928 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage4_8[0]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[1],stage5_6[1]}
   );
   gpc1163_5 gpc929 (
      {stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage4_8[1]},
      {stage4_9[1]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[2],stage5_6[2]}
   );
   gpc615_5 gpc930 (
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16]},
      {stage4_8[2]},
      {stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5], stage4_9[6], stage4_9[7]},
      {stage5_11[0],stage5_10[2],stage5_9[2],stage5_8[2],stage5_7[3]}
   );
   gpc615_5 gpc931 (
      {stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6], stage4_8[7]},
      {stage4_9[8]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[1],stage5_10[3],stage5_9[3],stage5_8[3]}
   );
   gpc1163_5 gpc932 (
      {stage4_10[6], stage4_10[7], stage4_10[8]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage4_12[0]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[0],stage5_12[1],stage5_11[2],stage5_10[4]}
   );
   gpc1163_5 gpc933 (
      {stage4_11[6], stage4_11[7], stage4_11[8]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6]},
      {stage4_13[1]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[1],stage5_13[1],stage5_12[2],stage5_11[3]}
   );
   gpc135_4 gpc934 (
      {stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6]},
      {stage4_14[1], stage4_14[2], stage4_14[3]},
      {stage4_15[0]},
      {stage5_16[0],stage5_15[1],stage5_14[2],stage5_13[2]}
   );
   gpc7_3 gpc935 (
      {stage4_14[4], stage4_14[5], stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage5_16[1],stage5_15[2],stage5_14[3]}
   );
   gpc606_5 gpc936 (
      {stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[0],stage5_17[0],stage5_16[2],stage5_15[3]}
   );
   gpc2135_5 gpc937 (
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4]},
      {stage4_17[6], stage4_17[7], stage4_17[8]},
      {stage4_18[0]},
      {stage4_19[0], stage4_19[1]},
      {stage5_20[0],stage5_19[1],stage5_18[1],stage5_17[1],stage5_16[3]}
   );
   gpc615_5 gpc938 (
      {stage4_16[5], stage4_16[6], stage4_16[7], stage4_16[8], 1'b0},
      {stage4_17[9]},
      {stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage5_20[1],stage5_19[2],stage5_18[2],stage5_17[2],stage5_16[4]}
   );
   gpc1163_5 gpc939 (
      {stage4_18[7], stage4_18[8], 1'b0},
      {stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5], stage4_19[6], stage4_19[7]},
      {stage4_20[0]},
      {stage4_21[0]},
      {stage5_22[0],stage5_21[0],stage5_20[2],stage5_19[3],stage5_18[3]}
   );
   gpc1_1 gpc940 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc941 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc942 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc943 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc944 (
      {stage4_2[5]},
      {stage5_2[1]}
   );
   gpc1_1 gpc945 (
      {stage4_2[6]},
      {stage5_2[2]}
   );
   gpc1_1 gpc946 (
      {stage4_2[7]},
      {stage5_2[3]}
   );
   gpc1_1 gpc947 (
      {stage4_2[8]},
      {stage5_2[4]}
   );
   gpc1_1 gpc948 (
      {stage4_2[9]},
      {stage5_2[5]}
   );
   gpc1_1 gpc949 (
      {stage4_4[1]},
      {stage5_4[2]}
   );
   gpc1_1 gpc950 (
      {stage4_4[2]},
      {stage5_4[3]}
   );
   gpc1_1 gpc951 (
      {stage4_4[3]},
      {stage5_4[4]}
   );
   gpc1_1 gpc952 (
      {stage4_4[4]},
      {stage5_4[5]}
   );
   gpc1_1 gpc953 (
      {stage4_4[5]},
      {stage5_4[6]}
   );
   gpc1_1 gpc954 (
      {stage4_6[6]},
      {stage5_6[3]}
   );
   gpc1_1 gpc955 (
      {stage4_6[7]},
      {stage5_6[4]}
   );
   gpc1_1 gpc956 (
      {stage4_10[9]},
      {stage5_10[5]}
   );
   gpc1_1 gpc957 (
      {stage4_11[9]},
      {stage5_11[4]}
   );
   gpc1_1 gpc958 (
      {stage4_13[7]},
      {stage5_13[3]}
   );
   gpc1_1 gpc959 (
      {stage4_15[7]},
      {stage5_15[4]}
   );
   gpc1_1 gpc960 (
      {stage4_15[8]},
      {stage5_15[5]}
   );
   gpc1_1 gpc961 (
      {stage4_19[8]},
      {stage5_19[4]}
   );
   gpc1_1 gpc962 (
      {stage4_19[9]},
      {stage5_19[5]}
   );
   gpc1_1 gpc963 (
      {stage4_20[1]},
      {stage5_20[3]}
   );
   gpc1_1 gpc964 (
      {stage4_20[2]},
      {stage5_20[4]}
   );
   gpc1_1 gpc965 (
      {stage4_20[3]},
      {stage5_20[5]}
   );
   gpc1_1 gpc966 (
      {stage4_21[1]},
      {stage5_21[1]}
   );
   gpc615_5 gpc967 (
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4]},
      {stage5_3[0]},
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5]},
      {stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc135_4 gpc968 (
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4]},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[0],stage6_6[1]}
   );
   gpc1343_5 gpc969 (
      {stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[1]}
   );
   gpc1343_5 gpc970 (
      {stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4]},
      {stage5_12[0], stage5_12[1], stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1],stage6_10[1]}
   );
   gpc1343_5 gpc971 (
      {stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[0], stage5_14[1], stage5_14[2], stage5_14[3]},
      {stage5_15[0], stage5_15[1], stage5_15[2]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc1343_5 gpc972 (
      {stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4]},
      {stage5_17[0], stage5_17[1], stage5_17[2]},
      {stage5_18[0]},
      {stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1]}
   );
   gpc1163_5 gpc973 (
      {stage5_18[1], stage5_18[2], stage5_18[3]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage5_20[0]},
      {stage5_21[0]},
      {stage6_22[0],stage6_21[0],stage6_20[0],stage6_19[1],stage6_18[1]}
   );
   gpc135_4 gpc974 (
      {stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage5_21[1], 1'b0, 1'b0},
      {stage5_22[0]},
      {stage6_23[0],stage6_22[1],stage6_21[1],stage6_20[1]}
   );
   gpc1_1 gpc975 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc976 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc977 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc978 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc979 (
      {stage5_2[5]},
      {stage6_2[1]}
   );
   gpc1_1 gpc980 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc981 (
      {stage5_4[6]},
      {stage6_4[1]}
   );
   gpc1_1 gpc982 (
      {stage5_5[0]},
      {stage6_5[1]}
   );
   gpc1_1 gpc983 (
      {stage5_7[3]},
      {stage6_7[1]}
   );
endmodule

module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor_CLA256_16 compressor_CLA256_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h91305fad1fb10be9c862895dece718a69bf03b4bfc67cf3ffbda78df3dede528b10f9185bc04f59c10cfb350bba48d271fb70a614494aaf4133599edccc7f2ddb3af404772486ab3fd42b2efc5fb08870070c3ba53acde24840ab41acfebf4b158c772c2cf9bc02553c846431c8a2deb6f3556accdaf415c04c9395a3baa0dfd8fa4d8b395f9f4eefb75d665bf63ed525a756bc77f7eab41c96c219ac875c4c7a44a1a2be4d9a9e9b708650029e003b59cbb00196dc4d3c765eea5b61a440c495bbfaac447bc76006fe49f266ff28048899cd5d032369350f19d77623372d14cf56ab7cabb3c92cb8730be66fd72875396ccaf2da06abe170042887680c42802daf084f91c0a531c1a4d1a9a2b73c63d3c6a18ce35cc4037f5befb68528b1df5d90999f27dc31c96b74e74649b0dfc8c08645fc5c6c1be1bb243a1f64982fdc77c1afbac22b38ca951c0bf9648255294fca31a7ad8b41097638cc3a02fab0462aca81b4dcf5f3f5e93cbaa1c8f90e3ef2217f297e45564d0b7046092130d1ccbf9967f5a3de00f252b72830f0fad914e28d5a5ca046de9104cfc52fbff2615e3c755b38ef4c6b60b850f559b8d1fc55a19d50bad1b23df45b13375987140b53486f45e0648174ec9e7461ba372f7caa9ad80698fce4f06270d7d0c1102d8816fe52e329528cf3d1f2eb3b77e0a32981dbec51152ed913ae399c865ad41d6221a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h42aab26fae053efe59c71d364a8e10829819482fa07ec053d6d37ccf6d1af52bd2d8dd997b04bb8c7275375ddcf477a479f60a2ee7a9b3ab9784d3bbe0fc715bf13c8ea42eb87a70a2efadab22598b2bc2abd1d09074019d3c82480664f73f56567c59d738449364575665e9866aae6c84f70012023f4a9392e63820f1b02acd0d5dec4640d78d49a9dd83e574a521406ad369d2dff868ba2d1dc84b21d545e5ee5f0f821a9521b056cabb4521aba1ba32cd9d8828e0fa42ec23b744dfb4119ffd7be1c1ffb6c16ccde2b82953c9de54f2fa89da2d325e987a2f8e0a0a337545ed9680aec3d6f63660deb47ab7654e0019ea62a1ee551fc520afb7e815ccb1367bfcfea818867755adf64cc107890122a40b17b55465100abacac66432be0ab5f748251028c2b606146d1b78a5c9a114340d8620ec8bbbc00967c841a4f62a4e43ddc72a203a6d36302579472eb703b64f269a2b1e4d90df26e6f33c8e33f6301e8b47426f7966d3cdca651332092939a55c4f280f4ff2aa61122986af7619fa668f279e0390dda63ee6bd17b6658c5079fe666982ff15df7ac223c1fc61a2e0f22319f648d5f513b49724f50615888c3a5361f3d2d95737adc102ce4f6c22ed6333524d1d70fe4cee64d99a587960850044fa727b8706e9ca566261fa1090b4010779869fbb4774d91147b01638814f94ec0901ebaeef666877cf1bdefd9054;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8641de93b0c4c54925c6db2b8cbc9fb065fd8f84920e158829054ac3823835c7721d19095d7c2c014c622d6cc079119f67246e0cdec4b319bb017044cbbfcc764c09cc3c967c8fa5f7bf9a583fb07df6bc3bb8065191b793710be9d16625d835221c735845f36a4c85ea08a08a4bde336fa753f5b593e6680e4eacc0092668fce8fe86b696205e12d888ff8c3fd8eca4dc580b336320d2ce24abd5bc5707cf846f92e9035551bd72d049246c85ba5b57416cf6cc646caa7c604d88dc93ef172044f23b8de50f9a80dfe260ca1f794d0d96369f04621146126aa9b43ed4f3faab9f5f50b09aa6ff2cc9934156ce550ee8c6c7df4e5a786fa68790f92904c23375592c39da062bf91c56258166b980095405f6e7617dd4801f5d6e3b054bc5dfc566be4803bb3648d20bb83476bd2025e68803e518840215fe6e6953c956bd97644897b4b303305d80a3552afd747bdea0b2c968c71800dac7bfd9cfc77df47a43de9fd140fd494d66ff88d6fda03717fa000f97afd6f54c203db4d251301a6d87f1e75e7c38a0df1f346608a44b1d97e7969c8ef4b9df0bf74684da5c68c7a47d40c8e04c00458046aba3fd0bc263683d4b6b69f0c2164dfe0c0a3f3011a5b82f2b6c7565156a70d6b4c481af0d3a33a00ab38b8a45ba4096a6bc156ad19d4bf6bff35ec95075885e46e0cc4d5aca3a5ef013a3c8cb354252b6eca1c03dbb419d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3304ad3864ac1f7585b2f20ecc11eb0ac677aa5b664d24bbd0834fe32465fc659c27005eee779f4b324e04e676590e5c539c30a24c465f7ba0f56ab78ed26cf108ca4e97b2bdb0e1410e4e1b55ccde5e6c10c4c63922a046b11aa9c1ac5d43e4dccbe281d6e801f867ce8ac9ca5380b34ef80bc84c80e506376750d36fec644d89b54bd00708a6fb1beddd6ac96f8f96c8c1ca3ceb7298a18c1d88a5408f53cf863eb0a8a188cb05c4b2a165d7511d9b4c2005d0f8f248f845983f2b00d1ebdc977bc5a5a473afadc531c8433a7ed0e34dc0b6457fcdcbf097eb903de2f001c0a96e0bda1053caad4f41ece7dcc18b369884a884b4609369df0944427598b3838a98c33e6a75e70a0990e7c9403765aaa8946095fee7d3a86ce4081d3930336c264e6d75be4d6cbf8e6fd2cbc4a4aeea90318e8c27e864b509779034d4dfbc2a14bb408303248cb1f78fe8a8cb817af895cf195b4df1ec91b2b157987f100b39059520805efd2c626c04f514530d8a28771adc0c0152bb13eebc7254ac500a7e96ab62eab307f532a96e0ffa5c3730bde46d30e6e1fb3a8af27ec3685debb2ff49f9ac7e3dd27d6af11c0e6764a4d3cc3b08c596e154197d03984c04774865f16026626878aa7a2fecb0be55586913ded77297c8d2d0948de8747f3e5ff9521bdf428c55a6985c8bf25962de5901f6ebb3d9648ac86c3315004fd0c14837c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h121c6525e31716c7e879009893d73f9d05795093105186ac14e95c22a6c53cb3eca806dbfed5ba0886a1edb9eb1c9d416ff45d140b1f3bd0e51924a3aeff713281ec077f0a58f962187e823e83d46333b9da59841d2a5cf5271102d6e1f17149b9bb316bc9d44444041a53c82f4288dd86eae30d8f794ea94089500d8688fa8416b6268be48ec9754d5c8d8a02c262c91609756f9f065cbffa2142df36fc95092a5baa84bf859ef96fbc38f22b20f20f354d8863cdc04a44da28d4f508ad31e9326eb8112f5306f51675a2ef15789d2f5592ff2bc80e329d71744690fa5f9f244996da317639ffaf35bd125393277325a7eb3e0daf662d0ff604b7f40655703062e6b0cd15f2d60e8dbda032c7f1fc8965326340df7f8e6383cbd5ae1cf8392931a351630ebd4b275970e23d71b5cc574421628ecd66239317fc2061d3f6a9b1c4f79b1a8d2f70edddfbb24f0df899434e1baebbac0eb523e1f0f7273e9acb9cecb5f81ebe7a1c535343baba16b822ce954b7cf72be720415979aad0ee4454960a4a4e85241efe5fe526bff61f44ac85b47446662315b3e045b10f73ef5d4e9f5e42b542479f319fa62094027a88f7229d1fc0c0df4067e3155fd7e28261ed0318d9418dd6bd1031fe2b599bcb46470ba462d44d0dce3a7a62a6f40a6a7053ea6168c32c3e8a75ce256f7807afdc4597bbe98f4aa95056024aec6cb6cfe95a98;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf15d42765d58588e11a57900f3443672d63998c274dc3f3d787429c9d0af992cbdc419117b9d1dd6fe6f0a03af02160bdea5d8b762f426e82f2660c5bc1af92c9aa0e4138fd65eb982b624a5663ce74fbe14caa3203d7935ff0536d36fbac8d50010b60b7aa5de335fa28815a8805c1719edf3cb2d5d87b7f5030cfedee75ded6a8fa8f76d345136f7b6c07cc8afc632bb4aa5912d1abf59512912a57faf91388445c632db4db5941e7bc9534363c00748df59cf09ff5cd72e6983d12250cd3d46eacbd92b9b2a257e402c9403eac3eaa82a181104e687e5c9bcb1452b04db7bc5d25305547907d5afa5917e28fdceacbe7499940cb9e6c3d6a9ecfff630e168a9673012eef7df7f216902624d063b16e5c201d366dcc3b0bd671b7601cfea69bedb019282cdf9da2a4fa814778af7691ff68d50a9280c3e9e7bbac0c5a2a1ae192c15213c6f2d57ed5d97255375f35bf6622ff0dd678e77f203c45c132718630145e2b0f563e81db0fd246fbccd06194d39b9d1f90b38bb615e2207bd28c48ae3b75455f8354cf5bd4ff035e4fcf90d9de2b316f67bbced4d2857aeae9da14d52000e9e01bcf243922672c2a7f981a07b25bb3e8284e5dddd231b50da482a5274b3be54afffe7152ec0ee0c48f86a97c946eea3b016cb9e2c03eaec6819d4576765178117fa09f8e955e590e44a1de65d8718ce7627e0598814d2a14a6dfc16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbd22ac612c600d3aeb2c4c4719cbadc87ba7253d0b7e2c0acd4d753dccdd0b0fa301e87c382392315266eb0d28e10e804811fa3fd6080b437484ccdbd6b8109066f67ccedec9e70b220a4f3661913fae6024b2c747333359ecfd5851a585e02c55176b02f8e552646cce9c2a2c93ec59b555fad17eb5defc32e62f6aa4b41217158b4dff686dd848da15449ed495f5742df8151fdaf5283a3e26dcb5f40eb60f1f3a0e9aced139e658d4b43e319a179801d6d8891ba5f3f96ab8b718718d28fc97e84d570b9c78f8302b3b3bb12bbabf72d228ddd057152ef51249f37aaaf2780d3b25d97678e401110c043f552101de7a34ea2b5373b4c7fe33a40a56411c0479006402cffe2d5804a20565e4b7b8ef3528be4d3fbff0861cad6f8b8611c91699af22aa94b5535025289beb554a6f485d442170295eacd98466bf64f3a8e87924e888fc957c28ba7c47d49ed405b0e323939f73aa53e92d709d78d5cb701cdbde06accc95675ae38daff0806f4ae6657f905facea20355e01deb366991786c67176535821dec7a035cd3287785dc074ff62c4667f65cfebcfe5836fb4bd986786a4c418e0f8fdfd3f943ef87d6533811225c4915fe180489a23e1edec37764f6158a53216dbd45251ec3bc4a0dbf5088ab104f41915ca07971362b8ed733855ecf816938127be9655ce2e9289f901b4b49bbecde11183247757426c97e988c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3256f2ceb48a7c7a4215d485a1e5bf0e55644ee66f402324f606d38c4e9dc9ba41da157ff997950d60f2ef29d4f6fe32330118cdc483ef4e3966b4be1862695ea57429988364e6b9512cb8fb2a8942fb293ebb35a6d798a50475ceb90f194ffc52db0d6fd5bfe3a9dec1559e05a9a13fec450017ad546bfb5e7b788a39d43ad407763ce9cdd159cf16ee4cefe378254aa117c64780a6ae3085f48f738103fcbedba88686a8eb6a2f4beeb96ed8806fdfeb67af1b6e23527a7f38d8c813ba7fac69436b58b84538a9660dfc91e99133dbdc88d5f7f87c8e8f9078e9272d366275c1c931ba59e6aacee54b6e5b8be5f5f0521087e4481973ebdbd8e43ea96fc9e1d4ceb304bffaf974f93f82cacd914c9d0367251f9232f6127cea39f83ad1b69cb5d91185335b2f372bc861eade1399104295d8a9d3a1c69d462321b39cc4c10e77e1dfcd4536ad156d0ddaefb42f42f8712dcf35912d73384e245952af980308500d39d9544713950d359b4373230efd9de562405421cf71fbe823f7bc5e0d210e54dcf0c7a3dd2983209ac2354d259e4fc6b561f6760d73b71d3a33c6e833cf36aa16dc2ca8df4ca3d3837160caabab5fd0658aa157b3a1f0bd29eab7a6d7febb92ca894bf9928a3cff0abcbf826bba6b09d075483faeb8890fdd6e6bfb7f65383a43381a4eb8dcc5cb36fdaaec0daa5468a07c29db4cdc8f3e709e16b8204a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h448d38c4771544d0e943a27eeffc2e1ea04c82fff199923de9aed0878af4731cd13b8857c690e60b15d277b6ee146e393d4e25160434a2446551692d8f192b53c4168f475b8490983073dc5a4cc8483d0d76e644a5ab490c17f0402624fca3156b072413f68144c80f227c58df05d9b34680a1a034ea96367c659bf16a88178e1227cf6c4a7bc8cc400bc5247ad01affaa701aab0d0ab609f50ca318dae9b882dc78c6d3432801dce01cf5ef9032d29bbcd2763716ea8abbb3464e15f4aa1aae6f8b58ba7349fa1c2055ec19a02a6f5266599526f835040463a6c54dcae609b8d0e6753a47ac571e5957029cd972188be5f3fd845639e70dbd04bf38ae798d391df5748659c72217e34332684cdc3e7f928a9192958b886aceb51ac6cab708911a9eb1e5485d9e8f72d0423f244df60f58d9d76652d402124b97670fd43221e45d9fd75c38a159034cd88605daf9727a6bc8d499c448d326457123b12d9d5e7c42b621f0e81d02f416c29a033a8c4db2a7859c1fff0058ce2d76560af34624d11bd713bfdae0cd7e40d74709d75e1d566b5bf2fbd7190e46e8fd0ad12a4e473efdaa3c7f1bf4c077c7034870ee31ef185b605551a822adf993373f3bcf96d44675a4e1806394d25ad954f0b144cbbd611a9a0d9e8b68f7ba32d34b813ae0efc787c7fa973cad3c16617d0be02067b71a6d4a9c97190c28880c77cd896918f4ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7c421e84c78df9362bf575a1a3e72b45cab04ac69c1506f484680f618659a8c7791c74bac6d78a3710f7c229a365fc25016ee37d5c18d45166ff694ebd1b5fbbed00835a1461537b1af77aa037d36230649dcbeba500fb7717d3b50acf2c7b1348aa71b46329f19d9b5e1c438b5dadc62a374389e5b97bc135468b38cce366cbc232c3c5c365a1dcef2e65c42ee39a67d09b3cc684a7b08384785e0094d2ae0d321c3800d8ec9672d52a99ffa80a4b388fc5aa4e0ddcd3e28e00b4016c687e8d37faa7ba23b14dede1e0b3f73c4e931269e2ecdb5bd58f2005a1a34ea04db42bcf2171a7b3572878b2f79dc723f185d21dbebfe444e4a039fe8d0b210724786b8b75214dc4fc6cb9a18523b19a422353fb3db2afb358c1097e4bf5b81cd48e05723423571951b442d3be8ba662c0b67d70becf13408836058e20295a3b823e98f75f972ec864e99dfc1000bd2a3bdbdf8ea2db4057e721d7267a6947506c0a057e9be02b68816920d6620cfeff8b9f20ea28c59ae5f9c683af9f71b4944bb93adf962d68ee63a2b69e846c186d94f990aaf3b66fa4917d20aef808d7766d99491df5b45e5c6f4737789b0ea8d83d0dd3b0ccb682a7c52389c3ce3f8c4ce60b50a0eb0d5048d205d6a4a8a48e9cb0c08b9b88cbb9d224df105631af72dbe85fe9db1611506af900fe6abd22267b70aecc4c25afbd26a264a0fa14f8fe6a51845;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h489e865954f38ae5ce0c6ffdfb36cc2f8ddbf98bc7996b941099736722c6d2fbf794a64045cfdf1c3943cd299558eb27aaa2cd1bd59bdab2ec4d32eb3b1e38f70228e7980f09e3c2f8b5172d1ba6e4f14099b5324a05179d9e0f9d677c40506ca5830de73f1370d10da68048937234269fc9046b9dc59681a02bcd765a22dd33d83ea099780728739392e9d864f569b81b0869ad29b7bf9e184b19ca91d4a9394fa75fd52efd4f510b55338ec0728e5328849416cab8d73137598ba041f4f8185d57b6e0690891b36563c8953397a85d61a3e86ed473f4929019fa6b525dffacf9580fba80db5e87a87c2654ed9105e7994499c3df5e62f07205954eae0971ce7a61b50f2039ad579f23a7b49a96a81ac709bfd2d7a7343d8d26906782f9c9bccd3e00c8600403d37cc3cbd36c2dbe55e696813f4fdd33da6adaabb96ae060efb1c2d780e427a787aeeeea79541c6d7a30f79a77d526dc6e5fa3d401f5f27aec76f3bd662c4b7af39100e79d498e516f104d6ac075425de0f90e0ac4bf350f01195b7320473022f9ff6621c10cfcc4c8f6983799b13d6bad329207fb380be6f207ad29741d1d36f44149614582fb993b576958cd09e39418148a2d2c9655e3ba90a6c23706a2a7803c217be8a5af956b7b13c1389032c6604b32d45cea8e39d5685315545e118a8f416d965ca1d4ac5b91afbeae9308f3319d0801da6b64e8fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h71cf94e7835fa21623ad2a371bcc247e86c8a2e5c6d52d2b4983d1b0c72b0ba89c25a22fb5d83c477bd48f115a8ded1b90980d85664a6c565c190d2693f6b2cf44bf331b694b4dc78b121ca0519075797926c61e8855119710d16e4d075f9560b57670bfc13976eb4896ad84e35cc3e40c8757987432159727a56e18fcd2f4f8cf561fd4bb22af5e2eed9b6d394bb5996800f9a2a88bbf4455391471cfa3e5a847e07ec7366b269b83ae70fde5a5a52d8d181ddf15d63e9220e526db660aa30026a5af24c43bdc1719cef0e7ccc382eb57127e2c303302a9bc7ef02dcf69ba455237626884287e3d6951a177fe4eb2f1698db8ef21f132a4ab0b4797229686bc46fd516485f0acb5ad5faee04cf08e97114bdcea5e7463da66d60e91deaeb30bd458ef2333808322ea2e8489dd27c944bcee52eed03a6b2b353eca8e0d3d766e522a783bca37b46174b3696f7f9d2f8235e22de4773c0740b7a7408bd890cbea787780d0a23fbc56e3765bd31a984da3e8cafcdbd0eaf81faa3a2fdcbf7aa569bef73ca1064241aa8614628d89eca16191d19f01f29a8f8ef063df2084cbaf09c4808f34e80ff14e89b564bf832e824fcfc343d40feb79e160475356c565c893623516436f89ab2f6c0b5baccd09c94f7c04e048204eb57a34d1157b4634d8070eebc31b05ed03334bd6eef1d4c4cc6cb21bf06879bb4581ccaea709a6a95a86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd24aaf92bfeded6b6d3568152d8c947ef7af7be56860ff185001b160f286d101b09b370da9216823a8b736266f7eaf200f4055d6a682749426dcf8211df31c134dd005595306e0a3f69df5c1774fcfabc7fac535a1c7363ae249af8c431a89220f10193612006965e86116c879b62172ca7db814bc3821873ec26e13d67fdb42fdd74514e368d79f6efa9f1b07cb4df7343841af5f91b9c050cdc452c0a0aae3f7210013455e22d5c750bcfd4f2bd59a2f4fde26f11e5866c1ce5d29d7e08669d8cb2c01f7fba246cd69afbadda41c48193cdd5ec7dee29b66371bc648ff65f7cf0846ba739c1c30d7c238f36bccca5b5d93419f9a804bc59dcb79311a3bc9d6f967fec8c1c3f1e215619c632ab09bc0788e8640fdb710560bb548c02c1e339104374df29f51b7c996d8317db5a14da0f24648b1e5f760057ce03cc2c2df5dd10f5aca4db51cc7484519ce1921c01b15db0f7d96135fe5e449e31fdd1318e625ea662f98b07ea5d2be77b62e8404402315fdeff1ad8e1b69c80bf54d46c0e8d662da4bf14dc13d2f597492b556515864cf86f5d3437d4c07a5f816c8bf0117456f730163b1eaa1e6d463651ef80aa8580d2d45d566bf360defa6b1864f4f02a583d7fc0ffba154e983e6a9781e0c4ab8514abf1c7d3148b3b080b7978d3b97e2f50286d14313e2f266299435567b484a05e660289fff62d82ac724e8eea2b1a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h779851378fc95c3f6cf1b0c830e312d83a875c1b2aa03ba449387c4a21c7678b06b00cf6ba4770f0c8857af91fbf3333cf08df0c0cc9dadc56aaaa68bfdacf39991b481004c438506da168f36e27bf70f1b99d4df761eaf4dbc4c21e274b30073c5b6aaebf653fdabf7ff1d99102dd12e0c7e62a53a1ebcf117b7dd3212993ae4ad3d1558089b053b5562ba8a1aaa54e3e7354cd07388b8a7e1b52235ea634a2d307d652e5632588dc55628daec9e7b1386488caf5b1a2de56356e9c6d6c2ddc98eee226470bfa8d3e348f28de32612be37aa56894293126666a35137e55ae5c84c9a6fa027e36ff3e311d0ff85a4774aedf0fb6b5ad4aebd7bad1bed2714347714f6637d98fe6f3bae42eef825ebccfaf3ce8bff2c167e93c1c250a32abff98930c0714d6e67454f514c0983e863edca80f06309311776353cdb13be789502d4e2a237aa82e061b6e446c7e4e41d1a19974b6e6859ebc4d1200f4f55c708b9da5f0ce2f95792ef1cbbfa7ef2595d80fd5b06090d471ffffd28800db2b11aa79e4881913ff772e98d5d77071c35a8e0efe7f7877e3208f393f3748c0cf93dac78d61b0058d50cf7688e9dfbb0dbcb862395be362596968962fd5369227ef395dce2fe419ccb7f7dd386d1c998043e012d915f6d0e1d872dd838d01a0b89d3fed635d35dd6cdf588ee86f1b55798ba560ef7e7afb78e28ddcad022dd62358954f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2e3b5ff879e249fd9a1383ae4e208a5fdb4af6bfaa045f38762dce87548d57c93dcb028b51e7bb1e6bd269ded21a4c6d10acb1476795ad9eb61df8b50a07d63e600a37f9b3d1482c68a7bd49591104195c682d2167d7a2bfd2da5815c180238dfe60e9b02ed84316005d2f627e623c1b180c0bade84944a546442a3e8a7819688246aad7e84a602d3c158b968783d94837aa7fbff59fd13b246682a804401fe3f8a1481aea3472b1b4028e07d424f2394f381a1090d286ccfe922ea40ecbe63b1a70aee18ff2f92ccaee5af2b6fee16f50adc49722f87df9164f0c6de47d843de80d0ddbaea6296187ae39253e27f589d72cabc07d40f5bd1473e48bfd90caa9c923bc90fa40dbb1de70540dc12b6f71dc4d71ea988a61ada250a349b7c366c92a3b8f407195b6f2921aa1ce233ce940f575915cc505f31cbd3c8615b3a755d388ec68d62ffd27eedd3fe5898eee6f0c3e771a9941188c241461250bf9983034074cc7c9e0c136d00894e168a82b2d6d715fd4d69ee9e344970a33e66e427dfec4e92cd8047756e4411d5ef0b4711e6595001792856f42d44fdc746e4a61e56b25d1034cc7bfbef85b0c50aa2a59f27b22fcf085a7fd2ccaaf167603aa3a83978b6b966867e8a9e6da1d62245732d79a5a29f2df836ab61b5d1111679f109352cee4270b0cff4f1a2ad80b1fef2068a246d694666dd66f4f37b05f3758fcd024;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h327e34195be914df81cdbdebf252ef078969721a4636ca4e155755edad2ba2dd62f7251b02dc27e1c8fa49702129ba2e372341b8b486c02b5fb126b7e9306bfc1e1c0114fa0cf7f5c495d45ab09a6e4d66206d0e888012566c1644e173d50ab9e8b5a894e59d1a3ceba848281fdf47d7af2c0476a71c2e5cf1d2a9b010d160c1686c2487deec076efe7e5c9ddfab72d308b56fa048e66c1774828dab12c900b0a4350facc458e0738291bf970bade9d24b10ba946170d1d2f8e0180a8e0ad02a895a07e2b4750d1d603395988d38e5c17d143387955c60460e6672d088ff53a424993450fb4f643b64a02b0ae24a74c48685676fb50a177ec2ff57407d6e49236449962d28ca3b8ea6a40d2fa24ef8562832d34a52e6d30c8926b9969cfe826e62738a79feaa66e7ad12f96422d9a43694daeaf9d276ba4e3b76e8072506290428a43f31511093c7e0161101bccd0c6d9992509f09c0fbd9e493e82f9d910af5606d7ab592f54a9d68df21bfcd5ad9bac5df5bc75d249fa817391bae2761aba1b4a1d14dd31e46adbf2d31eb5bc8b85d374d1b64970a9ef7ef5a5b5c83570820c591eff711e5457935d548c6ecf64ee20b75a43540ef25943336e9f623b9e74eb829c71f78d5f103584c3610b1dea72d3d75ba21ce4fa347b57f99683661f21d1240c62553048242fbcd77c36c3c2890b6cd1aa8b21a8bd95cffff34d3b703d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h57a9e1251e3e6615330ca3551edc721358dab72d701bc59be7dc5215d137a492f3dfed673dd096b9cfcc9e56f4056308ee38ef91d2351bec7d18fbf7c77fd5df7d427af21a0dbd35601d9a48471a8bf1d6922a87e63230235ee14763da995fbaef788cb01b81f8bfca5a664bf74954e05ef6a03a31390189baaa023d912749c1d08f61ec0635b8b30635c8de49b929ea3f12ae30959c2258d35d92f5afdfb9fb64797166425e8dcbdcb3c95161d2aad338bfe3f7f38fc42f7b5e808f21e62d26d07043c7be4055fcc4065c5eb3e37fd2cafb2d632a7de675642e3a367c2ecf9cf2d2b12aac749c5cf630323344209776ba31b2098b4ecd46ce0ff5c4743556cba159ba6e95f5cd195851b492adbc75dc33502387f603ddef78a9056c61e611d8223edf7f4c0ee25a3ff84cb797679807b135e8b24dd59fd7a22458ea0a6eed8da3fa95c46aa81d8e74cdd9bad7113e7ab3630423493e9c841b7deeaedeb694f315b7791e38ce49a01217f7bfcd35422ec247f06b97e5732e5baa8fcd717243c1a2b433efad3b4642da02cba2454c3f1798bc519811c5fbbcd1c83c8ce2bb311ba200500b157b795c8e81bcba89ea4e1c0c02128af9c3f290078c44097013854bb72e7e06db605fd7ccaf21b75c7eb93cb411b48167f5f18a87bfcebcabee3df9927c73ba970e4832401b04096777791be0e980b251e888a49d4aaaacee56d26a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb78ce5e65d80e2714ecf7b2e7e5066ca8950e2c5548208065a381b0702e93698775a22918d4831f94b89dcd00ecfd0a8cadf5918e8953eacfe1a9463a369e5995008d79858a0729e7bd0a0b32f21442e30e3310d9e15a6d2ddbcd7f1a3d1facee2fab6a483bf8c4b04e5e0c72ad6e0f7d26511e132efa9f8be9e85bf8724a8d12020da7e0d27a26181a7f3ae98dfece933d9bdd3d3165c60931face99a6bdc88fd71de632187c1a8258f8e800222154080b71fac26fff467f56145cef16f0e363a6b7fbb682fbd3e84f5ba430c583d89a94646c7e22f331a95ada24372acb8a57ed1f7aba59815b65146ae50f8fd38a8ee85b8cd772801986b3b8cff1329d2ccc23023afbb1a6701e2c50632880447974558476a5e90fa9b7b612fa79105d599705459b9ae51fe51c365b545b3652f08752d84c3e3987067b01060e5e08004c07e47ca8fe2206c58b4455cbc221dc407b0b2ea497605ef40db9482496cb279921b28f76d7e98baef4c8a6bd03299e1a61c58bd714c362df55dd1e788d62abb11e82a5c717ff79e88158a0ae7fde9cf86e202dc0e9d5618fbfbc1d74fca4705dd74e566b97cf84176c362707787d188ea1faa6c728f8db527d4252c8c37436eaeed31fec6999e1678af80eeed4b978186502abc885f31c9d9ce2867ac090c2c996824d57a862c4a02f6829d3685802776669e46e6834d50bbc06e558b2d5dc670;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf10640a309f92d91515c4ebee4ff98ba23cea25eca344234a25c4073f2a5e2349589362f6ea5f8ea2eaab73e6048e99194812a077c3b7e0739521bf338f539ec9ac948f1c1e78383a2aa6fa54caba8da0e3ca95908db2074c29d0a78fc3c1e1e5bf1a540b39e7a15cb0b763a991937eaac0b96c6bab063648a910c6fb1511f51eb69b8f79b7c4ea08ac4440295a9f3a5b8a397687c0d54e90949889fc136ecb576e8c84e83be35a1b05f0a04f7b95cf6dc3e20199587401119a7d96ac18e84df27997b6d0f7c0c8fa734b82f27e92aca5cc300a6406cc286d4541ad8f6112b034f929811502e8ff7541c4b245bfae7d6c71ea55d757b86c7899f8824c845b53dec4440a8c0b5db0a569491f9f33bc30da7a69701c51fa07e489929c7cb8f41dcf03dab886a57613f5c12da4669e6137aac80dae06b2c6c56d428ccccf556609535211391a3fb4a1a41ee32305133ab76a98da2f9d07309f17c2e5acbba338c02569d7073940aa0fc9b342bad9cab111ab33514d6e71398b0386985d6876b8f6e8bd2cd4ece5d076dd1a3d0be962c4b47b259ab54ac9712d147534ff6bbeaeac425a577f38b1c4d3657f3afe13bd10b4a001a2f248b2f55eb737a29185dc45d15868c8dab76afd873cc4b846827cfb37f3b89a7ea10534964cefba9cd82a6139230097cdd7f3b35f8796a2099f4b03b0f4475a7f0ba9e2d650cb5dc0883c2d2ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he57c3f2b791faa4ad980c3f1035d9c78724a581db5d5b028a1453f23f37b25ec69538bcb484625fffeb04f306d8e05e9e2a2ceec7e89c0ac32125f714dd651d38b2424f7079dbdd124c0905608d27a141b4f344ed39d792579ec2be65740f467c7b2be21efcf54ffac5e2cbbcb8ba37aed1c77af2269bc5c719932efc2ca4935fdac80f43122203c84ff5d6982c366aa8b728958e35ab57d320c66469c9761c08a18f06b6a435858e29252931933ad53979c7e152a508bf4f0ae9052187f53bb297c638fdfc8af47cc324ab01e08474875f859ddd6afbec74969933a86fac335a3686fff2954c83a73373bfa9b819d89feb9feaed5c9b7954b057e7261290552838634086e3a001b53e599b3f997dbfad43ed8118e4e9217f642d73c82f619ec400aa637523809ef2dd22b8fbc1ebbfce723a867c0f230a8607c35ca7082b0d89b1b2726a4ed4dd46c8eb7f9193230bfd05ee19092f5d86ef7f246d1332749c096201552f66bf93ca2f829aa284fd630d392114ee27c207af9d5a8673de8b672044f0cc0a5f62f99b19f91921f62cdcbd6faa7c64ea5f2207798208ba5dab79fac61496d619d0e52ab263ea4d80750419bcb4b8c1b2b6bd2782fe61ed2a2f34aa57f45c82a633140d2fa8826180853ebc89737fcb85760ef49337dcb96ffd2fbe3c21672a3d73494124527011f0e90c3170646335720114f66f511ad680bb0db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf6fd2cc5a990557a0800a6de8a9114d7139c9cd96fa8e6282929a94bf1ad0fdda23932b2625dbb8ec618f24e2d0633da8eea1e75d0cfbd0424cf9703d66380ba805541fb7cbe4638d71df1aab60a66afd0015e9a3bcf1b7bd3e74fa336ae812fe4fe66f7f56494f3eeba2c5073343968267ec6d352e268216122a5acd2941a59d4ba2f8aa585e5533691e2f0e97773e54570ba57bbc40173bb480cca9243f050b0508e62ee6db448f4e4ef31edb16ed80b6af35f0e4254e251be15cec9e55618c5fab3123a7ecf5501e9e38d02a83bd3ffd85f85f2c97fda4b0589322e1a45560f37947ac698889dc1787e0c3d4794f8b147b58118d4b518d80ce2042f0955e9d3854b35a968bc130a2b708ecf63acfc02a008efb09710d07c8f27c8bfea9288ba3050f40898cf9cdd546687bc278fae3fabab1044f94e540347c96ac039310f2ddbf5a843d9b8a0f841475502e257fb883720e4632b782d9bf3bdb44dbf5fdd0ec1b45aafba50c28e0eaa6a98922cd6b2a0ca02965485c3f7c2e06f2711f7c1facc93d39f70355d634e24f58313d634f7049f37f1c1b616d30605638f2a97c51a8bd66cc633bcd11c980c64b0724eaad1fc825d42c97ac9c7df1d3914c5a80a1e2ccea04a0ca604778c783c55989457f75990d6f7c52f06d9fc673c900d95d55960e06133950b691949ea96ae56891af54cac166581114e3bb88c315eabf25b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h94e7b8d0ac2324ced0d77b2fc04007800c5073656744102a680114b4a8bef9eaa974f3d7bf7f0d508b163696118a20ca68a73676d68ac4a759fbf900db40d08e730e01aab017a25924a16f52ec9010a6bc16b50c3b70556d52895e54fce421ab8d3043fa45b26b11226de24408a581e88ca80eecd5ad30b297d28715adb47f74281de2cdbac9d077b34c4737b3fc5132a614619d01b42996c4ebea776cd62fd7a84632825cca80d7f999ff68737fadaaad2c50214119a05b53d7ec512d9f548a1c8438dbef7e78c9c0c91e067074baa17c0abbf40e8a790e11622be60ca4ef0da842d5a631b398939ea2d3906c50e19648ae1acb725a214cd991817986f1a89da3411e9571aee90a2f8f0ec6885ffd88656afb91847fb62748eba1b2960bde0944cc6c3662809cd750770ca99ed7c07b23ce40a9218f831835e663691314a5c4f185a2b01be2acee2ab6da2334654d097b74785c96fe74e77a7ab636ca6b002a47fa0a87627e675ca89fadea5ef987e74d38ca96f62022da0715850a399bfa67549e835d5ce0fd17eddceeaaf445a8a6be51b5eff48520c9109f10b21a09574d4653d4661894ccaf87c03f5daf5433f5f618563ab00953e06e06925f597046663025ad105fa979a042500d117be32d6e49bc727542468fd5321b02c35c58db73177a040d608d861b9fe3b22283e74b745b8a2b991249d2de488ee1deb86f03f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7874ed00ec4446670158cca483237973800487d330fee03d6fc917a35bfb364267b350da0986c77052339124b2d39b68d247188bb754f81dd7d97d9c69633e2f119c4c76f7a9d865c56b85fc6ffd5d00abf29293325db38d33ab52b1858d4dc953076d953890729136c9eec83c3428324e96efda32c2c39ab132305e1035fb9320c9cff3f3ea5c25a7a0745a7df01443d4f0487d590b10256d61c602d842e948507c23a342e530fa681777ea2f03f1fe3ec67473f4993a0a3a852b102f72e0330289e4288c673ce6573c203929737bb66701003cce1f047243e2c12ceab184698512f0925a478e8a1a1064ce1dcf24a0740fe9b116281d59e7a91dc54094698b5247f28f952afee1105c28a3f38bb9037a555d127f750742f6d19cf7c2a569205074d226c762357a63645674914716c4a312d520b1ed7013dc222237c64f569e41a7786d2933818cf91038786030b10099e13304796f2e20d1c7ca61d66757ec252b0b9008b4411a41270c8de21809a42967be9c52eb1e06d0d61e07a54f69e61c3c2b9a694c49cb0e0f5d0b07a6c668d46ee189603cc1fb5da9c158bc542cee0519e7dc0a021d8dfdb626e93ee2ad4b086a08fe6262610573e7445c9e71729ec40c0bd6c2ecf3ad58cbf93e446962a9c1ef7be358aca207e4a2d9b19ab007a730a9251a1a5f15dad6b72581867a48c26bf762591b7ad525eba64292dfd2d29d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h64d4269cca3fcff2782dce95731d33d6d529b0e4d5c59b956b52803852daa6036815a7d07cda486c56309dc07349ad68b07d7fc7ce21434e39dff1b5c3c8cafc46ed1ef9d841170b255b59989bdbdcddf55da5f2baac32e409042a058c579f1e7f7dbd553ff11410ddc1db024de4cee32b9d1615e0e6fc4210f95d791d5dc466a9e4905cc03f4075f1abb7efcd9695da968804fea00d960cb7ab81126c643e4bfc8bff91e6c4506fe192f50143080c3353d94f694e07b6e308fd13104708eedb53240c5974fe25349bb60f07ddc0175cc4f0bf829766088579fc6a22d05cab29366e553ebc6453e11d3a0512381387cac08ae2c92d97fd986750c369425155a1bc8831d96ae51fb315027c9c4098c77f4c3aaed8b5eba9d27c0c9b8700876045423c91f227742bd78108273bbda4c7f5787b478ef11b324c86151f2849e4dd3a9651c1d72c54892358a60ddc316eae76fd8d65ca8b449c88379ce82250e574580a4e202c495672ace77c384efb69c1792708a28d606e670150dca7ab16d4e8d812421df9747a4df0ad5b5b55c32833fb7a998677c12458ac08bfa76214c4d66ac559fb8bc5de9afa2238419fdbced8e6a3b2150ccd9fcff4c70f35282c95164c353671d27f71729d8536c83d57113cec4745bf3ec10cc83a8793237c4eac303894b29c146b0675c7296c98111454331d4f7e50db89f06b1a2ae7254da2e8769c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf98b4166041aec966c08d52ccb61f6c7c9236305da9c3a32f0ed73fde46ff9a583660e5c8cc9c7c21c54f3145651ea6db687e35bde59b1257724f5bf473c77409e56fcfa068b95709e71aa16eb7bd0efbe0f12ab1f762ef4bb37d7a408061bcf6986a76036b94f8d93c4e5be442b6eda32e0238efe5cc575b45ebcea90a1967d55b1c94e0dbc8fd27f72900c1f66269927b7876a8a4d37e3c6777fd01f6a06d3f8c5c46c1bb3ae41b51b37ee28c181460216579dd19a82228dba19b5356983c67b741c7e1e57b674aa23922c29b2b3deaee2573c5afc0d9389b1204ff4ab09c4353bf8af035a0054cee8703886219b4c270b03f9c532b81e91985d7ca239f904471ba0c8240997844ab8e20f793062cecaeed1055736ad60196f07b794f6ffa3f522979152c7b11f51237d6d65460078af7b57567b04ac24c7dab88f00afc47efee3ffaa16ff85f3f95465a959c61d555f63befea7c10109cee5140082fd074ccc7102ea2282218a5cb45cb26ed5205458f0c2e512566f967848b206b6f7dd4ad5882f35dddd112be98218bb6af5d95b845746769b6809345de5a2245182c6c49d71a33851894b9a3ec8dec0313ba4046ab1b79a69180b406e70c8481f193d0d089a0c23de183be6804a789bb89cdcd92f24ea95fd8851e02b0f27e82db08bf3ece5ffe7b442450d17e9da708272e092a2b692f05e5c3680faf5111159d42ebd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h725db94fca9e97b116d14d172007bd5ae6bd7a063879327c795c899a1d33a54505ddd9d8d5d253891b11eb8e87f240fff442bbcd4579ee40fb55939a68519a98eaf7ac79862d66be8087bc4e36db5c87b92025f0d428152778f2c62ce037332b729c4c9d1b82f3baab7762a048d145a26a905229bb94ab738b105304226c85e97cd328ba725759a381bdc7790e5fb861985c106cefddca6bf4cd3ef07f0eb40ca0535f3497f1e12be9c728b30ab065dbc096b7548bc8ad5414111e2b8dee6059fa401159f3274f4f6f216fc8cb7669cc27cff6e364c44226c2461b903c9b8663ada645cdcded164867fb1883a080baf4035b771dbfee67c14b161e7c0cd5b509baa82b57f77094f42b4cdbde008ace6f5f7ee04d65adf11db5bd9051560a3f5a397641624ba90e61534cd76dbea8012da03834a6ab66032ee268ff845a6aeaaac051d0dffb60b3f0aafb672727bf44397157818a563238352e4b64fcbe3b5d85c98a5fa5f2228ee75272a0506e721fc7ec72e0cbb56fdf2e3fc13df3eac3c11cdb2836a3ed5464d5f7ac334278161625c7130cd5d8fea2d616a1141274a45b0da830972933e36a74175548ebf8bd90a6ca5672e9f8c78a40a1ce87f8ef93ece1b66b339abe6963d7c8191df77d512498c38c24beec6876152b284395362702262c672c0ec5aa2fc87175d2aa386b50d940b845467e7a5854ca7d845299643986;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h35c82247f811d9dc8cf8094277011c08f0bc293415254252d952632146debece0bd2c3bd38d3e5cb2415f1c04cacf4a3332a38708895ac566c9b26481445767dd5b0f05f1e0fa86d9bec3eda29a4fd5ed5635b3a05ddcf146956fefe6a0c8910977fd94bf7e2e5684b90977d8bc7808697950a3a79557b22d2df1d0cb10c0fbd8b2ef69bd4a94faeabc5356e7e41ea60c1ae338f2f53e406c7777999fdbd7a9186fb84b530eea8002064bd848efb85c43a7e3fc005765cac1f090e006d3d7b5ad14311a0157ec515e18e618801aaa8ad3b23ace1a0e2dc48ff57e9eeb6b424dd53ec420f00dfb3da93881bf7c089a69ccfd87f1a6217a1c69b9596366f9869dfef5cc71228194f9c1e6f5322d15be783a381f2a63c12074c8098227d16f0c19cad98c15f2ea5b606ae5d4258d9c5e9493d04494c69f183625986185af61da24f4f0ac0e33fdaa3347654cdaa5217b094947b587330707fa6dbb6efe6bfff96e8f753ecec06674b8a05cb8a89c0dbd3a28452295e2f2ce4f638e21b977cefec60c2109bc43acfe51193b03860165fa443f620018598b1013a2035991729c493d11b6f9e4b46488c76e6581a8d0bc64c39d39716c6061e7dce9176bd73a54f393cc243eb42828da53bd294308ab647139b510e53e5a8a4671ebd6591384ce9be021fd9d562ff8224dacdaa359cc23c0b59bbbc3dccedcec27c42ca4e7b7b4a9dfd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3ceb11376c3861f021cb0ea40f19c1b9d2c4bad405a050e8262075c19736215f74404c10501153d1f0cca53ebfd1544a596a2bf5aade089fbab3edb2ea8d1b014c59f9a5a774686c4104a25a81847358f867d7fc22b2619b62b350fe663568f475d70c1d7d17c14b62afc0a22cb3375741323f12da100e6da4351f163c0c36f55a2ddb59256c0b864a08a6c27d54a0e99e8d45d81720630ae9f7ae4e38c5143fcd13c89478f36c57e531dbcb0da85b977f96150f114e46875c74255d2752c052f7b426994d68350284c453e27725c342f5c87549b71558e5c0af4ac513abc69a988994be180626e58942fe449ed91ac4555cc8270ea05e5198fa32b41db424312d20c6d719ba9eca82f97cc20db99a5ad07a01b928cf54db5a30b112b0f5fd03b6580af57fb8ba1850aa89eb69cc073549ee01ed3ccc410d314fa3dd64464eb79af8713b4123bb3ea7efaa8753cfeeee8f8bd78b7e15a69335a0a6cb64d12b7ba2e9d61e23d583e944d38fa707388c7d515780bcabfe9f5b8c955197b76cc8b78ac63c9962dd3acb707914b79b6a911169cfa7f0adad71e38d3a8b43b0cf83fa716648a33971322adf8a78c514f1def3fcfed4768e31608c4951115dc28c03eb6785b8cd6b61d08a46e1b73e32a2a73006907a716890ae612d72b43027a7ba826924765f21a6c86b206b237e36b57055e0eb79550338ad80f859c949671bb5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf21f90e170a6adc84d9c156d337aa7279a83e3e6e13cc461309d53c8c90def196bacfa1bbf52aadcb4aef39c44deeadbd00d7dab994388c383f6d73ea8d75b3e0b881ad1a243fd7dce0933e87ce4a7304eb0615919ce705bc809e3e344532d050ecd9836876ea7848675e28381361dc96235676796b61fa4842744ed52002fe36823411b8346a394b6542e6cbe7fa1d0088a74104006cf5aed484c68d3aba5a048cda3b59ec6466a3b74e21eaab84b12236660aa586058efdb7c890050eef9cac506cfbb7dfdc1453890d573edf95c7babf3110ffffc446c04cb385356c1ce01047a390c2c68f5a86bde372d5a58a491cfc67f56bc43a4ed799f22a6e02402b194d34e98e8afe3e44aec0728a7c2b62abda180c1442b7d389bcd01e1ebbcc5d8290193c0c5d680a5a34bab9f6b994dc9d26e6871777cca56bb1018aa0b83d9ebab1a8fab3c5923be80917d8d96e86c25bf80642f73b5cf61f8c86b194a5be41f247b4d3c58a4266d5c30c90bdd485762fed024d4d02596f729c5b0ec6c45180938ed9c18202c20d432c2a3c9f688ca07a1b155663d4780e2387e97be9c9c20c24c281cf087ef16a78de497e9a322e37a708db3d8dcf03b833a89043a1fbecea5c14e0cc4154eb9950e2e513ac5406081847aeef1f530d3e14e0a677012a9e98f9f7ae69238e710b13d3555c804e6503d9e8c9f2d6aed57fea3f2e482408e430e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h47e02702491e991c9a3be010a47e6f29a9cebe8cbcde62f8b46d11914b83afaf164a048517d47fde4779e66c20e71c9a47bad1f510904b2e07b1a9709e5da6bb5760be9c0dda156dec9897c11b8c66dabf14f31e84055f10341f53af295623d00506c584d1c828fc94b47e597c81db711700ddcec9b61f7d90cd63f428dc234a40405eeba691e86bcf63247a127574e225b9039b5de409c59c4b7cc402b52b0097ca757c70cc0b28314deb7ff682fbc77e6d987313b55c6d04e8d34301ca381bde5ab180334c0f4dd83b393c4fb5c822849ed3f2c78a5f8cbb5ee9fbdb961ca6b158f57f539317ae65bd3dbe3e10767ae87711a2c0f5e490b4ad26be9882aa36dfd4beaa538615b8e5ab9137ba5bf8d62b4cfac876f2730e61980a2e983b8ad1748fd361d3f608735967754c44ae056fccb19250b63297d6bb26086109469134efe160a290fc45a9542fb5554e64061f0b006b92e49079f72a864c5dc301d5f06d7bd6b87b7312cde59a28989eb47501bdb380b79b278744d5e3786aa65a373be9874c4d57a82b56c9e2cedbd9c4f2e04e5e9675637fce7f7480decdf25cee096995190b482c13608187cabd448288b2eb565141ff55c6bd66fd47ea9148a57569d6e1e1889c063f685baf2a2879a655430350e3077498ccfa216a3d4551cb2b0792a1d54a7b3ab7be30bf6cb0cb2f39675db17c9fd4f46c3c232af31da898d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3c6dcf2f1da61fa22fa90410483158b462a1eddf59a32e3662f2d389360cd895e1bed7af9d04a504f18e541c285ecc4dce171dcbf5245e07404bc3868748671129115d578e93da64b28d96eaaa890149fa5bb582e64636558f6e5bc9ff54f39ee49a126df02d40206b48685e7def8bf6ae0905511f6ccf372553af097f543ba1d9cc10bbadb93671ed6e09ef98f049384775491227b59f4ed28a5a4224c063ac3b83f59c90ed5d52d01ecc1adb4b8b447a10898257c95054163474eb95508cce09ee7d6f20effbfbff8e77a1f3b487cf7250ccba82127b589c92a252dfa9ec5256302b872544557ae132e18f2543e6e38c19607c990ae206950001155baf838aba145c95da71ef9b59016427674f60b33e82770bb4ceb058e8e961549fcc73a2a12e8da97dbcd0d8da4d7ea35c07ac747a1f259baa01fbae8de3bf36cc03fd32c9c1dccffc2f925811e58d801ea27ca7e3949d62ef9e716a57fd5477186cde24197698da5c09062a79a43e7f9a5137c4624e0a7485012a8ecca50804ef106f99094b0f7ba9e3d0e5af449d391a20a5e446b51a3dbc08d84105fd31526cc7d5a8c4b75068e1ef7ee8fdea4d6ede87a6174706b5a384fd462e4a231f2b60acde7ded0816c316a7906b54f09411c4af0142aff177e6fdb0f990be7e1bbc7e6f08b18b2c8978b46eb0f830be5b18e26c4bacf2c9515f6aba069191e8af0ebe85438f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9b1399752bbff7f76caa1b25717a4a51cf47e2908287f5b3b454f6fae34c5b5819e9dd8f6069b79bc91a3d7bdd8b83c3be5cbde67e3f3d36485645993499e1af8b851f07d2b279028e137d35a4b6946e162fa4371e7bd0d4ad53a0172fc41205cd16d04d2ff84253b8344c13838ca719f468d48cf7bcd3a5bef4b403b4e279f562969136c0ab2da90d637403dbe051967d002b9ecbd0b2ba04a379f27bb593374cde3cccac3b86e522cb16deb44b628060b90f6fe1d897e86a39bbe07935bcb0c8d8f9a41c1667c108bd356559b72ef10ba4b70875a86bcdb787a003068c9e300db1074081b5536dba14ba073ea708d85da637510d21185f490e22e94e4e877b70af81b9bdc52dd4497520bcc8107da7879cd9c98ad00467e2fffa090a18387abf7ea35bdb5c830fe766b93f2916b5cdaeeebe25618eb7c9c0a9ecde825e5f4fd3bbae99af176595114064b4d2049f7be9e5d6b39f3664bb98591c790ad2b49149d84b562d8b76f339ea33e075eff2fa212fa6d3a8713a891d5f51fa5441b3e969942ad21ae2ad0f5627005c2f6d4e38127e31515a79a5a2b3d5c5dfbc6be7c36524681c0ae9583fb02cff2515e28ec52c639e9f1a03f6bad816515c11c3e33275f8aa5cdb459d6be32a0f22ef363efb6c215bc7605ff709593db50e4793db98bb2adc1e3be419b9f6f464fd4f5ebed88fd67138b6f7f398c81a7bcc7030614a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9db9c5758019d1e7b3b1458f46a7f6af96e28bff868c8fbc1befff9684eebfcb811a534d09c803816e395c7fa4e95dc3e3aad93a425879217e8a99cbc8702d81fa7cb8849ca63ca57a18f3171a42d829d95172609045357f7c51f73ab2373b7d16725f597465b9aabe6ece752785751a01b06ad8115716773cd8070b68fb0dc739b9a177c0d2ee71411d962b21c62e8f511fd271dc512464b296d96a739995d9774007202a51cbe64d33f12c36f7c5aebf30fc3281639ccda02de24a365b2c6a114b8cd408adc7a0baf1c222fe9289f4b9633f2743340dae7a831ba258800d89fdbccbb1d51b64646576ba49f3e409477e0b753a65662721b26bb1ad5ecc801fa45152aa2988b041731aae7276327ff8ed4ca7dfc86b764245853800c40329e171ca7d70cceb19e5e95c46f8fb98d0e95ca163378e4af36c4ca3a23b780be7864a69567ecadb023786acb51a40f658ad14e8058ff7b689c751f4c65af5236b2dddc1f01ba4921ec33b0eabad0f452f7b1337c2c91cb13122783527ac3d6b51a2306565f8651b7c3f2f0db11fcbbbb4882c0f94df9fcaf1d91567afb789a7ec966751e5bee14e116c95233f539b5b404571258f328bc990f12071b9f66292ff39c154d3c5cfca535a9cc8098de14ca46232739e1fed4c6a1e17623c36629052c54b49fd4facf939ba8a4c188f5c238ef67fbc10b1bfca4e6d737a33fe86a63767;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfc9aadb3fa283d6fb69f16cfd824af01adbaa8d33f5c0cabab13c0a296594e7eedf212cb528d2fa87c3e71f574e408203229b8d693706a50026c8a16b65de806777dd2255ba0564c77127782c2b9afde9366ca61f68b55289fd4b9c93d3d3efbe01e0a8de7f81106fcc408e3612ca77d6a0652ef4619e86104a452bd3a2880d0ed48bcaedce772474a3bfe9884fecafd47ab659c018c774b2243d6f798cd67eac8a9dee2e0b1b7d4a97a571a04f0303412a98812f1735a4c0ce8cc71c574637b0028656f529451239eb49b9c3656cc84f3a2a5a5e9d546fb219550b5e9a5e3d9b7a5162a14b5d8c03d1ede02f62369d62b6263e097f45784296e9ed1c0da45294db39d1b6c3102b376257a8ee9a60e25a0027aeefe5250072ec821b14f8c79d45c1c0f651a902d64bf523fb7fcf285269f34687c8aace4cc63fb9231d2519e0386d55776c6696bc6865571cc48f0d6367b3a532d0a17a88a5779bf2351d06417b22f8d41c88e72d2cfeee6cdd6f67b8ef75f01c658fd4475ce037008deac117cb8aaec7adea5ba729027f689bb569b3c21f49e648a85bbab4851b81cf68411577286f5a32639a918c76e6dbeb14b919a98c95e56d88db4a54c1192e24c376dac94e1322ffbd59490cf5042977f46db9f8426b86f60c37b34ff5cb6cbdb0747589c1aeac0405753aa3631b62fd359d7b1f24eaf22b25b48fbbc7a582f59cae2cf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb6268f1b5b35e995ce8e7272a6e1abea6172c4ff85bd8e50389a880cfb70b79c9d360e15e2ed2ffe5583e6331c62b74f3b7199660d70b1ade41c3821e8d80341932b01d2b611067cb5ac97d293185f7881d2c3b6b945a69afc9ed51c8d2e519980768838b82436bcd0f3257b13cf17b991a138d51ef05c66b5dc2525a1860ae6dbe1504018b53896ce014502906f38109f4b7883de77922fde75adcf902b78cc9050bf1d076c8f3f08aad93779a664f15ff5f91e028ad34903626c676c7c678a967c9be064e3f788b92e483c2d9bc89359cd207761b74cf44e613fd52c6be0f8b32c6b29f119585750e125b096e2b81bda022980b8362fefb6f73383b783edb44adaa32c9a2a2f5c72e081b2deef7dcdd70973ceda7e326df6ce274e4a9b6c199f1df8e5ff2db4c5732db8f236b925ae42e253f28d3ccceff642cdf151424df3af576876c3969d04e746579e37972ac513da0c564bb2812cb682d22f44744466a37998920a748fe06826737a260badaa5caa3076d426bed8c4e6847d3cce9e036abe74469cc48ea7f547d29b0c240361b5d787307c9706b61ba5e72584d1157de611d6f42d1f1cabf3d1679b249d4991293b118715170ace09eab1c45ed924537f7c8f6833404d7e92763a69e5faa84dbe917987447ac52f5971f22f2a2affbf99b1671a3e6719b681b236b7f5083816cde83dc2575660bbe7e0bf37c6b4f570;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9f39c09a024b5eb0a3227610988fad158d2bb4eefed2cda5d87ab57a55a5b438e18f2c17dbfcc7eeb4e384fee426422b48038cc93b5ea411e311269ae228058430b5f0d7c6374dd11bd643cd8e9da3f3a8ad7432d04148a3be2556ac11c9dbb1ec18d6a09536a945f442619a81d709fdcda968366acff165700abef585be16d1d5203f5210db9dba447bdbf82771ea4629f485cb0c500f9acc0242e8c931971bcaf1e4d323877e67bc66ba8a9326333e9a1150818e3b2aaf22c2a844d4296c257325442b33fb78f77e4cd6033b4c6854339782018fec67b497eb372ad09dede29cf23b9e99a7673959e514e86c9c90d8eefecd2836749b0e2bc9f15f38ab986baf4737e1f6debfa35f9ff626d82e892e3bc718eafc22046b72ad27f869567f7d7b3370dc825d9d8bc236b55bff0feb9557d76cde83326e5ba43644ee295fbcae3340a03eb5c32a584b062eed219ee2085fdf995a196d393229bbeed60361631156e39def28233ffd1f07b243f060b61c4dd3953a698490835b029ce7afa55acc870190673e99c85b85b918e58073d3e52648b9a6e7a02d3b77338d6406fdbbb43b6cbda74ac85e963471a405d1d78a8b177a037d10351a541821e21ccbd984a171f653aac9e66bc148a113d885c198f485567f8c47637102db787d20ba497756df3c144ae5d7e4f5079aae1de3acdad2c41ad21aaffe8b7b37e13f84673ea95f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3e10a2b5b78766e80dee43544e0b814c6791f2456c0da888face8ce0736fab3f0bc02aac557b687808304a105465f1383ff0e0e321651bbfc3479e19e47471006b35450a449bfb19562f9d4595110027c02ec85ca5a70dc0047a908f73062b42dbaa16fd30791048bf2b9008b7a501cfa09a864c377f08d3afc81cd92e63ad9615fb9d4e35ba2a5708f979b64aeb67935f6efc1e9184fc88f0ac24a4ff18fdd524745ac17f38067a2f4a2ba0c7c45c50caa7746ebe87e8a7c5a79c531332497632d15d3f7fb72620931bf372868df5892daa1c077c41fca0e898b69db4b05c2f98a5e815863b8a5a6841b3266e466e4eb42a3a6c6b74ef1a8b46d1a715612b220be5fe9ae31c42205f83bc039f85a05944da767d53b58f041c0effb7ea79cd80604eb7796bf8c6f6f049f82289a2ba3f3fba321320378026e3c36816ad8056e8ad10b762c838321d6ac63303b601552193a64a78fb94c638c4787888a5b9eae09c098e3130f7eef7f0c861df1898a618c1f96ac9d98e4702d97aca62ab21e7a5182c567850237f27ec543d93a8a28917c9d4b0be5df94f33cbe803308a59df79f2e8c28552e3db5c01a877626f638285a54e5392450de63138e63cea7fdd72f709ebbceedae637c0a1ac9925fbeee3121fe04d4cdcd9703654917ab5c0974729180891db3374e65de7579b79423384f9dbc6ddb5bf0d7667be4e51add7966542;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5693c657399ec0c47a92ff0a2397613e6f6e910615abf9ab2143fed37ed69d89361d7bac582353ce8537f3cca6ce777c1c06cb994b21f684641ab1a75cb1e182728e19d0d967e4941a3c83debadf54d39a60310ca9ec4e9f68f9c449bf479d2ab6b97caa61c4397a7e9e7bdb1df4d1aa097686bbb92d13018541a84248a0cb0c83bcf1bd81b5c8052a93242edb000d83559a77b417996d96a40a3daa9913a301aec2c14ba1d9f9b46c5d6a08f9c057c3395521235d9348c33aa9711d4248776ca576bbfd31b84a2452126950acbdc779cbc471b63ba13f9e293e3057d461553b987eb4e564cdfa4ce5640f2330946a8cd42110dbe2085c106e42150104c9beb57531548a2daf5353e26f68315a31b81f67de687cc432a2491a7382f2fe5851039301f4713fbbf5a3107e658267f8c36b9ea3a1864137204cf70257d507e834339544de12f8e08763523c908b2e898e64e3c5a2711371dbe7241b44c02ddba8a9e4607e88fc5feb7d98b0baf66974142eda4cb97d0e460094c3c55f4b6d5ad3fbbf26533ec8074050bb15d109746ccd95c1f14c20dc12215fd3e8d707d8a534bba3af447e7753bceb704e3014bdc94c9f84151e7df9591d44ae751b16ffa4c9f0dd719c2fc2047910025388c8fe4c5596d969b845323c341b9ab1e3d29a1137f34b6bbf2f66d8ce1fcd3685e27965d5ff4331a7ca6ed5b66219c7085785995141;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h54986c27ee12ff79e641f2363d366e58060467cbfb7cbfdfb4f0d7c736199482de8118b0b732a017524838a2f92f155e5637c22f0c0b9fd15d94d9f4b60ba23f62471ed536faac469d7dc9ff306c89711cc98652bdbb69053d5598784c99014bcb088dba3d2ee943657cc68064932df6775c7e18dfbfe53aa3760fb0e5c7e5d0f6771a3874b74680dcf138740a35dd70ea131ad11c410a9847da8f2dda5c6fd5aa8d3615a3ac44eb89316119f4044f4ebb9e53fe8004cfc393ca89353a4919323372e93afeac67d7b7ab55d3b20c2a49101d5bc7a0fbcc5a4d2de6ed0701f282cdb50c2db460b46a2da27c5b3747f8ebe3ffed845f7886f087d190b125b11efa18365de0ae8e5fc66ed9b55139ab9527d282dd05c1029086c8cd6244162645981060e682c8e2b988cbc8048b9585e291edb27c8e94b6a7d2d48baf98d6f3bccf874e05388e796923735337190bc67f4a465d89b568647bcbddddbe221fc404c273b3f117dee2006a9996fbd8e9f27016b6cc4e77bebc805cafe057d6140dedc73427f00c89c45ada12ad4e84683c611634025fd4cfe4beb1cf997364b679d0032606121342868f4c5650936a0134bd39952ba032585354ba9b79c9c314c92aa450927f0e2156bf0213bcebd004f60e09da52d38fc0653f03207ec36e4fb6d4c0354c2a34f4e4f1114399ce060dffa4dd99c737acecbc315038aca93721fd340b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfc7077da453e3300ecac7b3ab4e9912eef60339426d2722de5552d566c8ecaa9a343ff9e05b122d6cc32f1b2bec5945850e764eb8cf2cda070ed259da9d7611d3c5492ec79672e5350a6376a090da794c146e999fa11d67c6ea03d1eaf2f80d0a89ea1d462f54c35da4275d45a1e7f537fdbe5bfb74b8285428a5711db14884e313fe1b3c9a57fe5212e60ac0db622b86e97a5e351c6397d8c739c049c4e8902eb171f784624a0ba7a5b5258211fa47f2d1d80e7b50476925b568a791c5f4d6ec4ada50595328d20ba5153acfe34fe93f1abb34feec18a7c18d3462a4887dc91aaed94a6d348a2d170cbb461cad919e36f45670f7a9600686fa67fabd441244e4e2a5ac524f53cf34d530c799bba043c315c9de1d9d9f7f8256011bc7e6405e0bd04b1f94c6a04c5aa81ba8adc968d3b14ac6af6e0b31deeced6994bb84bee8a659f022e1f4a74fc593d8d2902f34205cdf8c11c9f3c90c75d2548521114e3929c77502c1078e0a89a3f51159a0ecd5251f00325bff76805e28d579037594a353f721553e5eab5776b592325b3ac34eab965905c23c74a4388a77cf1490dfd740aa6e5a9393a49549467a7a264acef9e5e78efb6252e85b4b6d13a45f5e811ed466ac99d6ad234fd7dd5a7b152a7350c3bfd95dd4db8e798799dfb41a9bbd0052021900a71263b458b910e6d3793dea5fe1a41535e33f18ae46045364bbf63dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb6d9afb33728917b781f3c593ca0fd8bfb04745ad909150919337fc996684d5b023564654243153d2ba6f958f00e9eb0500ce5f8a48ee5c9c45864ff92b0c13dde7ae1a12eaf2f1f6564a63497a19dd114779f969d4fd36d4857e38502bc846743f38669151b234c3183ce4dfc2fc302f5dc1716ac80151e3ccabc3eaeed36dc26c81b2809ac3fecb3a3855890339f655cb6735c53e3025034e9ba75f13d9acba502ff60e0621a84b59dea85ad031dd134732f9c73235231b3479e92075003c2624ae4cbef5d751c8fd34889dd4b2500f178e8b8459d09c4a93bab73ce47dc2c97fd694de2fce4d9eb424b6a5843a361f82f60d1bef6e71ae984c05c0c70562493dbe1e1a1652c946aeb4b32bc60a58c372a2fb4ce55d272a45c578afb09b987bce0f2a6fe77b22c064eb8034cde2d767eae088fa6bce135319c2f3a97f22bd3c1204f478ad2a4e0311e989b23f4bb1749f619e22d12435e10f239ecaa88e295b72a3e20f3f21b8a5f26867a8fbe822b3d03cc026877563a058d33730d6fe49c1867e18db77f0f6dc9d174ef6d788b9cd441174e02f4e2fbad2caf8289c2c2cf96442263db31683403112395ffbd3a7039c95ac64836f89aedb7aac8e9be1fbda6fb50c6586374315f3036baa160dfaf027331300756bb4234a180d8e41aef65b8c91567cb2af451625c008463d46eb89031689a4b62648ac6700e8032af6220;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h11f3941408490c6ceb81906959f0b3bd34a8aee1e1c67092731a355f2d804fc7b1e545b23d701c8eeeb5ac140838242846525fae86416e315bbb018232a5b9f0701f86207bb1e1fcbf72268f7725b1d0745813dc8225de33bd54a13929a876294a43c69deb7e79f66a09063afab2739736961c7163feef234fed29ac6688ff51d5e273143c26e7654bf2d9c4631820c8ccb1e916bf5b743425e426f31eb7bfc74dada6fea2fe19516ed3c34207bad6e6459ab7f9ca358654b7513b1da3e365899737e9066629832336d9981c5098da8d4073d86eafa942a78c38f23329404516eeecdbb5fd3010d403346a078fa03b83b6b707154f0f89c5e7ca40cdff7097a9211a796d1b220f12b8c08b87c26b44b902c92362db9f546c5415cf47b82161b7b2240d16dd0589cf8c55ee107a2603378e9b065119f7d6c20ee6d178a0fe3148f7fc9fb0c7025d3439da28f8ae302b2f88a067f87135e57268d9e89fcbaeb06e9dc3a0f6e64819bfe1cccfbe503df5bdcb149c8bae4d3a814f29536c015c596af654dd59564a1936ec60d427699180c22a5f42c3d803f1ffb1cf99c5b437cc22dfb59c408aef865747e81920460f283662f03f1d0cdce34e776a2b735d96cc7f2dbecb80b9c4d75a6835397e7a536947855dddb8c1673938717cdabd308858e0ffc220efefdb4c4b117035acbd2247333fadc795d5e49935ef5bdced37d8d9e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd32badef8c9fcd951998c0c413d8c1f8865c87aae87643b8c0d969b6c889aee5d112e50ca99b96c2fafe8bac0d6b5830f55dce0bf47bffccf9acac021eb9bdc8f7cb5228b876a6adf2bd32c3bb0410372d7739a68a874470a88c69fcd14f3cd0ef8c530926a3e15028ffe1e4a5ed50fee37dbe59f768b102fbfb16c2ed197e27010286e9681fc89308e4a6825850536fcf4aa6d88e2e05d944553ebf3adc46a36e60142c356f31963cdde07de98e85248a1d4cbb939214322d8d38079a5583ae234e1648bd4eeb9e64e9146db4354bacbe65b1516a2e0d0bacb1a03fa6848eeb8361d1762111ad9eb124a063a55930ba45ab74f9f9b6f1406bd4a449979bd43549a62e4da57f5d41327aed3bfcfe5c2f79cd0ff80bf55662da459b6679d42c22a7399b0e487c33514d2ffa3a5a280a71846b29f946b70acf791f06b8071ceda779d7d2ae8013282d0050843b17320574344cbc527109a67d51785a1c29a490e050db06e3df24fa95240654ab72e8f6ca17d558a94f8438dd5f0c1736acab12ac959506d473ba07d75ace121f21b476ac74ce1d094c4400bc86d9790fa9e35ff8237d41c8f85bf59bbd9ad5b679f04d318ef28f85cf227dccf4624c434aa502cfdf194745cf3d9aa60fb3f0e4da79e371b2b153219cf7df8f4e38447beaba1dd1efe790581036cc726785710667dbcc10334c157ce0a6b1b76a92942afe381be5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2c826b1066b64b98e66cd6672aacf4ebae9304b53e1fe69d33768a802966ef0643fab8b5529fc8498fd1e9514aa542ace8d52fa50339848c47b0a7f3e7f7fdc120ecdba5402648fe64156a1b88fc15f788379d620393c6beb62b46818aef1f6afe4086766680174c18f70ab48f79d3cccb6816959220ddefd1cd075094c89d4e910ab3aa15e12a45a06f013356c9317e8d544bac8c6bf737d8a46032ad010f470e64a463db7e264d6986f5eabf54a99397f381cf65d2bf5526bb7087174d15b000965ade32d2440df6f58989e09541cd419c81c4710b18e2d6b8c2134bba01254185abb25b774fcf358d5bb2a3f66eaf59617a08e7e3a5ae2ba63384e3139fb8e57f939daa44eefc418485bf40d2666e29f4e3805ada75097e88645fbf080228d1c8f70063bce5169ed45e6f51e31b013b1ecad8d39ce976d73557bbaaeb8db07125b340d835960408c2923d9c04241c4daa5886a5c2f02bb4963704dae73dd0d5952962e082a24a325b31a6691ab1b96a1360b9f979a35436e4c6905655efd8cb02fb8f61f3300d539dd723b8f73ac5c3b4efd09dbc3961637caa84eccfbff2a567d6ad660facd3e435904be92d043886233a7a2139fca48541efffe585c4f59a6e406beedce9d87bd461ba2bff90d37e3d3de9f59ae1b756f49bbfc312054d368aedb63c00d48dec2bf1b38f130053e3b8b29015c0df8df9bf54d2df15b004;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd82e32c0b036bfaf53e76e069ee6b825d8c83749db2c52b642d676156ddae31d7847442501a5cfcc494f512a867f6f8d53335cdbf469fd2d3e2f0ef6f73b122188375724208011c765c7c1f72ead8df43acee27da2ede6de52fec5ce465344af18aeb7377487a70cc2c5ca12b9c7f0b441cec9f03cb5e631b505c7ba2abab59195182153b8496be73f9c385497796f7ca6a1ab5b7fbd490a202e475621e6a0c2d3dcb57f928152df80c41531d4c95e93cc998df607c975589ef9df4c840b60b400a060ed63058651f93d23fdb5356d6d72dbd838bdcec46d3b37ce0d841b86de8a85a27849c22f6d568233d964333d4bafa359030e1de7fb55063fe4a9c8a4a1aefef1549070979483815dd0128609f233a94246c97683696c110cdd12debf9ea1f3474123d39e2d7c85293740393c17850a6f0a5f739294b365860a8f8b9f591f2349337af53eea41ae5486e75c5b474c128441282dab8e90fe6851fa0d4fe84fb7f8a96c74ede397028e3b24dcc52bd8c4d195967bc86d551eca51c12ba4b07680b95d64d574390def1ffbeb1db6e432b9e57ee27ed598dc6f97f60e18398eed43d5131170ed02cc48c0215b8faef4f55aa9cf7bd09a039b2501514c6d9e359d10f99945406d9052d095eaae9e972bdeb787bd1d0255be1cee2d5daf8b37851c3b692fc3636c19b00e07b5338f22814afbfc4d53f5923c19479dbcb2a50a2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6cd003670ed2014e76f3b810e8f41167fdc563d8101e47b8225c27c8faa9efc4fb02f7930e7a5c3ed5ec885bde2ee88db19ec457b9c41c596ddfe67d2bc412c9988faf8050a88450a56ede6d8543ecf3016e64f4c522f258116e8a38376ec64b88c48d28618747920e901993e2be8a42c4fa82186aab180cfb10f0f1d4954bca1cf9609345afa30e26f6d3c0f51e4ca31d944982143ab5db47b6b26db587ef39eb8115b10a3f3876c35cad57d0100342de9e2f2de66128aa7c14c07a25a14973b1d1699c43a8bdb0189fc9d62eaf73129ac82d27e19971571ef717a13c6a3cb602cfb687b05c856a4e3138af63219fd3b92d7d4b48d5061d92f9ffd2aa86890758f07739ae429db08040b59cc2ec363786301c4077de9a2ee415822762b808f182872d842370afb79da1f2dd59c0e39ba86df4ad3c07ccb6b04a63e1fb9313ac3c9713c1ac6839d6d36cd6decc3ccf3fdae66247cd0b772a26ba9d2ee781c45c5baa873c5235f75f7ba65404b7853dcbaef28de4068c5f6577bb64947ec23fea796237b4cdee5c8c180432c9fbec97cb5c9ec53f993da62ca5d35ad9749b5d371b3951102b76527256ff5ac905de30ac00c46201d5161ee834110e32868e15d8c0629408421374223e7dbda301c51107ac086f51bb674392695187f785de80a9ad81c3ce08bf47fe6ee0e1a19487eaf675efd255d14f57ac70039934ecb4611e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8bf54ed3dab430889003055302c0ccbe89c8c06cd36fcc4bdd95cc4f131fe5ec7e0d368b4c22091c2aee6d1b5e3f4a989c0e9f03dbff9f149196d98acd352f1173513d9b7b084aa3ef8c5effdefd3c33ed82597f57dcab4fc64fdc4056d4cadb39b5f439a6e031861cf3c9377b56419b8fb7231cb80d5fa31578f9abaaea5318f56029665bb276807d11ab45ecdad5ddd9708097c1272d4c572e097382361478df555d507debae4f88b68e9319679d93b1e8b27bfbb1317095b3c1c5dd000bbd45baaad5ec58a9cd72c4324d39bcec4f6ddba8b127e6b73119acbc2fab99238571c08fc1419d220a777ef7cedb1eef7c79aa557a452bea4d37612d6d629e7dc5ee707adb89f93e492c791733d3b77832d1a22ce022ce485f1d388c198c55b2c0aebdff85d645ba4d39069d59a94651670e6fa7a6a702a711039be59e800e330ae3f5a38872bf35e8b7d8d48a6f20c68c987b4916eb2f4638d5c917b6bde2dfccc370c793bd779bf5c163f1f7cc9cf04980f2eca8d3f6210ecebfe8739b2702e50ce6e23a89653c366326daa197105bbe6f0a069fba269d623b59d51887dd45b0f0cf982dbdfd11f850dabb8e46f7ceaa8e9882b3013bea9f61bb0696311e7beac095ef9dfc6332e5bd2ade3412ef8abeb147d14ecbc0ea09d12e0446dbbe27b08cb41ac53291438cb964536f59104fdf6749437a8b73b1d46b65c7fc73665352;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hee0b5874f0809ad1e3137119c40f13dd16d06851b81c20113f3c185ad181d8a63c0aad4f3e69fdfb24123ca413b1dfe13bd2dd2c413a751d218ae2db0bdef19109535f329817149523c557ca2c3cf67aaedb6c18e19340eab13ed8d3499073f3db17208c2d95828b2d010652c58cf79df6aa7f9c8182aa659d3db07cad7990878e47c9a618c77b69d79e1721863c1130c75d62c15044d56cb12cc12fea76f767827dc684caa03eecbbd7d59546335e21fe28432472472bd629d9e610de2228b172d9ced39cdb6bea6c18336dd1f9531200624ff15804baec9f561e06f5c5e8b24f55d77ff4ae504668c26d424e23d02ffa8c9587f13ea630c98464be9b2b1e3dbc34ad2d054d32b87fd70fc7f129f1d1acf0e2ed83d88cbfb714fdc4928a663b6323abae99de4e3d4ee98861634af9ca3df0367ec98e8fef331b6c5b48d7418739a2239b167cc983921a648e47cd799f93a6ffd70980369aa1631193eac3f277a79df1aca85c3ae23ef3ffb911a5e62fa0c766c1589758e5da99bbb44427a7bbcd62b24bc28102382442d74960e5ff705801fa57493adf5559f5306c3408fc25859dc7fd6f8e397ce7381e0e0aff6ba63dd3a4f5afede63eac9f97eda5c932fb961cde584b0d36c9c0ae7d3114a5e424e9e89e1447572a3e6488fcf1dc88bd5c4527e04a97a4523a5a61d72871f80b24343c751149c7cec4818c53fc984549ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h661eecfaa83065045a5f92f1cb6aebe38542097a92d601b9886532cf9a43fc55f4accf18bdf0012a4eb3a04167fda6e737db9baa5b8e7b3b7b7ec2fed3036d2245ca6631df316cb57d35239eed8bdd6128d6647867aa3d15465841d9a9f73dfbbd1c912d9ead2364ba5ee44e4369c1c8f16ee19382d2c92cedb2f202e3d7a28b3fdb5b3eaa66845acb45ba9868cc43a3e78db9fb81e8c61d9afbe4113b1bee4df5f3e04bc9efbb59a994a03712c23b00aab34edb39e6353978b68b41df921c037bad437d1b55e5eac5841928c92dd3d80af606d8a7d84b48179a54fb1e2d4fb2abaced3f05bb6ab819a49e07f947b95c2cfcd7748d89ca477821b0402794eec05c24c5be0975b6c6ae9c1c719dbc86297d600adbddf7433ee1b617ed65e0deb26622cb6dcff6751370eb0e179ccb8b4074966464281bda5193cd250132b38ff16a4eed9160cc74c8eb8a4949da129154d632d3ba4e811f6348888a1cc48cbf7d24ab075b905c79d28a387854d4a03bd1d82feef13dc08856adeda6eba5cb91852181aac1d01226379d61ad51c2c19dc4a33359284351f939d47eaf3b4d7d8bbec6bf37f36bf17cc81040859c62e813e8f8bbf824106ac4b3553180fb09c200a5d6041015044d5b1b9a0a05b1d34aff23751d56840e665b209f9dda45eccb3b1702d26648389fc20aa5f7bafa009e3181eb3f520005a36597c4542cf6d350c0c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf078c4d35a2359c0adec4f100cc073be2b06f0c9fb3426ba971be8584e7f04958a4d32ab9eabbd6befa2c81c67ad71e4b850aa06e2e5456bcaa6597d971e08ca32d819ca8940d1287698903e0d51c8368cd18846b859c868c0ee43e0709bfe72ffd0548dceff5236ae05375f858d7ffab3b80504eaaa861435e0eeac55aade70030cd3fb6a8925e4865505a3eeb473c6d225a163905388d6cf759dbac4c59c0c26d71b4d031c1c3ebcf0a1af9a1fe5368e499602d8654bede4431639d2b527c59d92d8f43b6d89a7ab1006b31c5a248c6b936dca15b22dd751fc6a5d5f50b89ed11d6273f9083e1f90996dec777772a8d7f3ebad9464bb8bf36c10d898ddc66ee5e6730c54b5d512b93219f32a915f546dac85015dd108f1f70c90eadd6921cf4263c41808994b4de84ed76f70e4645e386e79b2f0214e74f18fe4a0f3df668991747d8706affb248bbc58e2efc767dc4a70bf53eeab5771437fcdfe7dd9fe8cd8d7c1abf9f3dc81989888df60508a3b0327fb9e9c7be163fd9fe500167b1c04d5a8dc67bb5a41fa1e18ec313d77813312d5c4436d9e59765ce92cff0c52dea197cf3325067bc1662e8525fecf9f22d2a5a331d23a0467b030de54217fadc4b098020e4e11653ca8d3510b0a3aedffaad41a4d7064b52af7d5323820a55f102eda78e039824f992ca92067b07193a45940383c9275e274382eb42b10ab7288c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hbeb5474ed48ba907c105f90f0a897f6d11afc51098accc380cfcec2a8ee77fe1d08c93cc48e071871fb02fffe521da0393dd0e2438bf7dc607d5f5fd8301c4ccba408358643bf745bafcc6d391300dd690b21aad59f08588afe1af96bb28663b9fdd637e9b3a6c905a37aa1aaab3a6586cebfa0854facba3c205eb4f8ff60d51dca0b71a79eda54f7e7fc1c6a55fa82afbf0477a5b035b92f2778edc576550238c788a59e38d0ca84a6e8ba165d2d6ae4d10432f36854e66008528ec15e8f859bb70374bcf8c55db03b13b42df296e7999bf67afda5b920646db19de5ccea07d525c0ad5e0c4d5d212366b607d4f1a2568e788f5de55d94739497b1e4f44edbad680b33e654a64cdaffec655576244091595994be97da8bac7d7195ec76acfbec2073cbeb1e9cb9e9f9523f3fe05a7b99315d92563fe3a962bede043e0721ac9f8a9597db3f206ec80e9b9cd3f46df1e50b1f464fbdf86402f344529aa32f49231b2c8930ebd65094b44b2fa48dfdd74b86a9f98300f50db5c66a34e1919ebb0671e60b1ef4dc1e538ab03ceff00e93ac84aea8c943bb31361052f31f78c77425d8e151590e6407204da20cbaf370bf2aa7789e4ff696f1a75432a6cd15c6223ccfcf5594517b95719458a0e1c7cd858f9afde750d290601b4c84107393eacc71c669dae033cf0fd60c838aaae65cfd525a3bfd881f2d1aa9df2af13a0a6a335;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h138caaaf17b43162b6dc0634b6e7086d743a01a84c5ab8413528b2ce126135dd853d993d5f78d800b4fe00e6a0649800a3beea45a67891d6043076ca96d247d2be7a6f2d2529c090edaf259e26bed4da41c073af13f4dbb384153a049c78fd36bcf7223002c383c31528f80d0dff22abb9ad2e96d9e1a9e7fa23df31e136c924bb66a2d5f45f82a056850df5414ba6108ae08c5de0c507474806a8fd0155bc97d4a36b083ac125445794400aee5e20e05693c5ccedc94211290bd915db0ae324b173ae485aa5224d2a42c0fd83f8523a78c6d47031b1a3949f9c3cca3de65f69529360ec1a6dfff30c1271956d0981b3c19cb7e51f424b6c3338a36623f498fd17802058086c7b1d14a141c5bc99737729a6d8138a17e5b57dc54535af8db98cef4db511b8f442c27a432b6a41e4f3dbe0cc54fbfcaf5cf967ecf278a159441284a3fcca307c90b80beb31a79419ba01ac2475bcebca110e82d09a95a09ccb0d907476cdf61df42073e9d23c906fd4617dcd39ee081151d36e996d9cc3c4a7692cbf511e10f5b87f24db9305cd496d1021486477d20474114f4d048dc2a7f8bdc3184567edf9d21c7467e6ff6110e8c967806368b244ad67ffa4dddcc2db02e6991cd554daca5a70d31f3543ba26e14d46df045043f235efde4b34d3e36719e37cffe4613995b9142bca31b28956b558d3b29aa78653db55a152f26273d1948b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h79b559f2833d266e896ad4a510a2ed6bfcc9337294e4cdfed1ef29ea17e9a7808a880feda6cfbfbd9dbf7a52490cc0af14d5be0e40752abdb721fc03f5a123de7ebd57398b037b986eb6a298df8d62eaf784a1b01c2314686d745c208aba84baf238c1efa9b32643d8c0a76912cce0af05ab72b49449257e2d9715d25a47b506d60110df5ab33748ae33c978c9b057964e8b9a27f512066ca7032f399646d2c03d6263fb6768c87c2388446d51b3fcafb958f4bc021b76a4c512b2ca8602cbac1c541466fdf6c95152098cdd1b9601de301407a2413801b1b51cb949ad3eeb5e9569f6b0c2f0d216957c7d3d1da59a1488e08137f4cdaec68b8b32836aaf0538994da64790a729358a0ef7ad78b814e450ffdd8b665621561c28eb45499ef5abb2e7c82696b79eb787ff0ff053d07c99ed5c1251ccaa15a2e300d1f6cc1bf6f2af75b842d8988d59b72f567c198683ee2a8c17fe983587a3cb4fece240419313a464bcf598417b22b7f5b714360b085471aed5fa258e1d372c3660f503b354d8dd6b8067fc5c753b675a0536ba7748a98d94d0f3b7217a4e1f695deab9e59dd5cf71d629d14e5847eb91da21b43a539f5400bc5997f58079a2badef59b35c97ef6f2cdddbb71328a717340b74dfe2f67916cf2a74072556ea22870a168cf230d3ca63dacf8c1f9dd2f36e7c49c956d876e33a52950b8c96476e649f357c5fd07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5488d1c1e9b8ebaf81d7116427752781f03496e8bcb5a1de6e040cb718ac030f12cea52edd47bab337db13b24097acd63a209d51adf2769215d82ef3132018ac2e37dc55ea5401b670432d60895e3a070aef937e00f9f0b5e577b7ef3b0e8d536b1491c241de0fd674ed3d00b4283296880d7ec888494c07e3524e5f6545fa31c2c3c379c57c8a9ac6156c9a0cf69dd3b6aae2eeea1cf8fd135b039d4117f56ab3a7686fa03060d5af9db4c425df3d66103b52baa47d94143181f23198b6bf19123da1b661bc50fa38b6886f0763d03c9b72a51a3cbe1043043c5aefbd6705576a763b71338ec386b40720cb5ac966f028c81cb020c31bd59c898e86553b64071aa271cdafcc4329a4c60f3adde9c000d89d4bae477642a26937a654f48b0d25758796d146d989dc32646aa02011ccc8e809a09d16c6045c90055a27cdc4c681210324909e6c2cdd8057a81d056af92a6bbf0a292f4ef10a4fc3c94027c3822c41eecbd1c2d99b2d02027d30dc83887954af84de0d20625f66d92e403a70ba1f5bf2891a482e5b898145f08ecfcb74ffd67eb9e94ea082e8580ab462d439532a81b9706a2e9aaef141b8155d396e68a36293346c021f1c9547897330362e87f338a2423e5898c039bb5311f6bb07f93082908144c9e20d5af911651db633feb5fb48a10644f3aba70985a03d47431992e7d92589f6b7f8950042476afff74776;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h58c78ecb2caf54b02fe9944cbcebf9a3675fbff2e94812d0a5115c53b1f94a9d05f534e98289d2f029467e15acc119893eb61bcb5e59a1ea7049727c6ea7859a9ed0c00155190a44c0d372388bca9d1f30f9afdaecddc99f06ea3e996bd5403446f5be67514ba4309e83867db2f53bbcd0c7ee5791a9999805e6eb9acc51574fc436fe3e9ebaf8da010fc6c75b225a505f636fb3f72698159c028e1e264f54308ec23fc4fbae65daf75f61128778e9dc7e24c27e0a3b19ec21aa6b2599839ea249a65739ffc915badb48f3231d02b24284b4bb98e94c9221f823f29a50ee91ca8e6705f263a7f731f5b9f589ff39b977b9aaf94f3b75789a8d2027c110cab3fbb9406da35de2f67074ae46bc36ff3a594b9c61df0dc4f80e4234841090d878c682574453da8792c5478c3afe79d288540855fe336c07664905012bc894225d1f9cb90fc86c104441a5fa8cbd86484cf682fe0d949bf507bf784bea86c61369bcaa6f0a6a9ebf1d3bee0ac37b0e397a82a5a4d4af6fb70726e277070eb3d6b9755bee434137ed43c2c87f240c3667eb76f91009e0010157544eee0e9ee6ef7378bed3a8b4f2c95b97e70e26bc8a87d9bfaea4c738c4af03358207431c808db8aa0d7d3690579df2f53c313648f0e314b4a6a9f5ce7385db5be5b0f451c95b4f8c8fee0e1e1bdfd20b7f72c564df182eb96777aa3fc787e62c7627cd38e782a2a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h15df0a9e8b8ee7874f2a579121393a222285ac4b65069216a18e1cd47b5e92a0e7656a0373a40feb1627378ce5f622726419118456d4a7604713d71a37a1a6ddc2904b052c14252e60ae14cb7875353ef4d07259677e9971cf58c0aa8d625c8ed231278c4c808f4b1b3cd2c34129ca6d5a62edc06148524c7844ceb369b8d7ba8eae3b2449bbb062d9de373c064c1da3f07bcb80b478db01ba93bbb960b5fc7697cf8dbdaf021ff1d1ceefdb1111bbe4814d88ad88d00eb102887839349e3f165d63adb4a5ec9247b2bc44f459625714dadcbd9564b2cb93711240ee507534ca5cc76500caf47b041d16d79de87a68d2143c43eade90de7237371657373ca973b5b31d4ed96aaed56336b4c84527e830f4c967cac15c978f0d7488f8592e91dc40418d4b073f59fb2d7163cb32b976de03854967ed284ae3918b3802b910f75ab6acb742a2bf286b4170ac264de7c36f85d5a2ab1108d5cb2e9b81b3fe1a6b779937262526b0d2ac26a0b9724dc347b1af5070770a73f62111325edad7dc1283d182012be1995b3fb7a1654703511b07511ccf1e159f4a5b456c5e10f9391da620216c2f427cee45d64b09ccfdfee9d9583378d79859b42acfe206dafdbf22ce531c651b46a27380186c534c2cc0be4a4e3df13bba1d09df8135cfdf73c9ab7fbd4fa24f495762077b91a7efc6f4b949bb63a54df5e67e704b4eff08d2126ef6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h161d0785ca9d78c81f934827ad5d0e667c0391a0c2797796b6dc2dec92e3b36345d47ba46f54150533b9c1e80f0bab2cf645354c6beb8dae91bbbb1ac9b3620a3b5eba0d395237a5bb1a8ec08afa80447b36eb43d2a3fddc6cbf192130660257641ee08ce1c485f4ef84f3f76f284a043cd5e1079aad341c795e83af86e7c3f9a2231387ecf93f3077ab3c356613ae19597933be102bd36476bc7a0b923c6d1daccb4d7f754929e15993a5990877dbcb50e404f4acc350cecd1aee57c6425fc994d08eb14ac4f5915ce5c8a9495aff42f75fd0c86e346e1c9f97536a5a44e26275199626f003ea40d0cdbfa8e9f33383bf39a196d99900d57556c3bbc3f769aa2eaf16851d18628c299ef025603befe869f3794d6588609e7ff28d0f7a2133e24225cf49b1afedc27fd33507e78dd9a4b707c38dffe48c93e575a0998f3e1acfacf4b8fb9e2c80cc098994b5042f00caf302ec7be260badf8a3eaa2861118fb828cbfec961902acf35a02a380b26911a2f8fad3b58e2ca9367fe3ea09b51ddc493b3ccadb1e016240d760db70bcf63e6dbe624655eaa85c486010be40942c1e9cd95bc398b4e25f63483dc4c41a04c864b80bc035a837f95551c952867443b726fb3ae5d84e8b58f3d7ed02a9373ecee8cd529b590e884ef23011a6c3f5851ab515b609f95ddaa53b3e5dfa3dfc582d8e5007f6678b7f11ac682401d40e7ffa0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc895c752f1542aca2d95b501f07c27ba562a4cd5b3ca9422026f09c3fe898f0730b32907bdbe6af60b69cc1b47e7f938ea80c50a5463c1c27618e3d4bdd2d63a3992c8ddd75800bb1a4e32d1b6deb4c35e4694c8eae73b2f487b8b5add1f74c22d7fd21552ae66ed3f740ae6808bf14137c0e72f065004afaf1cb3be25048562b58fbc66e0988a5902685d69d765cd967701c988470ec518aae9fbf819a5993828408eb004b125548d0f05b1f118117107981202612e7de6bd971b270f0352e9a84203540f3cbf14254d875bfa45750df19ac46d3a3d8b67132912467fbd57130b52f0340fe48b0b042184cc2759886d4b1a85a51e137106b4eb8207f20ae1764607d5d42ae381560b512b6e899e6009fa138c72c4103b78cee904571b30d00031e66647122349b7d072c7cb6b0e0931568f1b19e6e7d9dd0cae989024591541494f93de721f76f7480a45fcfcd3716da24d82b270163f9bc22dcddcd296213da2acaf08fa22bc0aae47bd5d49519f17f45d9f34cb28d42dc21b88c84de9301e0f8856ee62ac0e9e87fa3ddb50e9182a498576b158f02442779da2101e02f3597cf1dccbe042b24ec31177e049fc2243389b52fce2ba0764f2bb0f31692bc8efd819a1381d3f69e59e9699708ffa7881a0f6ca806dd523ed3b74f1b50ef9ad349aafb39abe9667788a26598550df987d65b333cf2420ba36a10b5d9ac82ebb32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6ec44547c4914bd02a137f033956bb73c1779c73eb3656b30430fbefc339e5fbd882a2709f781ef141918b12086eae9898c95a62c62b60a1c7f1df22ca8de04c4f6c013d71ccc7863a85add8bda435dcf734265563f635ebbe05b0c04ef0cec3bb704dca0fb46955a7932792e123f9a0b8759444d461338c52c728980eb2b2affc7dbcd1f5143da761c7d2d43c8eb62bfa84c242c38c5053d2272dee9f4876394653bb586bced2ed7c447b7451435472151ed2f2a7da76426ae362e12dc145d9787e7e79a5751d20a94fe86f4f879c1ee95cbd7780f2084a378f473d61c389958929473a3f12b080f63f8772ba20f57deb84058cb31353f5fe72b30cf037a084df3ea52c23477cd8ebb75ce4aa0e68fa7b793763730e8587b65c3b7c82b270854c97ee30ee2495c7c04cc1c946bce5be11486ebaa37834b009cdcbf64318170f182081423b48000dd7bec2b60c87e8a40af5378feb1a6be09ebbfae114c987df0cc55b3898f0bc1aba82a45b4864382c155158433db78233f5474df0ce500471ff1da8d2c919bff6e007b72887b4b7e02f39077fec1b5cdb71c6e3c02f86d4cac3df9e613afe9302718a3a99c4cd8a89f72056f6dd56b591f729c6235e0956ea7d282522fd135ecbf2602ae92d91ee2c1455977895c5c7cf5be67773d3e5315a93c4c619511917dff37ee601cbbe41189cc3bf5d3bdd076b6673d9543ae1c783;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h24a7d6101e9b4adf069656037e9ee05aa396f900e145afb4add89360b7e221560ed3763b7378e8261c12d6c3005b24cf81488b3242207bf4055bf6f22717fe0ff932ce946fd5f69fef9bb5619c3a3ba8f87e587224f5b107f489007e696f2270b3b835945823e5c92146af8023a9311daf51fc87e3265f40ece863f35207a8f78b415944922a23e0950a9a26c6d2f1882119b3307480aca2c8642265e9e3208695535ebdf396da3ced1b583859e68004ec6d1e367fd17e8472c22c7e93a094a44af74cd6edb9cbffff598f0eeabd9979c38571a611a88ec4f53ca604020b09cec09932056c5c1c34037b4ff22299bcb6c0334fb0f3bdb732bd0866c6d60d4797c56253baf3f2d6dfee0bff7b7a42ddda32a335b787a510ba89108c2ac391a4dacca117bd72b09eb12c1c2b21361c7afc5d457429ec5f5fb7aeecefca3c064ed977a4281708d1945afd6a4ef4fd9dc607505078b1683da694a9acf206632ca7ac76c4e201911c217fff8cfa6d8ba89265baa254b86db1b25ad0c386e02b90bae2e32c02ae7d8c42a8ec37bc20e3bffa8d39c847779889ed8961f34ecd41971e70a0fd27bd0debc86fc3b197717b1338fa301d0c29bf178246a24aacf113ba7daa4a8cc1778acc1a241e092cca027688eb7968350fe4515fb02310a2701dfb90781d1efd1b42815f451ef19313f39aa112bc4b4bd9752899b9b92f43b5c767fa71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc084a0fb6baa4270ed0eab9cc0e1572d67a683808ccabbbf581b8bd741641cffcbf67df9c7d467c246f381f14139c8d28f766089d438332730495154c9dd728449db8bea26a7ab4cfdd48e7b28ad19117cf50605cec1b0ec167bb576491a276a33481b5f73d03059b8c1e078f67093657593d08d2dbf9f9f4fcf94016bde2b2fcae943e9199647937c916bc8aec20a5701d917d90f8f7a1704664e389c9cccfb9e19b6203868a4cc6e96985ad34a6ec80a88345626d27f938c9956a11ca1716a684f7111e50960870736be9867a2f280c481bb408c4ecfbe4d4f1c1f6a00c33d33eae766ad9ccd5b232f31349efedad3f30a4ca0cfcfec7e96a8731099143d7728d1fb42ae3fe958ed575bf4442b2e024e78b124c0e1602b3bd9fa407fa295df6274cc249b021826d33eaf3d85c0c151143fbd4dbe9fd110e384cd15c383600799e5fa03a3f8f99a61296d36e18a5399a31a74448c8873d7236f03f1d3db46573bc0dee62956af1dd198e7e074db24612128b0712438a1af4e4ec90cb3a6c9d7174f04fd74ece3d01cd0a1654d415af4da92187bd06b9b383d12ab7bbe3eddc8d928155e3f23dd6a110a6baf9436cc2cb4eaa27fc757091725286a6d45d6526fa5b7325be324c222a06dfc6b26d3eae085302066c156a3bc6e9a1f21598a3fbc484333a1491ec0079ebaec9bffde363830611bc23c0dd485545eeb3b0509d894;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3f429be1fef67f88c6a118327f8348bae8a66ec0185005d67f49b263b687ea5febb18baea21fcb6a55bb35cb4ef5e43e732d71bf85ee4c64edad2f21d9dad7570473ae6284b60b22ed59d525638ba9637cde392422aa01afcb728f6a91b6efef8e90ac1e840b4f3746ffb89d3f85f8c5e4531e59f65fbc32d36af7bbbeefd9ed750cb2f99a6f5264d9eb463a505b50925e2731e42001b8f6183965b417432922e5acb0b4e533b8bb54aef85b1df8a1618daeb8e0397fb39b7690e172b1559d6a4d49dfeabde6db4f251a7ad34a8965c71071f73cc28bee9b8cfb6a997ce6b9024f924d702e8fdd4596c0716ddcc084746a24e311af2317d2bde674f14dbdec00f67a06d82b4205672da88f3699ff4a461684f6f4c8f06880f9369033345e0355fde452ab9a0cb0fb336d0a0491197d0f44e81812bc60c3e14d8024521974c0ef619f27094941f451524819c2bff7eb15d613b6be19cd1ac5e839e19036df8f15fed5f49d7b311f84cbbdfe31a79a94f3b50de531eaaee33ec83011a1510f2e6a0c4438a45bb3d67dbc92bbf144258fc88de7a73e8c35b919831bfe3eb3728414e87d87cf1d4eda84f64bf5aaa85e335369ee6fa784ec6f4aa39d73110ab36a5efa421592066c17cf82d4b29f02d7368493f96ce50f051510650e006471143f4087a776ba2ce25ab66da2711e648a70ef5126eb9a80d394878b14ae8979814fe1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'heda051c5b1056317fe6f25e8446ec1d9fa4608c0c8358da809ba38c306eb937b39a9277c986fd5eab329f46e26c7fff88f8bbecb4f902f3ae160a46bf9d87e0c3659906db2b89cb561566626140afffd180571e6aa4b080a1d7433433053002f70c8ea3b0be8188ea2e2786ad8009b5a2709bdbd52988e3cdd1dc6e717fad7b3da2e4f9d3dbf75904e05496b4736f8d3e07ca90f3495feb8f10d6298bb2131bf7c8eef04c85d3561b24bd1677e39a26763326b34fc5f4ac1d6df51e28afa2460090efaad737de6de1c4729f9a1fd7de84cec261a1a09adc653aed2ea6a45ce1e97b298221abc17da34f1af6a1adcccf2b2ff6d6d13f3a22b44f402dfce5bfb00db3fae0f2fa50dd71e7cb8cd7b44014dde91aeb552c03e2c416d7e15d96c438c1d8b6af9ee3aa7dcffe49dcc5129e3166a939a052381f4d96bded7508e37846498c83c923e7aa203c43f94b4ee3f8d487b248532fce0ca95c8bf9de5c31ee6cbd2161c5f388ebe926d4e51587235dc355357b3311f439bc735c86517768897e3f0052a25bc7d39776dd64fb93d03664590a220ecb70e0218036ebcaf5e727db0df58f0f9c50e4665e60a5fd9152f03a77795a46a9a6d37dae68739828b1d53356a512a9b0ed5576205af29c2f73bf2a6f130cd92f798bffb455ab786d7f655b9150c7b94a39a1d89a2e205262784b9cf367ca65b6a6c9b7c1d940f44d5815b56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h43b8092fd564eba8be880905a98335ad92ab676275ae3b6d4b2eb72e949e13aa47f1febfac27fd9f35b1dd51d19e2c2c2cc440143f64bda066b0e5c8f52037bf6cd4fa46161fd6c02114a89017ea711e8c2aa041e374c6aed785e29294a918888ea0539929f16c98481dccb76882d6c1b4886ae249df86dbc006009c2879068f20a2e61836aa03eb135945d09059bc1876d983fe6671d437b63a9c33af4d7262a17648f475fd37ec850fd7f405cc4428a5b11c8d05aa520570d88373314db29521c7be880c175e9b5eb1a1ff7a747c16cbc15188c766cdd40ebd1e3289e33b3fbaa1d700e169846483127ddf95a1d826cc81aaab28d1408b120eb6810d2620d09e462c95f2dacc3e8aba80aca3df59dadf7f80aa6abfcc3c1aa329c8448e010b60ef05c28e87ade64a50084dfd2ecf362570e69d83c1264106f9dfb09d1dbd2703244c3793b7b732ea63903806113aa5e39ca74b352f67cb15f171ebaadec51943044cdff73969b02f7975d3fad7d4bdf39a0bfe40af70c7670af42bf499aaf64f3c31bdf183d8ac121f5aeaf3bf4fbdc4132ee0df954f9b6737e97537646c4f4884503eb8848b1fb367c05898f262eac4d7a65dd891539fd5400fd1856ae169b4a4f2ef83b998cc31b6f0e7bf6418b4f35b8b787d633e424cc9a3c6d52a2dad826d5cc1603abc6f6544ee4eff9e7e8a444e508829933440051945f6e4c5d282;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd3a67f3cafb1848e6c799fb4658a6fa3f11def19ff102925148d8b38241ea4b3482d5fe448ca0136438efbe7082d67e4b760eb5d0407b94b0628471985235f1b94391c57b2264abebd7ef951c00bb9c05e13a5c7a93a1d43b9c029cb44815800337cecd623ea0a207c4ad25f91724c0e775d8ed5c59b60fea198465cb2269dfea3106f2758355ee29c95061b830ce50dcb388e6dcf638eed6248a4204c71c898e77af1f878f45680f62d12099e020967cb95668ecea9ca8f82360127b556567c498a5d3487e733bed052a216ac13f494a269cf197190f0f5117102a329fd08b87f03044db6997054ff9f8c398c4254629030b8b4b0ce631e1d7fcfa82efe78b494d4d48500d037fdd9db76343062e8fbd87eb05f50ed10d9a1786efaceeff1c009c55468acddca3b9f5b06545052e2a97624a3f55257f40d1723b14487d690b624ddbece386765a1e66843ddea09163e94a041a85f088c28031555a18ae7910afe98d4b63ef41db3155121b9c0497c8e6b3acf8712e3a11b7f2dab729f647be19996950bfe3c4169f1a101d15159c91fe233b906c755516c2d1d0811886feca29ea5fb468b2be267f7cb4092977ebc8c11928a9a184631ce414d27a7d7bca9b57f2e5ffb9619b4ecfc7629cccacb51ddaa161893f2ecfd7846dbae826c49a30475fd162b6df66f1921dd119c8f380995cda480f984b67de99826ce78bb4c378a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4df408c34839dd65efc8857c7d230ba4e152e1693a6ad15bb2fda17f252fff1d67532866945dd11ca158a813e2e68e4f6f9fb917e8a653face50219e97d4755a57db13f81a1ca23902529937bb7ef67f305b29db0ce9952b398dbf28da709b46aa1cbc86cf57d475b6027c876ace400e8186689dd4406bb863d4365ab009f22e77e7574d4f25502786704c92fa1634c9a1c6545d47cce08471cbfdc02852f055e77d904eaaa2d2929cb2a990c2918c3219352c97e4c1be2c1adeb356b83e98bb9c28494ffec2556f2ad8541736bf9c47f1caabb5fa17003d518c20ad2abc69a8d924544f00f92b45d7f74fa5bc8b5270abac01c8180a9dff5a600f69aad8b38e1b489f07fe1e6d0cdea55bb2471519045d3f356ac67ef687c9645a70d090481b234891469cc9ab9c5f6699f768ad35c3da5e28a1772a4080c79cde874dd793c30d05f6030c919de65d63f20651b23945b38b9bc36fb7f16e187e912ee63e0891c46f4a2551f71eab0acf19bd08343e0a140ff3fef813c154f4dddadfa5569b07864e83272a99d5e13f7603653b58a20eed9451882059d148dc149126f608392f089995a0a575019a5204cd6e988c0bf33bc4d8e70d2b1e5606d71a9e575a23ac138e729ec64b9cb4ce791b2f1b974d381191bac4b3f1f7abb109da15f58fe311f116fb060bd4c301b10096118330c793aa6fe7ef6ca9a7315f0ccd3fca9cbc74;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he227aae88ad80572a1079a1f0711f247b42612608793fc37320feee63efe9a1e1f4d7eadd416dec430fbec64975f802b1ce525588b228131f73a3dd84ce964d4cacdcd286ac51d135310242264e852011dfedc2e1cc7870f20d551d6fe4bcfeb11856228fbdf53c3000d4d7f458f417a3ce99ccdba62e74707368738613d781c66b7319e014b11cbdce5329a9527df7c59a72118e6b6c585bddacc2e499817622126f0f4705103ca810f0593f7d968d6cb98d0ba95f4cd78f1508f2aaf30b74dd2d965966826d1840ae04c802bbd1785bb4de20073bcff94ff6f4806f4523bf770161d30fcc0eb3ae81d39d43b185dc00094eaa8b5d0cdf94b835a0cc2cdcfa806e1bce01c5624c5effcf386f43eb04a7848196597f61640fb3249fbb2e04c422fcd60808dffe9b30f7aed887fe6f4d37aa808cbbb7393d763b5ff6b6b00f5d40974483c919e1be9e9d9743b075debc37080af25ea47e1bf3e0957b27fcca38ffd41987ed905665131b19fcda30ff10f3a2b5a92d742d8905e2182c603539db3b8b0a7febdca285d4ba6bca8565395c52691e25ebcbffc48aa998bc161b90cb0d87f85b9a04559060679b1a783c58a6f26e0ccbc0593db965f54fed43deb91256afdc0a829202abb92b580a0598ecf2bb9b23d998747b2edc09138e3ca41a599baaed07fcf5bba38538dc17004d1cda757956888526947af2202a31c92864d4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb7dee15e305b3785781ceb3a7491fe5fee67480a8264e77086b10d190c5fea185e92827a1617584be8e8b21cf1edfd2bc3faff0fc21768f2161ac26b349644beded7409e66067b730598e85ea1ceeb3147069fe6861738a2aa396bc97281743760e7fdaa723ccceeba70f691b1509acbe4437a260ee26322cd1fd3a3f85096ee71bce612439aca5d59df13aef3ecd57e6926eb9170a6664663277775eb3e5114267f7073ea54caa5147b085f3847c46becb3900736f5995653c8da0477e2190e2eed3fa1903874478068a68b53f65c7462af35914ea3749d143874b95d3665f014a2f6f97a397eb872ae11c9e05d7caf8034a685bb70a7ef9ae3d713e34c7fc8575f05065f12e47024567d3089ca6792e5b03064d92119a70a6f06853d5207eabb3eb0d7acb76cb90c9c3b99058729b61c4da33870a45a7f9639fc6cc4ec32863542b261dee3481b4cf18cf72cb21c3816e0b71d503cb151c8fe0efa191026db557209036eeace18423865675718eb72cfb1293912071b83c280cf44f2c2bc381ceaeb0e52a2fa23cc56519af2c7841ac3f3ae24b379afd90ec2eb0e007009d82870ac4f45c2a920c9f4f427e4eca0a8fbf95c97425b1b0058c290f578b069984c96f7307dffec5ad2c2b24b45627fa38865d289293c0af952bbe67715451eb8c201e441323f3dfc7a6b1673b21cde4fb37de51151acea841440ac89970cace9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4467b81f715c9da583fcd69b1738ca9cbb611869155f54a1b7cc4f3bb02568795c31407df878ae2085b9c4e3a939d6148360bcc3f253dcb79f29f0e1059d06e8384600048a787ee8bbdb3aa099bc031d27b0184fc01f51fdb9134f93ea4194963b43adb7afabbf1d5be40ba0f50bfc0dddb3fd5c1666621845eb2fd3646951be044d57b597a9f14f99d5edc7dc1cbd0e896423469303327bf845fc7e3289df4ab0fdc3ef8551501796449682c8a5ff004d03cd9502c3f782e248f17552ee70f07d9284ccf7c82d0a698c482619630f14a64eb73ad47d5fa3eb80978aa6e142cf50bc0e1c4a129e97d8f751327e6a891678434b962a2a1456be85df7a938fa904df8d4c2464f2e754cecb686aa27d4c29b6ce066286c761fa508f1745c8b0ea3e7607254f5e5f57fa9d62bd12292d5b4b53dc025c21d03e001afbaabc1e646a8d42437231d9ec4723d23154b771501570b5a29eab5a2d61ca96f93af74be13a4888dc64f0a92a68f0e68907bf7980062860ff31af7d8444524ae11120b649aa54240664462e902c29cdd6bcab4190bc7f7a9dd7e3980cbcef471adb1df2d7a827be2497234d3183ce72049132fb3e0866c6f0ab6fba67941064e8063191e70bba2132fbc5e390496ac9c73e5b87a8ec0e202958d043d9d026b77eedf915663c14f9979160d69c1123ec691ba9c070dd2b88a761f1b40cb35b8dd1c1192e6907eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h713e91bd14d9b3b7142a0da168cb925ed602a8410003eaf6a6ac6639c586f2bdf92c9d50fe54cf8d89777632be95292e770dbe21bd3ac38719c4afd520054a5fe1cfde23e6f492c942c5e907319ced466ce5d4070e52c710fa457d3b1018f9d4a123e05ee61e4994a138cf94425a4c12975b256e58d44fdb3395f4eec4119bbb8841dd17d448e82fb1bb0512a86edb1b47692575229cc9d4a94dd6a19a16c0bdff101fb80004f97ed41f18a7a680d13cabd6864dc4da250ba480caf2ce7c68e8411960c0c249dedd46b9675f5cf11f7dde30250f331845d775f860d3172181c8a314bc83036dc7b27735cae84ffce3f4245ccb08220bf38af50544f21416542820c38e57257c8103c0af4adea3c8454d94db0e2e8c121c8026e78015ffd128e67abac4b78f88f02b6c16da7012ff375929af983ce88f554d811e1c115a0350b9231133281631bd1d03977ecdf4c69b1fa6a0b25dfb6401d367f65566910507f8dd4a732b3c72b26dcd09bdbf6013e8edbdb934264695555c2511902e27457c378003c87fd60e26d86ed4d9526770df457aca6c9dbdc7dfa2e0d861c4cf4ac166d4bca4ab43df308256518305453ffb6c4b11fbd23653566fe9ee20bece32da078bdf0257c2b41e3cc530cf896441668f754ca9974652d4a1cb2b1b42ea78ce396cd052dee1f829a3bcb3e69963d34f7f17bd4eb265d6411c06686c0882e146b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3d4937a0321f7fe8764ff85f767d553e217b770560f06430001a8f019309e8585f6137a4b725ff078883735bade9f3c71c5b5740321ea33797ee2119d3e5254c17d8c94dc4890daf0e6ea6ab887184a19ddbb16c53f28ac1a2e7e505ea525c854fbb7a591e015aebcaafb89501cfecc928cf1958b24232ffe89c89292d225170b249d0f93cf277f548e1da047ff31d4c4e50353ff14dff022dc656f3a875a48aa5b655e49dff78c2fb2ac80cf212eac1df5ec157a1c8ef61187b1cc8a9b19f3f165095805fad54ff678cf00bd74463cc04fa3bf5f764081113eaf5166510ff4c4c38a194450858af87b973a8aa34ddb976ca7493ba0e9231ae5ec6314c7d905327cf0badede2c57e0a9f7e44dfc36805488687ad4a5ab100b568c8a0b0c49204a183455e3dd22df65e0f6e0ef2907fea54f187c1ecd2708ae0a1d69d3fae86759408b1b0425ce4b411ecfe38c4d3973292c609e0845f803d45baa9c0460598bba1f97637284341195c32ac402e961b80a76512c86ab5b29900a4f8874de2c589e3c89a96170abe646bd8767e6505d98b839951ea78c16c72011dc4543e7e7fb2cfd9e29544161e81027510af79768571672ebd47a2d184ab1e98a4566cea40ea174064075d3c1ec77a4b00ea82bf9c71c63266c631e9ac34ad7a3b6ad52c372a036905e68eec19250227c52dc0c72c5d0e3acecaf0ca11121ed18b70dfd3cbe4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf8d97aae3b7d5bbf36e3f7e77bcbc121fd65514548db5dc0ec0305d7b776d95a6db3d25e0b6712e591079b59af39a82c4185dd97a57c72914e450908c054b7a7d4a134a6fabef536066627aa9dba86e657450b2802f2bba97503369f2911d56e6e2f76567575141796f55ecb208da90a88fabdc67de2943c8d7a20ff34c89c85ba65ce017965781006343514c7e3fdce78968ab28a4d193b5cc5e9ca5c3c3fc95297827913f2981efae44c1b4ffb00eafd5459b078a410a26a1c3ff08584245a8fc6cd58c0774f2680602af9f64d2bb7915266aca237e8e77b8e33f8fb2781e99acc672fcdbf5498178daf873c7ad545cc3d3ad0392bc25857a742ef4524ec5d6e4f9d8a17a6949b5911bbe1fda03e9d7bde0d869828febaba0fec9eb86e413cbe97d72076df8a580b62dd1c73dcaabfa50f99c617c3dd26735af2267fce14132b891e6dcc12822901071293d3d266f2590706d9d3f7518eab80361b83a9c35e9f771b432c2a225358d7308d8f70343fb471e9311f65f03f278ec3e38d1318be18db3083a011b4943e7679ca7385b213728561d5b7729233917f7e9c890a423d1f14471a401ae65560509ea95601d8784cdf7a04d00707285e8f8041031863c5c040cb44e47d23680892accff9b0ad01402af05ca779520356e3557d5ab5e0c0feefd948c6013889983226fed2c53640d9281b4ebf848315283a207415ba0a70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc2bb6a8ecaae1b73952b38c14c0eb500599df72712fb866134f9bfc6deee9ce47b14f8618242b0dce240c5c0e92941cbcae139ae06f2fce5e150cac5d94063d66415f779109ead817d1fc4b8e3325df7e3c3aa1877342ae204d675e986784efd66b2af734aa8d4e40976851d5602c378895883d774ec7cde3865bd9e66afe7f9b6e6b9178c2d0aa1397a434133060867ac7ef4d8b2ae5faf3edd4299702c92c9ebd4db5dd176fc6e6572c24b6e87ef6bb779e18d386dcc7c0dc5628ab0edd32c1cd971ec7fbdc4d2ca7493a6fc5e120eb35a5f3fdf65a75f245b2b48065cfc25bdc022361033eda1095be4937ad889dd8f0f6ea8f6a1ad42b03482481b2a1525a457436b249da8519ca9a47d54fdc73adb5a4ab0a52f7abf39a8edf42db913f9c8939708cc6b6dad6f1434703182e26fcc05a31fd558db4574b08eafa5c94813772feff5dd3838c158f6231993e8e1d0d228857f168f821c5d6bf44f5afcd50e374008cc89ff043740178cadb5c50f84d4631cfe684c2138ef68821f6fb884a73db0b7f3df4371497a9e4d0e1b44c8e727c01d6030cd58e192c19522ac8fb3d70fb55017e9b3af046a2ea70872f9fe6d792ade5739a603288736ff4a802ee4804128fc3e94aa1c3c559b9a9ff120fad8063cae5da83a335de88a888a1ce01e1479b4b9b1f32770543b6f0d847237e8657af67b7a6117931be099941dede1ff3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hdab9f302762dcf6707fc3a3040c33dcc6a688922a98a6b8f2d5726ae9b3090a6502a043d5fe6d2f1e690b54bcb3d9e481162a589e024e696b68c4ee27547d85b38b911e73d2bddc8858c950ee26f8f2538df6b15f7c864daa8b3560d2aba9dd02d963582c61b04361712b10acb476cebe3f6ecf6639fc0fe7e1b56ba189e5bf7d6a9bc76b81a8b0778f6fd702085c86ca29417282481ff3be5d3915dea709433a7b1fce97557aa8fe5acbb5d3d5192eb112e1b521f46c87cd24f41f86b78dbbfc2bf04f863d5b29f944baa468cab00f637e2d69092cef62fb90cc86054469ce984a7d1c0b5d05c9f0e7a5a97f8f2e92fa8d8297688ae549fae60b0c083ef39a0f789fb8701f14eb482cd80345a5bbd32689ef480e6fe8eb0aed4660eb7dc1e1349748b0f9f8e6478b4c5dfba24eec018d6dc59a3f3a9977cfd087e02e80bfccec6a26443a0d891307c8ed1d6edb3332a18034e2314bd129fd1030463c9f0de89634d3907f5bbfa639c8b1f1004318917fb6959362e40de7e3c35df4fc0400e924ef65c62a8bce9963428f5ec6993c6baab0d5cdc959731ff460aa1fe1cc2dfeabacaf77bd204584cccd4a21b64b08cd9eb337ceaf0a42d731141c96da7322ee92738acc91835002f2a29a8a220dc337dcb0abd4c5a5becd674c16285462e1fde3c0d356f675f7d763d5d100ecf2b96538f8ab94c6103d18d866505155f753b57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h838ae53624621fff0f8ff5c23545ae5cd1f33649f52fa68104d0a80db138d69af2d2dd2877d3f28622f6c2281347afcb6651d4393c6e696da12d9d3de6aac5c8bf497ac46b762951b4d2b79ab22cb4d3a03d3f42be3c99489940698c32067d1e34f39183242f0082476695531b60f013659b1ba956b7fbeaeeba2957e36f80d7edb0e0c5bfb97328aaa7ac2be600dc4cf320a214e707b63d3054943d834934f75a20f05d3d8e3be1a904a73d7d7794fb3e0446c3e5b8350f2f2936c0550385d2cd2ee007f66fcbb0608cef05c151f6c45b546da05ad58dad7db6ae275ea024e1d4ed5c417fd2cad807bfd65cd91709b5add86a60f1f39dcf05942dcd242ea6dfbf017ef0cea81c50e11f074dce4fc526767fb70db9debd857690690b8476af8d4fd347834df00883347f53f6e6f5e39c69f2f3ac2f641ec26cd14441f5e532ebdc76620dc680452983b553a52ee4e65e6885b53390cdeff9f5d09349e2de52e05c21426a40c358e61be07d015108e0df669a2ed593c9c105d33b9ba68c547073ca62ec4059d3fa66caaddafc51ac06bbcd82e90c1d9a941026143b9cb2cf60303ec502f2d6ee448a027a99dfbc9007798153e7626bb05a80983dc6347d46fcffabfe67e879c28d398c05a7d2cec8b4fe3c719eb0072c2d8b2ef566fd132208ca1dc60618f0545c73a389b74bcde96d0cc9f9da4c5b48ac187f773a58a1635913;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h28588d132f93fa0cbd4ac005649e5a610d53849bcbc4a173a22d162a0bfb6973e18ff1cc79220c2b36a4da1baaa417220e5d64524bf607fd81d1aac735d0b5cdf3fa846930fa28d8056e9e0d0234492d5db098dfe7e112cb73998fc2f4e93de1a679ad7840a5acac2e1705fa56eb39a7171ef1faf33c85432bdab065ea23af0bbfd077d65edc8dae7dc8270484b9aa35132b160cc5a6b709d48efbf914841078ad34fbe62924255137c335d66000382eca9741b5ff40f8fa4a9dd822fcb1be1f425bc321763beabd605866fba76f2a34a6be03b1ddfea8f1b130899fcc412ccb7b1109412568664bf2e685f975183f14eb83371a56d722af6c268822970c5dd25bab5bfd8540be11750c07f4e08774318fcb163c685539291b306dfdeb42da11329c2515bbb4f4caac72bdc675e7ac8e35a97346048f7ef06840cf4c0c0c3e744715fe954ec86830a0bfead9a8a0669d06df70acdd8468e8bd3bfb4bb4d2507792c6bb46c54abb5b996c6c53e4ca387cc6ce81074bffb54d0f698445143813400e0de7d27246bdf681490fe51ec6a181a96a2799db52eac200d30523befc9f572e1878d921d0ab57e05d9b33a5c50ed89e5df578bd9f39810d3662592afd3f43e657f24016faf08e77f53b4cd67618fc2f2f704801af4f2bdc891e26d93789671e3541b072748c9d24cacb5c19e8373e478c49b53ee4786789ab44a3061445fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h891c1a4a398602c2f97c6fb1094280d1cf44895df98e6881e542c19ebde4554e8179ce5ff2933d4ab2ca137db8c0ca4c66b64ad34d6777dab6d7893909ddd9e2ede48b444368596ccda22804ceaccfad44de5bbfcc1c88ea986f073eb821034fa262155390ba7a5ae8e05d2d705545d40d60168f97e1c0d3177c1066132df4ab0a3882adfdcc33178ff411e20642bc62b9c8af8f68f52e602d348f7ae1ce8740b9cfd29ad78278d8f5b0427c4223dffca6c0e34161025d68fc8966648428b49abf835e149bd07c1cde93c3558620b301296cf2f65e8480969c9bc3213126693c9965c67edc481aeaf19dda2d2b8343ecce0014dc66a167392ca496af8de25d3ecce5238ae6db26f9ff7b607b590f12a5cd02c619efdbe27734508dcd595e1fbd874bbf9a4c375e5283d6a4e3a8491a6c80f845dd736e1434dca02c31ceea7a75d3690ffefb32f5340da20c364ba57aca0ab01d3fa2b140be29f0c6ff1717b35e6a956edde501753a53e20119b59c9d41187cf87b43a85ea75231a00d8bf38bbdd188b135af93cd9f4848554bdda76eae916eb6f1a6c7c841ee59960adf77645abcaf8280b3d1462e91f866fe2ff2d0234ca3f582692afe1f60ef6decf50e7bbc8024b2777ac8c0e45424cf1384cf825978c7de299ff050fd812202248381cf8b60ef2fde96561e83ba8e09e94b78a32554d8fbf6b9c7cd41a64cc50b8c8ffad1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd41f5330c76c134ebba785750a22eaecee338e4750d0d1b13ff69bb22a9fb6d4f722b8a790d35e3df3a809291a420465162ba395457d2f54c1c05ef4a791a56f7f877740eb4561222bae725f37757c17725bf69f5caad59416256cf35dd6295cd81b5d6b31318300c0f0fb20c4bbaba8950903e78077ba5abde4dac9598c66ab7c0f6415bc08c29f743c8fa8c68909abd915316e02e14955111265248545f476c34a948e6f467a3c25841bb2d7a336b9422593d9bd61b3d40d6f681892dcbfb1963dbfc7a71b150df12f3f2e7fd9580990ec33df1570cc90a3a299dd2a5369fb587faa7c5ceb1d6a0615a65722a5f610a5f0b9ed94a1c12cf54df65be5a7ce26af67fd5b4527aa20abb0ca3b6f1327944a495687491ac46ccc995cdd0bb41ff39aa69b1bfebc362e534b0148157d3a01c03979bc73bf3bdf3e726e9bd754531eef13557a78cd6f9777949ae3d1d3dd7972e89a98718e9494953335ac1d5c52ff95d84ead88cff2e83713844ca40d1ebe70c3413714f9f6e78fd843ce3090243e7bedad763906cdee07fe7ee5cb48b75728c959ae1e2b6b9465e38b8cdf930355b5f3582829f7dc4dae2416af345441a85a490cd919a7b80f589fceba34f6b5e233d432a7a0d10a0f203d8e4cecbe59439ce68011acfe15b2ac562479e4848b4a5c1dd8fd216a99bdd19e7eaf6266d3a9a95fc8db635112ef31cf269958a30016;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h47db79fe1efe8c31e233a00deb9fdffd2ca8510381b8a6fc5163589636fb5d2ce54f1aee134d7ba7c353714692c2f1cc82ea1a03f9862f23b74d96eed54af02eaef4dcb5185ba211df9c10a274f3e8d067f388e2a5924eacde50c2b4e0bc64e0713f2d1723d32947b220914dc95900a5f4dbdece04796a7e43ad3fe592b062cf86b1819931f5a3a7c2d1ea19dec630ba071768a35bb5940bb0fc8e1204ac66e9f636032f90c1e41888a85d06304d66909ba3066c375e8376565b17b944a30014e340da9ae739ef140b50d6e45b38b4d062e54d054bd171a9fafb3c542b7a86919226a4ca416aefd5e167df0834f03c54e35242f618b484464652503f85e2ea0e658eab7809165c7af306bb6b2e274d6c8780711c6ac2d5fd16c96f6eeb56bb89426c0afb348007682f1b2874efc0c4efc31f21ba33ce01ec8fc023dfa9f601be787cd54741680abae4869da0a1b4d6e5558f37bfe13215ee71da2763ec7fe4a6e494b315837fa54a395c1552d3cc5adfba52dbb25bc37b1708ecda0e3af8ca07fd69e597cd1f459e6d48fc8ef4eb98dfe9c15256b0513d6d10be6c907b355b83a13aece03233901863479e2371624f007793bbfac5e118dedfb4fb320228804ef65bf05adc7a9796aee09527dbf04626b79b0161805684b206c3ce2aea5276ebe5b1168f5c5a85930f1067e2dd0abeb71bead1a3a5c5a89b37b4b14e9b3e2076;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h9dc9446c4b8cf5769f982b51fad6cdb750f14aecfd1fea64ce61df5d1b86151d4206fb12868a701e64c2ae23c35653b059bb3df6ef10608bc5561772aec87572f2b22465a8f5c340482d4dfc8ab3117a23dde064d0ddeeba9db7cf28aa74f9e093769e1be53f7e4136470a6a992925c947643031a7fe541bdceb1c098e7359de1c38aa48b8a64d90feec1bb9a1ebb112909d5873d4b07eb59db3e882807527e180ec410fe0f089807bb1bd18b175942d00965b2c378e2a8796b37b44d5652ba4a64b345ce7370fa2596009717d0ec9c0e0a1a5ffb58fd8488442bbd7e6e6b10e12b7fa40791c89b9da240facfb4861b7c78511b49539bfdb11ef63e9248d1d1a5f3dcfe74f9e460d9fe8554edece36fbfa02843f7eb0061f4bb404e197c050e5b2cca5bfc0364f3e9a2d0c8e38da7772aff0880e72149d29174d3405afd42d8bff21a2739399df8c11fc6981100fd9857193c3659026f6be2ab39e50e8275b401a90b7ea3cd14d6a26c02f9e2cbdd281cc1179ce13045ebb7e28e85a9a1b475dcb840e9b807ae81ba34b83f6176bf49cdc9d6c7df2b72fa69015596b83f5bfc646f15a7c512e45fe0e8a6016a71573dac50de329b40aa35d4546d8d87982a15e89294e9023ff39d6173c3ddf3768fe7506750c06ef5799a126a78087a0e7de31b71e8332c64e2d9b24acbdc21cb8b6a5902f79394dbc80b347acb59bba3d239a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hedc52fb8fe9400610f665f6a150c9df28ca94dd0990d2f1dfa3d1a9574189fb717da4bad33e9dfb140fadc1cf2b4a7484102a9dc9527eb3e1627b44ce9ba7c4c7cae04f0c201357e112dbc3f95ba0a4684d93b1ac6924c37f3faf8d436c299027fc534b3809abdcef1544bda7b1830ff7909981a298c8406b938a4afb7db0e103a62da51399b012e03b138d13e16e333f169307d1e3ed4d7c22e36ff58f5ac587b8529e74e2ccade10230d3a61a241158c5e25dd812491fc17be68eaf7850d9e54166f4f15074339b98c26446a185f1b1db1cef3e567e2acd2e4cc6d2731155ad26e1898296e858f8174a2ac3c174145e42a86539515c9605ae063b62c16305ebfe503427739634122df0300671f1ad30c9a13c1a3a641e7dc4e8c86dedb0a50c19d762b1ad7b3b037918bfba52c81cbe14cffa5d1f8e8dba840f834b4a20016a9cf884694e183df793d3b6f6cef93afca9fd2dc41fdf20736607a3fabf4560797e3011e2849dfefd68163bf4b844571cd53e3b3b290d2f264c67c5a8eff2fba392d9a2664c42c0520bd8762c49352da6e77852f61eaf12c63dc6eeee998ba0b02df208e9ded34182ce57b7d76b2cd975994ac13d9386b2a712e86474b7d6ed885e6edbf51525f0c057b73fb2430719ec8d0cf79af2280fb50a36437dd205fdde53b3588f0da9ccb968d81b3c8828628f8b8ee30a9c282feea0656f3d5c79ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha56e8dc1290804efe06b807fef8dbce6d2733c4227db553497a651de79837dc0c2add9caece234ccb597fdeacf2ce48e26184a5e5e1abe4c5ade9c51f67a7f08a089c1d6c8ded5d5e845c0b596124182da72a7d8ed51db38d16831fa1a8285dd134df717fc128d78100c5b7cdec5bfb9a862409efcde62a0837ea4cbe3658b2f98ac819e88b5a111ec8bcbb5ffc9f93c95969067a42425bfd09c46c1a3a163cee57627c2dff71cc9f3a01d100dee9e4f30dda70962d0b14654884dec4050c8f958acdc9f7f45aca634ba1e200f6b67c898632a8fd2b84a54b29e3dff26c72521097a439674ae0116ac76b9843f84863e66df8107743a1b885894afcaf6692d8bd34923f9e66fa799781e10c7a433fade6b176b2779f62784bfc8fcb845ff68abc9e950bec1fb6c62614dd21a1e20370aec97fdcb34aa7954510ccaec39276feaa647e61e4a7f63e03edaae7e0d669f7c9418e9e5a2286f3c90d7a9783e6ac785f3520a35e4bdf73271b398bffd17431f988521c4303fcbb89df549f80323aa6eb0959bdd373d367275fccdf9a66e32930e8348e78ddd91ef7ced8549dd08031fde6e32cbd8a9710f7ebf8800b57fb371a0fa1c77f92dbcf5c7b99f6cb4319dec3f6cb43e1766d59d3d812db3e2bb159abed15580c39190cb5c1890ef5d4d9631e1259bf8dd0340da0f03c72a7be9d3088616ceb6e78fa492872c6795ef1421c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h33395487da98dc1b9c711eb41eec91a7545c483359f2a0ccf109c9c6e7aeb38fe4c54bc0d12b6869f8631322f702e72027ed893443ae3f788dc996939338b6be4e9d297120ed125f9c8db4b0a76bc7cde1115c67136a4d5c9badc896ce2ad5cc3f06a6f0ca7bc1c11f9ed2e9d7a00e57cd75c44f04a41f0bbc81bb8cacbca7204fddc5454cb9905f63bfea07b6ebbff70163361f807b1077ca6d7a1cb37a157e5146f05160a976e8d074464e12ddce07c9ae633f39e8a75d63ec9095295312aeae1bf7145d0dd50f8f7267f05f02ea50a39375747d456736cb42e890e6e82bc46a9e60b34ff6de99fbd5b6d249cec032a305dce79ec215eb8b386fcb3f47d2a59523731a3076bf76719b8d6d6c508274d6e74868bd097aa733e86395d2f71e9ffccb203ae03e541b41a461ec3445e5dad08f5d47723a3256b09df226caa79dc277d17af884d7d7676601ec837a01ee3111cf976376cb362c8ed1e9a6054e1643e2640806e011d723bbdcc81d10a806fb6f3f6d49661a0aa473b5e50e61c9965c48f9cae1567de93b82dbf26058543babaa8cbc72a2958037e9531d0641ff8484c4c239ab9a86fde6db11095f6fa229ebf42edeca90b7bd7812818801f5746a5c2bbf8d6b6adb7431d45744aa6e1b29cf8e7272f8c44c0e560f7a640fe7b9a70b3c3571021ac37b6bf9d05a8e74dc32010cc099feb4a46716bbf6ea0e90a45131;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc8f030efbf4beedbd8a0c6a5eb27b16221fedd005e3d33e6dd59cc01aaf4dcb86b23713ba25ed513de642bb6e79c88586c499a43affde88c7fd57656390cbbcf6b0fc8c1629ad494f1e2465a8f9a2821c5cc43c649d309c623e5b0af356ad185b81a7397ca2506b9bcd7e211b9072715043ae2944360301766e9df25a888c8fa6642924c9bcbde70aba4f1b4b8790ead4c14407374e3b30959694d68fcaef29a64dde25b0fb8be8d9862a744c872fe0fc689f38882525afa8d7724e54b733e299628cacd1a38576ad25cafee228240c99e584f18fb479f627ea2327f0f355f0d26e17b58dfa52e7f010539e246d9ee6294a3e1602eb4efcfdcaa1679539f3886570481e220509c24807e889dae8ccfdfe8b0570737213597f46cddc85ace9304c1350892c17cb3d5629c56250ebf0f59079747f4934322f624e0087652616868ea030863a179acfc7e5fc715f969d7752eae026b9c5f69046bc69f858c62aa7e4a17ee356b318d2d24082297003056d9d3b5094f5bbc87a497bbc4df323c1773ad16a334bd85b4c57b1775835cac5ccdf474582f905ec6b3ec2850d5c403b253c7a768c139c3509eb2e603145bd88955eadea87920ffd9f9bce806f64295f9652ae1d5c866ea155d6382b4dadd4aaa197d4b92d5ea7dca13be364e4d29a0a88dd7e22e30d7c0b9da6a1c9ecac5906d4841ec89db07cf87e1ec52daaf285f168;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h52209a46daba6574c12ab2515e25d0e1139db467c922c96dcfe708ad9c246207524f2aeba5991bd76cbf5ffaaf5125fd5d375a242381e6fb18887fc9f8739b4d204d062d3fabf1d31f8593314c30798a98c8bd9f25cdb28358e89fe2d4b090b93a34cf548b959460c823bc00961186bdf4d759a5f366786b276d39f22bab4b7a40a021e52d546a47359049c4537f011c49f493c009bba1c96b51f15e4cdf749747169b6100a454d051f5a73ecc4347aecd1ef18bf9f0193029b088f7f1ddd29ef0a147d495e31be356218a5c54e7209d7e03babccbf92265b3316778a80485a505b4dc6c677c5d07bf38d45917a382904f4317420117970715f8344dc611bd7f7673aca6c9029951ba1630085a04d4058dd1af515f4986d12a5edc7ac6fb92e1361d70bcc13da415992a0b6bed41401887b91754592bbc585a6ce8249c18ece1a017aa9007a9e6e27093fea0f64c2cf74d0c67e9aa20c774107ff360c4d3b61c0601868bc136917fcae33f9ea9f914bb3d0d3e2ed5ed2056d235da101eca118087be5f07f51f434997ac9bbae80430c2bcb8fa3611b55b29abaf532cd728d5007f2c44e168e82ce10d4b411df460efeb83689afe71744c1ec7cbd171bd6d7244f6a9a61cf0de46b57ebfb345bfab9e0ce6f4036ef9e1c7948a61ba9865b3699ce739cd7f82350e722159f6e257dc82b10843d6c77b79a990a9489612a079f31b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8e15e808e818dbfd6cba61ee6fae4f3362a59e18050f9f6c86e8265b09ca3bc394c9f8fe2826327b81d8e0cd32a293442fe6973501a9a397f6d41d7f2da56e55728e2261bf1c7ff15d48ae7d5b6df814735cd0f2ddac01e2085a10e678169f11f137ae8a66de037a79a128d08300b5cd42f2e87b51e460052b53e773dde480ec5fe42ef5c5058483ef039e38dafa65b5b856caddff63db6558771e17153c6ba51cc430be79ffe3858d9c6e4355cc527730ca90ed14667c67e7fd9f21a15b1164f6811994809eb237edc8692fbc3cd76c53446eb29522d362f59ca94ae4a47269b3cffa702a2e269fa9dbb39d616b637e9f752d0e8ae5474ea9abc62223f1a53bb40412ca0feccd6718e961e7e4b9eb446f654ee4b9532d05179acb7e3f4d0adcb5859149c706a3cf8e4440f82cbdc54878a5c2b13bb2994b44948a54d5ceb2c4a4a543990d655c0a046a3addebae798d479e807a9cc7f68bed2d66282d8bb4308fdc98acac78f65fbfb4470552aedbad9931885f4c0f13e9554b4dec2c6a64e536f593c6d83bd3dfd737fc05432c276959a6ee6b42546a67e917fc8e5eb5872a1d8e981c028a3ba4216aecca7c5ab8ee91509d37289782272eedb5df4548e314116a377183cd45026b264fb38de6732b45c43c84d5bb6f030486dce2772934051469864ab86e6d16f4abb8f31640d8636d1b5e41b446fce551e1095d38f09e06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hce6ae26e91d02d2f7ce1b60619066415d3e9b6bb84a54b0ef6e5d7566ab87948d7c113d201806921b5c190b4cc0068067cca847c50d60c48f2a47d6e7a262a6cd2a7c0488ecf08c4c4b5b426e82c2ba8a1d5e370176f3ab81aa7814ddf622d8889804ab75833a3b71e847970d0a0612b9b186b99f9955e2e514246b2333646d96824b9595e2e98de62832b1f51dbe04fb5bf48654e34b1d3c5aa1e0ee22fd801926cc91c7f85069a9f4aeb3e1c9d70c02b759631e626598f45e8234c954751b2d857472908c6337e3dabac0ad75a94572b0be8345129e3ed67077d777d9ccf08416593d1953e8ce759a533e48d5096fe678dd5a3d2f9e629775c47b17dd2e0e922783bd478950842fe9e068e96a4ac53697af3a28bfbf98f70f830c9d8260574adfe9e29ef21df5bb3377422b93cb170caa9d2f7ff2c2d477a5c6c6e465a8e6c83838f7bd8c5c9f79a28236a7bc84cce9af03a0de3b6ef523c496362b07a776282af6272f09f71dd9994da13e42607ad0728b020d5e6e116430cbcc4952522200e6f2f6cb4bd771c793d3c696bc94dc61050e81f31b1aac5b35c13eb79e48b43d53eec3f0af7e1542ef1ba679ac296726dede58485e9552bfee6f081b4b83f985fd824afddf3ab15336ff0bb39f6707911ffb1e41463c0e17111a81a5da5889037afc0f3e168a4bea92dff5365d3ef3790f43e0866238f3544accace6745f138;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8c08887b978c286d4e9e72116a36c96643490760ff8e2229b73980251372685c2b42457e8ccc7a571c0550f09f2df5feab6e7707bc7b1db55de2d4e601b2633f04acdabf7e995ed716c8de256d961552f2c6e3208ea24836a7d00566dea95b80bb5ad5a06f41a48e720bd4257a44de2ed5baa9ab35c3dcc13e3a85eaa70f75fb87ee29d9c497cba70006c080c055d18865341a4fc112724b6825d79e1e17cb66e440ea218b9223ced918b6fea03655b3e27b5dd2d9ff9d7d7d99fa4d6069d4a08c577e9cf905607a54084967a6fd4da284d03253ff682907dbee6c43c9b87f3820582c2f59be34fc8d563056eb61df0006b629cbcc3f784be0741e1102795b3013fb68c336e7a203099db221b88472f98b6cc107f7a11cc7877a59f768947c267c32a0158e10d2e0bf9e4e2d839a8f0e0198afa641b07f3ffd09db2b353629caddd5333dec78cf40b10442a7453d8321d8c13cf17b043fee32a79809419111cf0dce5660b32161d20e646e12e81282c1a64f59b148f8171d9966084d3abaac8dd9f3056310ce5e807905bd74eaf153a8114a12de6944ebf8782497c8da54693a8044060fdfe9235171974cf10b5139ce78895e73fdf0112d40da7d02cc0e764fbb84c197880b39c7b97745036bd9eadd5a04ea1065f705b71f08abf489e144dd62dd50b04f47af2986fbd848899d7025ad73aa66a96578389e8e41b1141b5235;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h76bcd67bcd50b8ff91b2bc88b381f6d50c927b7746a423ea4890170704ecf3a0a3ff466993fd54a1b5b306c8c415d0fb2f99202798f814b73ab443e06aa1afe18d7e83e00f2b06f23e90352b1725f8f8fbb07eee8bdd5dc31912cc49855f060c7a267f04fcb093dba1dc434314109ca2a411487e3e47177530c3ae3e2a067e26643e4c32cf70d8fb9aa756ad050ef52bf4cf3e457410c9931d73682949125e81834ad49319b26a2ec9d27a537062c86bc24a2f82e41312b0a5f20f3d486fa88bcc530ce2c83c991eaf3c8dc5fee74c726387979870317084ec6b9f7fb62f14a4dfa5390ee9212bd60ef40730c156c95deafd2c76c266b152a5dfb41b11b214c56391b7a24bdb9998acf562029ce7396db677c713040f8a5a25c9672873535071e75017466903aa5d9077695c6fa9affa6d436f0e8357c330b4e560a9353185927c5b2410b44c944ef8e5a8cc1b9c411c18abebf5785bb981082f5a80a50737c89b10cc881e7647a63c76ad7ca53b9bf40d1cc578a81d427d8c8c65443ccbaa73dcd762a464a7e7721b4fddcd8007fddd76a3102abb9310dd33d17b9f354c41a8b1805babc701424a14233cb2bfa56f135adb704d2cfce6112ad4f12836b64405af17cb213876a1f77e60926e828ab15a9820ab78177724b8f1778d0a8e8d8a5a0ad821e9efc7b57129d696c6962b682da4b05aa2ebde521bef6bd12962686539;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc6d00eccfcec612804fbb8cd1c2cb3cb4b21590d6294c537d194b60c5a79d00eacdc3475a3aa79fdf477db9dad2e6b7b4cea7e3cd2e6078629741a55c96016bc062a4d9b5042225072d6ed16fc1e197a9a08ecfadc901d3ec0405f5db9f0df7f48e5c6bcb1461482456689210c719854b13eca00fc84179a610e936c0158aab58d5539e579f7cefacf9cc65c02f012596b9663ed7a0f920d408316acc0e03c9a938d2f2b212fc85240527563c4601b02e7b7a160b1be80799915415406a931133bb85be02a9bd98d50bb6dee2856cd1cc6b2cd9513eb86d4dd44f5f7f814087b1d4938632d2f6480702beadb3f41cfa787535630256e533fa5b1ca5bd5e62ff9cc4db7cde308d66c335ff68bdea18b7f8fa1d911909e5ce13eb776082d7018d77c25d5dcff66714a2f7b17f38ebac4a2526ec1efce6e508c8f01af59eb7bfcf0200b2e30472c50d1830ad8429bf14d25bedcb607a0832c2c8b02b3dad5bc20a70bfc74f0932965f51b0e2b39c46a50ce147abb0360304e8cc368a10201e20204723e4e1c332a20ba5419a9f1fb5c7c65ae75b83097a36af423d4a36f6c8ef81d4ccfc1418573353f4e0eba42a5fb59e2e45497f1a4f6df04ac152ed7d7ec4dae8fa4f54b460618855d72f1a07dee98f306cbb9be8642afe64099644a3400bbb1f2969441eee125b3522017596d54c0419e0067381da7fe7cb59a0e6e749e6e19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3a027611706291961261489e531a0e863c5a339f790ef52b2332dbe49f8f81e092b86c7496aec741dcbee185d5f4024c53324bfbfa90b93c7d2c278ca46418b0f9c995dce0648c4636ca1b1e1ab30afa6438b2132bc8bd21a5c7917fea03299e0362767b63b303a249875a30473214718d1dbf57962bfe7032377a68155646314730d25cd7d94b228f5af977b7d3f4c084eed1c4f69c971ef36f5da7a55941f35c03b676940e63ca80042fae95d7646b27bd563d72ced5dc015320b0e469fca2116aa17e9ef6283ff3616d8f4992c27b9a0cc85f78558d2dc012078486adff2991012433a06664398458c5be1cad60b8207b49a3bb7f2f5d92d004f8eb232fd4cb6889cbd968bdd62e76c130a8c57410e378005e42b3ad59c59a31ce8d162c9e95c4686a96463c30368a1d2376c60e5a814e2bcd3a412398f140fbdb0f01c86414265eac5862496d34e1055e57e61c461278166eea14982f7d69818329ba7742e411db26cffd83ca0299262a6ab0a88328e5f7ca7cb5118942c8e56b5b3fff6c679d93312fc8a9f28258e760536ab2fd79335a2b05e96f9b3fe7e3d01b34e4c2b393c9563eeae8a8ffa543d242ff5f2c733afd037ae9505067d203a2e9d5140226dca7ae181ccbf5eb8cbb907ed67e82399efb7884bece88656fc3749553642dd3c9ad2520f05b9754c5605dfe43f22bcedb1974bdf6c979b012f04d830e238a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h14d44dc743430369fd55c33bd58fd6776c9cf107add32c30894d4f790cbb8588e7d70f638b1551cf5a0e4c65fb4853627ea530e5bd8ee91b8e3a9a8c617c29938c9b6c455369d3536646578fe6e5660be386e846560c3e77135cf795e372ec7f3e92b3b5d187a8d886efcc04a24ca54af60342f1ab74d9a5655bc0ff5b6c057c2f930ceeafe6433cdb4bf9230fce4558d2a8fc23d516a0603b118756511ea9b2f1eec002f40797de1ba3217185711b5fafcb2c013482eb2e792bd0a1f8629da40ffdcff7b5719ec4ec3dbaf163ed3a55fc7bac523bb1a235d8cec2f565d5fd8c4ed5dc3c6778ac9a7081e0c695f60876d1919f1c30041758eec1f7e4269150ce81324cc7e79bef08d9c54c71bbe1057ea2c3c745f300a35dcd71062202925eec38bbf03872ae927b4b54f59f8dc53f4ada035906a5a5732945900aca7641886c79ab48060d998477cc1e66f2e94e3135cb622973ee0ca9d76f56d4bc10004321ae7be178b5935750ff80943720f1ec4543f4b05ad422b78b127710345f16267ffe91b4b56c33de4bc62c8e3ec676d095aa6b9481cc6491387ba7ae3691dacd809245fbc39132ad672a19927a7bfc4fd6c175473ba3740a260bfcde83094319e48ed21c5dcbc124290e6e3dc0eb04bff438fad558f9d2c9e611f40798a0e55baa3a0b81dab17dc771ea7999fd02b99d64baebd400b08c88858b7a02766451a24a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h77824fe2a9ed27dbcc56506f2dc9c33cde85c4715aeecedff3dc33b91aecbd235006100f1bb835b295aa3aac2e87afc2da4e42c7050d52fef4272d09ef608af485e341caf84937fb14904366589133fbbdcca9b542c20fcad42b5713d7082ce266121d649c2172abec6cdfa587267d92ef533ae81ef99a6853d6196c76048c93504ec5c3e9aeb10cf5dbe8e1ffe7dd4c7287931217336d4538be315c2a9d77cb12c824ff2f4f1275529aac04b35ae99e795f3d3599592d6909653d0da9648d26dbe20cd49c415cefab63bb23925ec361a09631bd939fe1a63371320109703c009d5633b259d23c50ae0598de40817caa73f3f70ad408573a26cfe49efdbdf6ba593e6fd65e32df0f5bf9fc32ec7cb2bd22cde2ea95088d55d454fe5fb590c447f02adb28b86620342fe48cd0a1295bdb8330002f536e4448e68cbf22f23901e725a8f4e39128b1ff0a510d214840d674d87d7c0054be20e34f36ba777a3830eb2920ceec78c45523db2f5931bd2a50826667bff4f1b8b89a77bcda46c91261433810c80e8d3565797e18127c670a029650f1e51a7961d31c1c0bce691eda25c8d785923444af02a7391fdc780e89ea7296f39bbb9d6c285e2e2c9bfeb9c04d990163000925b016ee8dbb8593e043a291c2a9403b365ae8e790a243895420daf62d83baefeb51fd8ac31ceded413c7350f0e88265d5d77eef6e3b1a2ff4a3d4bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6ac5c8cc1eab43c1da45869a8147450de20d7de3cdd922d6917699d3b14ead1bfe0a751c545cb79b2817c354efc945f42b83f95d6cbf341fde834f463474ccbc0e31693c95940b21440fcd4d57d5388ad4b3e027e7c03bb57756c0ff4a8599070641ac36773425f5fd1f146f4a31d8f5b2c02af88b2bdf2a270cf4b340e48fee915e6e34bcbcbcdd9a63a186680e8cc2fd50d624d9ae93c7e52852ac556f4afd63635aa7ca90751a62d320b62b8c288a8ae93938d36b01206c7fb2e17b7df3b4271fc3b7dfd6709dba7cfd25ebfb2e9d9f26a62a3acb151c991657570732a1613cd18713e4fb8a4331c0cca5c1c73d9670428f85a509094855a0fb404f8c9777d14b472b687e5797661ce95727ae8c22d725debc10f48e409626e7aeeb9c1de9e1ae27bf5140be5e65a111d72efb67243f446c772167c26b24f910d8585ab6e3714627da422f34a91e81c976da748368d3780a655ddac7100c306d999b8e91c732a4a67f13bbeac51b782bded2256ff5752c104e14fab46d65a205515d3a1abc3787da94a7c7bfeaa3ed8a96292cd9f5237c56031e654837a750796710d141d8200ccc61a4ff317ef6597f7912c6117e8d3220bcf6b94590cae0f08909ff38160a712ee89ef810af4f09cf7f5e68bcff4b25d61f580c271db2b137bd559b4ef48bc366a6f06d39fcdde7c6bc156b0b183c3fa4c6bc1647438387f4462af52c73;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5a8d7c01caa481807b7122dec432be33868caa79efd7787f760b63f0dfa7d5de0cd1f20ba2acbc8ed6e04323736a5e61655dcaed61a892b5f6566979c0f54471502d6837cdb26b231095e73b5919cab73a0cd6c3b4b895f86d35d3896d096400aa3bb92c46d02a46923eab3c8cf265d1dab708e184e6369a342a679ebb66cd4227d381e908c65dbdb56e8bb69400dcb7090c94c03037d31342401bc2dc557001c1869923985ff3b0d456ba4b813fef5682090ec2369f1d452aad2e17655035655248dded1077800aad875ad846cb11c6721ee3dd8003b2c1405d94c0c54d584bb8bfe0fda6bb18be1d2e5cb2ff0115462b63d28e74b5d6818acc76c2ed95ce4ed60ce82786636b04fd7e5111d566dc00263552bb35b3c140f24f237e2e65f33f2190d17ed07373b45a64997b3950dd631f20d9d09388a6754de79034426f8bd3f8b21771f2cedf5063adba194e7ed739314657b75977c0e5668d8226bf26d360f8be6ae237dd94c25f24846b03a5ea30520b30cca6b382a2586810bbda6c9f421137f94df51a4d35719000582003a72c847acf6bfe36ce137cfdca04d241c9319486ee55bee3e076fcf0797a61d52bd335ca0e9a4c17cefbe9c03ca1c50ebdd6dd224c46e7b6e0066a507fffb9f593f401b4a0f4e216505acdd4854ee64c9e3990fa1f5c44a7e8618330077c7c4cda0844e0024c7c4f3d53a8ae576a8b1fcc04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4891a350d4d8aed83a9cc20ac326d582a0d31299a9c80ad36aa155724f04f647dc9b58bf33438c40735d09f2b136d851ff2d6470b2d00258af1e133c15041524cf2dec16dc9d7dadda3c4780c977eb5ff253c312533517633b4a79b5e46374ee0e997f8ff796955c7f7c21df7e11b0253d9d4bb0e7a3043814c387bac4bf21696c59fd238117297ce6d2417703c704c7cc190113f6d3787a4e88be11c6de51d6c04304242ac2d13e40ec32dda1fe55d38334aab85efe417f31d493d6fd3606526aaafc6864610df692a06cf41127547f9d7891c2dc696f2626294bc5b96b46063fafdf1d9a8b189d542bb6f690edced45ecf5d369a75b2b46d7d18c0345407c6be32e329a1f16d59394db1797c479c3f5015eee79454ac23c39f7f049a2dc648d99600d42395c31dcd369d6988b05268c192a082e98769d85fb68bd5676f03d21bdfea0bbe9a24faea99bb5ff6767098bbc10cce435f4be37b5dab5e1821b793bbed10275150e2fbca31e9b4d7a8ba645408ce96e4cfffe0ce5d3ac86cba651f053a3ee7d8731df70c5668284aa955ef7f3c79b8cba22b0f8a758d81da36bfbec628556a130be6cb917f6c2abc2a1cb728f88089cc30e760a48b0590c82df82f015a4728bf38595dafef649fb900ba95d426ce998c45d0bdad2d276cbc50c357bf55a14ae94ca8bff3d3900eaa92f847ed77595881542bd85a8732887c3313cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h95cdbe1dbdfc11cef6f0c8b48ff9f87882ea19e570eb3c4722be8d334563b924268fdf52e6fc5e0e249b777770aebf9afffd2818739293f16a2c24187803c20231ad45429fea32dcc3169f3cec90866890e71af672469d14c01a6ae7c54eec034081441fb233cc88e569a1efc580da3d4378def924abc0003a7ab83d3cffdcb7e9f5b03f9df10264235846e70fd4514ef0b8f44e41e0a5a9ce2a0a783ff373a45acffb49783e8aa73143aa0fb5ba4f9d16667eb359e6b7a1cb7fc88721366375c285b3407103361d7a0f02baaea27b5c65c8187b96f59530e96273fa045f3205690995ddf982874a99e2e0bb044e064b50c3e2e7119ddb0b5d23181017fa3932a9c70563cbb552009866eaf7b7f641424df378de466377e25b4cbd50adb4333ac01155d2685d8bce4c3fb07e32e84b1318ff9902ca126596a27b7b6db6da6a1814d754e45f9ed7dd912ed53d6d439797d700c203974c2b97e4524a6829e119bff12bd4043074e919f0af7c0645ea0ba774d83ccbe3271e607ee0f8a90e70df1b4a3b803da69a9de5aa7f96c86aa206d3507403ab08a63b4a616b51d1025c27972ddeee150c94532012922e1c55baea958574d9d7154e9c7424477e6eb84bb2235687919418207f7e5f87f69580dd6db525978e9262d2e819e0d5b2ea075c620ad2fda63a91b37546687dd2a9d919f48294cb6afea3e929e5beb3fbd1095cd78e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h303b6017540cecf24d6e7c30bef42b5f031abcdab4d5dc2ee33f1d61e621ac6883ebdddb3b330b8928c4312bce34e12bcdfc7ada79c747d168931ef9678dbe2df2814ee5df2af566ae606bf98c6f7d8d588a1a4e63f29e52bcdf52902c7f59f3dd069539374d3de081e73622dd1f9c8497a2b834ad4a7fed07095fe7b72e3971b0ed885cfb28d6b761315eef8445fc840218d1f27d084abf2868b934b657eddd37469a9ebc80105b0f64f40f046358d379a487cf914002981bd5f2537b206379b5b6ea0d95f50340fbe9dc45267f24cf05207b6e8e9459c3035997c0a2894bc30739d7ad9cda653efd9391e2560ff1ee568066429a45a9ca22edc2459a98470939d35acdcc30f91d297be70ad0e388e9b08bb262fa7fc3abe84116cec2fdc338dfb2055f9b356fa4a8fabd9f31a070709f4faf349647db6ac4b300ed7e5b3f90dd9e76ffb8d807d5433436b7a151782702f6462641f884eafe7ec58871ebd6c88093aaadf9f58e2b3c640ceb3d80b9fc4e917fc50a350cda3d8e2dd2e0c1f39c5a12089a4607fde74503c0feb6e3c1b72a88ecadf38c4a32d56cadb2b0a2e2a2a5deb8781fa2ebdc06b8da0be6a66789d9bc1edc6904599d1760e76eedc4a9a01efdb8d420346595da7d4444adb6a1882b916fc74323bb95a4c0130cecdc9cd95334da16eeb1e55d1fe745e7a1086c1da91c81b9245107dc3c0ee1dca40c2213;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he222fb22a4875c97b00facfe2f8a512ddc535a0a9d7a4776c7229f093035afe862417bc4f07959c83f3794ac652e7677a8d5b37c0ceb68de60b2f6f48243c81682a5bf3ba6b1228e0569ea5e1d131578f8ab6edc980b92e5e6b163403c61c2f1b130819f6920071da4213ed04fb1b05ae353248c961ae7a83aab7e3f7b500e2daa92b64967e23cea62b5df999a479981a07ecebe8a8556429e4af5c5bd0152234faef7a0056b02a20ff97b618a5db736bb524a4ba01899ecb327a98404691ac7ddec2791ba7fb14e96a926992d86befd8442a2cd803e34bb764b7d5b30540c083d545929030615828c27af55574c5555300794544b017f66c7d38c931c4c170989e9dfa2b6ec5cd7b4793cc34254ae03c2c4451883d2086ef8c5bb6a3cec5bac9c3dbd9117fdfe4a18204a9254640fbf6ba71aee247e137b65b2d59bac3592f67125332a22acf5e08e0569f1de60ad5666a44542806f48ee52c359ce3aefe037570a222ea1e7265db3973df3b04310c53cdbc4359c906a75f1633a9c6ad4ebf4b0e8393d79167c0141f468a7f799b011602ea31746380c0f49b94e00183e370248c1262d255aa74dc6dfff1e890959101f58291cb8ac4d405eab27a088751c3fadb451fddfd2b038ee7c577fe023f2a1d06f9d5655c58c1dd64419bcc78c7c3acee79a397bda95ebb74d5db723824950a83df1aabddd7610fe0cd520c7e3bf4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h766da97a4be23ee61c911d44b33d3de612e116eb134dd00de324c123b31d96eb9b0d2433f2083305c4145c5cba278277cd8dcc30ad63fb78d841c63395d6b2935d1a76f6dd23935dc49e3d51879e5ffa08ed3d87cf9d54978cfcfc9365c7dcc1583b60a1afdadd0cda492e7552455e0991f630859002e6a32480ab269ba95f8af8535f910999e4cf940a49b8c9fead1a38567507eace71239f4fd2f42c707a2c18c2652af4bcf0d761c0ed7f7c013760df20bcc28ce6e5b68f90d7b8c6a4b36133f179408d7ac2dbab0271192b8d0d23d94069cad7b6b23d1315737519b782696669c96b97e1498fe04c0ab27d368242338b4df58418db9c6562c724ac575611246d329c3da644e280b5b4b6f04cbda7dba66c6a49121895b56613fc165541e2c5b6a32937b7ee1de10e4433529a7b1843b083d525fbe78bbbdd6c6c45057ac191312d28e63082bbcda7b4050321d20ae0e9eb4b442722a1f92795237eb880c3c9b46e8a63ba54fe18a5f4a103a32f92a037c4bd07727f1d451b76a96f322a3627732760463bf579c4beaf6fde6522c7886317d7d53e943422e207f23f44c6ed778ec504503fdb421aa919d9058e2aa4a90857b793600ba1b08d712003d51b48644747252e5af448eec71a0494b5563d3500f2963eacdf0d9457dd696669b2eb380b0d68bd904be24c3dcd7b016ae19119f9a1fff95cbc8b0831e0046d3cff23;
        #1
        $finish();
    end
endmodule
