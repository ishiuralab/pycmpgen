module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [21:0] src23;
    reg [20:0] src24;
    reg [19:0] src25;
    reg [18:0] src26;
    reg [17:0] src27;
    reg [16:0] src28;
    reg [15:0] src29;
    reg [14:0] src30;
    reg [13:0] src31;
    reg [12:0] src32;
    reg [11:0] src33;
    reg [10:0] src34;
    reg [9:0] src35;
    reg [8:0] src36;
    reg [7:0] src37;
    reg [6:0] src38;
    reg [5:0] src39;
    reg [4:0] src40;
    reg [3:0] src41;
    reg [2:0] src42;
    reg [1:0] src43;
    reg [0:0] src44;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [45:0] srcsum;
    wire [45:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3])<<41) + ((src42[0] + src42[1] + src42[2])<<42) + ((src43[0] + src43[1])<<43) + ((src44[0])<<44);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1175d9915c2073d4a1a9f6bb97584bed8570b47790997add6daf37b8ba5898340d8ab2777d8262ee49baa6895d23ed4accccf376604c7f4f001e6a1325d1774a20926;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182cf054247fcb5c3bc28652e24b89b154cd01e10ba43f7a6edb2ebb95e04746b7bc847fce78fcbf067c68685abbc5d7f70c400555f69858133ea7a755340bbbe58e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec1fb81a614ee6e324a1bfa4f4f0fa2e753a084321bb2cb447d51c45cfe7219e265c863562cb8a265a94152b8d11ae34055d2727e3c58d6585c3045845593410032b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8e12e21d6a08a2748dcd9fcae8509fa1813e85d239e02a7ea72b92fc404af319709451d8891213cce341cc5147a43f685e5b45d75cddc9ba4e73cb8ae547596b5f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7834047192e344767016edd34097fd5c89ff80da1f8b6bf36499ee59baee80440ae7bb052ef3fc45d5fad49b8b5d1e3a6ed87ef68d15e2cb2e7a308628945836e63;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65da2bb00cea01338ac2369290bc93a9d3e26d9d40bfdcb6368c27ff4ac5975559fb7c45a64057776db53d36888d3c3b0db6b4709e41d368a0e6036fe4e9d9c6142e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3c848ab427092ea6261322b311d2cbf55c558f8b89692d1abf79f8db7ac8ca30bf4dfc2de9cbb163e87c52c4443ed63f68e9f20a289c37e9a4338a754cff8d4b733;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0eb6f1e379880dd0dc73453db8e6bbef5f559383389a7bd9a5a04b13fd830f3a5c494c7c6a11a4093b1d40d30789707d04c96cbc6bb9185ede7708810354a41e4b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c96dd798aa286fee76769e95cee3b726ec83e1b307e08c7236a21f5526bb1737aaa809afa6c9df4c08ee68b28b8055d996bf35d97e413d896e2d2b7441d88f68ffe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f43772ee9eb7768303ef951f770fec2bbdc1fa4ce5ac8bbc92bea1b80b8bc0b035a5dd69960fad7a560b1934864795a9f7b7f9d9be5b77347e2b6fd44dd8a28d566;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d381314dd7d533671366e3bf23499d3d20d9d78c5889c09886a0b55d66310542481b303c5fbeed8a87f095ca3af8ed232ef49db4b0c51781a7c067d85fe2929736b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24bde0b1b891fbf5ee7c64f117ffd6930fccd258f6c4b4c4a5ec8afeaf7d04a88712b7ad0b162678aa589148f95c8bed1724c3c9a0b18fa38001f7be94ce6b7989d9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2dca3c2603dfaf8d4e939cb14a2990666cb7d96ce5fe860e51db9b170c7362fb82b97c337d23f9cf3ce306afb6c6baa26732793f77754c76ad8ad26df73ff09af364;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h149144d00f18b291041260de68bebf6891dab7612372bef70a96db68b5d48edc1d40358b4cebcffb26fa7d2bb4e9e4f1d57465875ee2aabf0490ffb07be361a8b1bd7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e1e12f5c080303aa18dee9b46ab49d713bc433bb38ecc0b3eaf2bca7457284e5d3cde2e7c935bce938219b42dfa8c261867a7fefe270e45835fec263ccc134a72be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a59a20ae3c3d9ecb742f853b744e60de26757dc68a48c5b26316f1e533bc0ebe4ab7673b899852f0ef91d93b808c6af2ec55d0548989febae3ba98c5c88aafb9b44e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47b273a38504f7d17d0c20c6884c957274de49d6f8262a485eb05dfabbd30b445e3240b77ea815b10acf06f8632db3ee992db085547489c780e6117b3d142485f3a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145e9cf5b7c148d30e5d45dfac22e0d6821efd3e33dd1c7cbbd9e36c484cfeed639bde6c330ba835de75aea187308de356a77d8e205a473b7980e2248467f0b6e2b60;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb85a602f7f4991a5d9a40dbe53e11fcc5a25f408b2c2a9a268bdec0a692a24ab668e5bb62a38056497433ae2f1ce1f7606bb1ef34e54ed929d5d18a3c97d7505bc6d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174bfd1bd005c6ecc90dc71a261f4084c04e7f04a936f3b0b08b56eb4df5fa990dbc80f4b3a40ddcd126cb3462dd19fb922653299d944935a50d3af17f92e9fd758d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cabdcbd29c5e341faa703f4bdee22b1dbae6c91bc19f86f5209256c98fa79271ce904b582c877cfc1c72ffec9b65e75a3f3251b20844a9daeb7e51d285b4b429cada;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f22cecb09454bfecd9152785bb622e4ea06ac456f2cd35bf441adf1fcf1550d8b4eb36b8916a8e7c091f57bc8c3d74b5ead726036c05d8aaa0a71b2f110e73832a56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1565f5cf4118dc34b4b13dc28ee452b12a46523820798edb20d7f4c9df8e99ef816788aa00a7bfe472f81a28d34d4ad817c5ed925dcf469e197800b590fda32838f28;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4d2e767fb45b345df693fbd03238c19854f67385d8f18cd00d4a57adc1bc384743cc4cef0246cb82df7d77400c6c08eb34a7ca945fc869c2c97dcb5a6c48909b9a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc8bd63d501dd8fc983c698cf7db1f831f32e9402401ebc1b290dd9f450c78f91a8b2e927febe7895d1eda596ad26712f8f627d5bc7ff79653da9549c28ce69f1f31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f4a32b606644c49fe1099c7755ac9c400f33cc8420fd6c66bffa157d78923270266e33d3d49787a234628523107e501037065701c513d3ba3cbdaf21355f00bed0b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c488bc753e90d6829320fdfbadc2b29ad15ad2e2b272bd05538d1306a444c85d9e02777b4330d776a510b4b199d7c2c7b9a15f54d6a7c18451a4d192765199bc414;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc79bd20be5862c766941e1de1c2c3550cbe50f3e4da2616825e9e71c94730c643d23a615de081aa6d54ce450fc289ef688cffe60176af4d193a7bf9a776dfe5ca7cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103f17eb2dc4ad69689c69edc38d979aeda18c5ad9b8ca98203698b5f916013bd4b08887dcb40b7f79d7709ed8ed71b0ecdc931d10ef2a14c7fb2e7dd83f6425400c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he895990689586316fa7dc61b27d01f123c68a2173c181aace7ba8c8a22f8d58a639a0b4608fc54351d049c6ad3f1833867fc924594d5bec8714e517f7ee684c52aab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2875f4e33117618270c2b0186cc4c9384388c713c3892a62440cd201ffec2b7be08824884ed5164e76acd8c2a203e35985a9a3d66191a37d0934017710e16a3c3419;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a33c605a8758012aa15e56ec52f90ce06a1c1fca63c3f1867e5c42a87402e8763ee0a040b879bac89ab6e34ddb163cf0befe548e3b57cac8d790d734a80ab6e562d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h355f7a30ce6be1ba469d634438b23fa72fc80f16d07eaf8680bf270be57185defd565a80e0da3517599639b1d3c52b0eee7a3ca7bbd72d889afccc282810b0f2a3ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15eaa281840ee4f88e1425d819b6edac07d80fb231fb1f2a04de534a578bbfeba710b3518e4cc0bb588f768f379af36c33126d9d51a55afad24bfd5ab8133f3d0cda4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18174bad11b9ca63265ddae221c02fab4b4770982a635dfd2a9dd007263489e0d478bb02bb86ecf2fd82cbabc963f3ff716f31a890a49d555aac0c86ea46d6bf6b087;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1901924213f9497c6d28e599ccc088efe4d197eee9fece64bf0a4ca034297f6b25885742e0f12845e0ad4941fe4b46a1aaffef3a7bc774ca9b32d87ebe7143ed8935e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d591d84011538a4ff964ad1043e579a038bd23833d6c3069414debc6abe88b30757d12ffeee639e0dd2f46832ee040247b4286363e5411ac7638aa734ef28518e2c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171661f32f83e93472cabaca75aca00361019a43eb25f9bb9fc8287542295c6e65bd8f84171947bff98685ef3d79080ef60e684c5d2df555c1021bcd10b536e036530;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1831355bf1536b055f11727ea35046b8124e7bda73fcef669a86d1347f57a2fff0e4ad22dc4ba63f7e816df42dae3d3f1a78074c8a289867660fa0505ec06aaae061c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h686098acd115d4fa99b58f1fadc1307c575e52545494a9db479aafeaed9e1b0ac1dcae85a8ea362a9e8f05f14af02d9e43659d9a27c23b6e6d48a4b4bcedc9aa4dde;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fa7daf759c152248adfcbda9e1ef43a3ed9fe6bfe0a03c8c562410dccc2858cfc41d57ce5fac039b93357b2c9fc4564b0566fa4082d6c284208d8a1f57162a658bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15931f30ef976fe1256b72d07cc10726cfe5e114be63000d796c45f727dd4cdd64334521e18f7a693729f9f39bd371af419525a8153dccaa47995b5790a4c8fea8fbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f243196774bf26ba403c508f0d225f6db727057850b03bf58e094ea47c85c854dee2648b8d8c863b36b2679983aa45de967dcf512df3d97dfa15157ead99d3591a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1932f43bee3e35a77dc3fad48c22f6ebcb531e68dc566e59f503dfc4c812da58eb50fc02b1874f99c316688bb70295afc7527942eca72d8254a46095719e15ce36762;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27494bcf765c72e0a0ced011db42cca084c50e86b10bac9e76ec7d62c132962c8045b47d6f13cd8434f89370b7b02da9090fe9b54333c6b84762d8cbf355d974e343;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2aa7d8229f75ff96e490d75971aa85230b519e7a58163462736334057a3d76c4e34642ec122457928bc94b900b60d8f13f2d612075cd366ba820a22c0d9971e59aa2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h601733b5b81a1f09de1522f181d7be26b0e59411adf8e9b13275175bb644656e34481830c209428010a35bb698b6d241022f95dc28d856e9598918d3a46a3d54eb10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc649aea742a4bd612a6e6e7a23f1d45ae473523419cf4a2f08bc4796d170fb32e6a1f2fec5c531fab14ba6c557f87d863537bbfd7b3c689c5ac7129e4dcbfdb339d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he90b6436053336a6005a5d570659e09dc6423258a4a4248f1c2c1105bf1fae400c2a4319c18ed1041759d4e1cd64420d6a2a971795aa5daa2f486ab20475f5b983fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h183fc747fca90cd969f17155ce509956f19fd4afe49364e49750f02c1af1fb898c3798203e7cc23a27b1eea808fc306607b59b7ea2eb8605e001b5134cefdbef1ae1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a97e7b445ef44b07e51848ec71565f4a6a817512241145c164aa16fb69157999f59efad08aeb23f31cc83bbe05e0650fcbeaf0794f636eb0a3c9092e451ec8f2e0e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd19a7f3fbed9e03c219e62f8a83f46847adaa33a98206328ca8386bfbddc66cbba0fafa5f52454dd1d42b89c0e7cf542562150534e0395f02cf27f38e8fa664e54e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfaa6c498a1ce0025e7a518a757f50522835da7904c79a6bc8956799cdced5da4561e515d31d37ad781818dae8582dbab09efe2602d67cbbf461ac16c9d7cf344aed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he384ed50537c71cb06b883e3ac625c86953a2cbb962ea221dc1109e0b5ca913d0e053cc4bfe417bdca9613fab8f99b2ec64693ed954b33f9277ccbf148d84cf02692;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11d57fde2af7c23db553d4123b7f082dc74c1f31ac499b257aca5730317618c1496b9dcb5bbe6219909dc26d5d18ebd6d9b556b23d62b0e9081f96c787457d66a66ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1375e4ce51006dd0329030b200e55269987e1b3ade8efd6e2aec9e4aaeeb659e3eae8546103581185b89582b1b51feb193b626dddcf6d2e0792db7885f1e20f9e0bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14516e66c3aaa55c84bb589c1b6fab0166bde0fe269dea9c7353f550aa1aaffed23f6665e46a00ceda893f0c94f26fa64e9133564d6f70b63e9407f2875b85b31f1c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h122da513a64ecaef7d5c3d49307d9d9f6c72d834f6a49b11f9b9437218a8596687ca742b091369e79068ee418cdd06f5a22cf9688c2f6a2741935700ddf9551b140b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haee4060ad174272f6373c1df3d0a3115e6b6629b38aa516223a909dd6201b6d18b718edf9afaf080bb24efd16026a8fe7da1d8ac2f4862c937282510aa0d7705fd09;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6040dbe559fbf77a4b7a75718e59a5e2db920ec991d87741864db7d3f3e688bb8ba97d072982561cbe69c9a65320032afcdb56de641f7b57ccaba81289382e96b44b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f5bbc5044af9f415d63e3fed80c6e93ca6aa6583d8ddd5267856bd6eaa76b3579305bcf70d59e11fd4ea87cd25b96548e4a56be95cfcf6ff042451d2ed566acf84;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5aa3451236c7383c0ce72381f8dbc802098b8350fc354656c0e4e41661d9737741aec888eb7b2f6d4a2a780a4b5d188ba5db48b14f83f7aefd69bc4cbd5bfb8b0c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83a4cc1339823230cbd8aa2ede3be234ea2a3bb65560ede64a265490605a25e80c44b6d7bf8e42bf6ff587c5078c30255f72789bc907ab381717d78b4978043c4021;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd6b7afaa2c6ee8bcfe6f4498bbf4580ce22685bda38e15db7d0bdc73426c38174eec468976fc1a6ab716f33b1bafdc386d9982952fa003890d9c33ccfbf0694e3a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfafcc699de945e26df5262ebe4ee234d444524384567c7e2891bb9525a4bad5baecf4b9fb19a74ebbd780a91462f69f607beff426fe25e8dd9f59a0faf992fd74fd3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f318058c132825437645907c691946ebb20e1f3328ccf900ab1219a56eeddd0d8166875bfe02661183bccad805072d3dcc479daea6d87efae93df47aba09b020cbd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186eb162aee196f8710adcde6bbe72e46f676858742ccc9ec78b3955f3a21d140a5954bfec2a939c7b329ceb58ca083285b50116419548607dad253a58b55f2755b1d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffc10a6f3a48193e036793118d36f8f22676f50489a7d5986f9aedc5d2897992cea77a77af13de655ccb55189d197d85a6d7976da5e1d84cc7ad7a663db521b3fc50;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145251fd597bc812f6faaf28cead50ec10077de6ef1acee97420ede1a3efc4e4cbdd8822ee2c8e27aa93594229d27c903b8b79885b0c38ec966bd204f9304b1ea70b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2ab81a8d3c90d222bed5b5f8fabc10e50a02f886bc6aacff621db1a53c844b3abe89ddcbedce6cefe62c95ad1e6dc00c8583ea68fd55961799124ac29826d9aa7ca1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13dcfe0348b9d9ac65c62f29f8ce95d968a5a4de7a154d8f40287755ff7d98f924911618459395db4482eb73e5db88751a93951e3b10158a15ae255a6dbaf0618a99f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d9780ec86b2fa4ac741255f952c0c812ab94a6e4ac5d6f424a04a0596eb5c9505f0f5b8632cf9c7f207d795fa5b125a6d912df3ed7d40ccddfbc278eeef2e777f235;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ce3c7125f411d1c993342652d657e1fa345a59f8f0b852648b7a59ecef7fc656312b5e148cec7c336bc5cde5630746b80d021ae35369e13ea827c36bc9d1436f19c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h370032b29e8fac9a6434eb6b9158fd06a93c43083f0496a607f092eb905d4f300b66e839b9b618a0ceaf8dc8ad46207215424701de22963c7cb6545f39fcb40436d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h160f406b536b1b5ade77ed3a5d5857043cad2e5ba06da66df93c0368aa67d18450021a9a998af583729a7a697905620abdb39b473bdd310cb3fe4a7bebab1465af535;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h206abfa2ba239d3dd486963257c165d3be458992e1f176b45385d09ef5623b62783827eeab91001e78a4c925c3549bc9d92515017ca816d8f80996d269633d0d1f4c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h191a452e625ac51fed357d5756b8603b76d5ab4b2b7f3267e0baf78124cc06eb03afa492915954bae115d299adce30dfe1f1b4a8eafbb94fbba9f289f228f90888e26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54744788f020628c5c238f9b732ab774e624c509d4ceb102968843dfefa11a397f81a49884944164fad31d6b5e98530a3ee3577e3e26ff12490f2c6fd86298bc3dea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91e415fa1a9b8e297370dda94dc90f0709a1405410fb5b00d216dbc778ecf1aad18591b159c693a2efbd79bc97da6d7fe85020f65940f0124589d210fc65538ab3d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61b7e6a03719c971aaa52471149e1d323881bcf9b6239c3c2caae694b3314fc40ec4661d83e0534f655f5b7566750be354ea3ea2adbd76992ff11dde1e7518ea4cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h195ec5b869a2656be7d6e0f3e2a25eff58d0db51c04cf98885b48200ec25fbf0ff097b4bf267d930f91a750cd308b1167e44a7abba81ed4f832caa5793b6ffcb996bd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a57a4af03e4f53f32e3f098a1dc7b18a4c9a4f60f48f22f71442d385629e81a424452b3623a8637fc0855ca7bddc5fe190bb4a415026adfb9e5dafb1f49fd1cbaa81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1196292f8789e84e6ed3a6f43d56f26ebedfb3a628b96bc796e82faa5576c98eebbd2a7d5fdd3bb91df49085d0ea850946338d34371fb0fad30396d682ea27d967411;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9eca09353239842e09060dc063aea2a02319fa9f44c4cc06885e2ef6a4bf0273a127ecab905df41b97029f43692bb21f20e2ef7e4096e71d2aff14e8f4d728a0b9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8055105c5f9aee21191ccb1bd8e4bb308b9458e882ebf631b3bf0d98c979c1eccfcc576f62d133788e88b03fbcc0b965b2e0efcd0e87fd2f6e00781711b27c78d7bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ddcf579e3ae005aade109e4d9aa0934cf8e1e9672766a21066697cfb0e0f52760d20ed80a8b3c404785f0584fce6eade3718e8a78d9e83418dd951e2f028e3020acb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110238a7ece604c0360a1de2f18c6b13b1ca22640127fd9b0056d1d71126d41b88ff8fb91816ce089bbb3e8b139cc594851bf04f58dfa24026f96a5791f5c17149957;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6a5b4e0a0e5679fb08b53bb074205c6cb3353eea396e1f0b421c7ac015b25a376c8959bcd1178b3c55369bbac8fa41cf2a6a6f71cc2874bcef0bbd9098b301bf4b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127ef4fb83a7a7ac7406f3e7f0b57c282c39be24480e99aaacf8611d83585d0c133b9d528b284d365fe6feef64150c6eccde440b8ed5a1fd1adabb478b056699fdd4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f73c802d840bfa0d4f7e027e99c1c7b7691b961c57575b2376b89b4b9e16e1f4f15c3ad6845c6faf21522af27d4ac6f02b1ef53f26b4e20ff3ce3d2a7dd02735637a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c3d30298ad61db215892fc9a4c25dee5a8c2a1c5dfb03163dea76351468e0865f0999ff4adb9bbf4dc97424da2303fc688f2ec252506a7fe983dfb88e9d02d13ac55;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h334966ca0ef502d25f6b29005fcd1cce0861149d0e437ccf951385a01052a088215beaad2003506bd8c63ac00e16569c01f180df0a0d56350f131b249b2da04c678c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c910a4872f222600dff8807f345c49f9e7747c7463d1a828426248bebfbdedc73fdc37e53486e95fb78446495c30828381704358f6e90202e9d202b8390a2c827e29;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1427727b04d43e3c2764b4dc83cf736a586979cff0a66f9ce7a5dd013c509d2d2acff56b5980284a793e98b7a6752e9bacd388d9531348f50dbcccebd39b285d28559;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1301b09a5a787cfbf71ec448fdd1361707af032c07db1634e89ca5f156ae610b3bfbe42476ef3eb50d8855b48878629ca553071a63ccee73b37f906565e91d21633a7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d1651f5f5f89c0770eba423c4568adcb27a2fb2b7bb10fd6ef4ddfa439211f87728ba25814f470432456b3a03b62aaa7ec3d9855f910bc63b9e647c551377fafc182;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf5699f02894b8bd6519f9208332d88957afb07884d12c7536f30cc3327bacded0f18f27178750ced7d1fb81204369eb11013b31d1e8c44ad836334b73829e85db06a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d924f003bc540face0e65820075ca8f12cd402f21fd8c3f7a60d0aa95527d20ba9ed6707f9dfc30cdedf766adc44498bc27c59746c8919356c4492e2be7b80c6da61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73d3122dd73bec5e5697fa928544b54a166e3f6c14ca6f82fe58435c97fe29574d23394291995fe203a88f6f693436a5a4e26a5ddefd2abce0da55da5365398b6642;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c41c735a87b1e29289a1f6b3627390922d89bda87fda458fa73eb65693ca0a31e65b3ad238447d9b8f4b98707bab4f1261750531f886410931ba5b4b1eed1ce5a733;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe711320436e3fb4f924982f4cb6a1ef94999f59592d37a7352eaf3b3f135c9b6fe56660a44922281576582b46a1b578198af87837dfba23ed0d0924e423e1fc855f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb080d3fd135b79ef1234bfc2feea8e29dae0f952a01a845c8e4825166e0a729f097eeb9a1037edd35366e3fa9fe7408e9ed5a26e5522d84f60fbbba1fb30c1fe2ee5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha382df6c33778dc913955074481265d65a3709b9b21e4f0396f3a049fd5030284988467b4b10f31fbfafa9b86c550475682c76eb1bb16f551121fe996a9598346dd7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19819a11473480d092b95378f1e2061a88af7fcecfac8b74959c8b25d30df23cd15c820119557dd644d30744454339b1dec24c0ee901c782f8cbd11931790347efd56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155569cbf7c8e4673bbe471743b39d837fb4838d4c88b0b3e1cad0a005c4d931fd78cb65f304bd6e9b96b878fd781b2a5ccd5061a04b34e7a193d3ae98936f4971888;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc22e1a3c01adc3a7dc2057422c1b3678c0d2db6a07a38c822991c680b8ddd89bb1f1f2dfa18c91eaa8e40a95eeafaa67b5d413f87fd589c401682196571604af084;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10edd0340cac06b8fdc11a538efe6541a15834cc7bf3706e1a7c64f5f2a293db0e0f498d552a92d68d3330d0240710c5c2fcab30829174fa328f7ab2b93e602b29a40;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h375c89d7558508f9a237971d051ff513c7ea9aadbd9f9b5840123ee05874ea5a78ed5c8cdda68739e8c3665cfc05e7d122262b5c83f0b9afb96afde32abc422e640e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce320efa8b43696cb1ee5b92654f43a5272ebd409c5e628b7995c20e04d2f3a1cfefcfec03652fb8495e91429c6f6d7205462b6e850b9bd0be55f710265d9dfb584d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h158e1e3354bf310e2ef44f0a4a8b738f59e7b7fd9a5c32308a5c216da488665d7cdf7aa753715c0bd122d25851e6b08b23b6f11451d462c47d62a26eeb1d0e8feb2e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h504a044acbfbab81f6ff381efc460696b53fc8e9160ec55861483e73dbfdaa045691c68be89932af2145754549b52a0e0cd10419b6e4e0f83064ddf89a369a4f0c21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b719e40052c6cc0ff6c90bba1f1af57135299f113eabf72b4d6a833cb3614a82427dffec8e91751820ec6d35f352226aa551af29e8d3fa176d34e05eaf220b55cba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d3b47d717908ac1004bc605bba6872d9d6149ab369194a1a98cdb6dc2248a7e7715d1ba952f1b004a8dea2cc1055363794596daf0e192b17e3b42e8cfb88ac54986;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87cf9d454ab305980065777c24907b83f969757f2ea8be0d4b5a53c487ad32354dbc14975e15ae880178848dbc2285d074122924324c81bb3b4de46494ebfd723766;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1787eb6a5e9bfa8528f9996c4aedddcfc8278f1c89ed512a209205c14cea1a81075f18936c81bd9294e1d9275eefa71eff535394e25c350a7e816fdf535befcb965d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ea10d4b3abca8068b32d31b78b9701c6c48b59810aaddd3ed846dc52e5f7b54a2f3239de7b81762b685d84787ee0f9004d109a5cbe5938e55eb3cfc2f492d3d78c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h84f8121b41d997692b2b9887914d7d789f4dfd13389c16a06bc5a21fa5ad42e94f3234dab6e3431634d81b42dc1f8d263810b000f6ad415deb085041cc615da7a7ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha2f6eb659cab98ebfa4ec4abf70eee1c81b5ce08d2374aa594a963884e307e621621d93ae93420c8cf9219ebd596fa9ad78f3d56c0ddd7529b799d7c007cd013caf3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bed0db04fb9d130845b4869e30ec3724b7709382c3fa06ab4bb579acdc9a53b4d766459150b878b5691c3b4a2a954915a4dd6d563fee9a6ded0ec220020a3af3da02;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15822118648e59b895a4c4bf8e920b2747f2a3c1e333f5e3eb5cb2d20566678e2f5b3bd43825acdd6e8db8ffc7fec4e8d977b7e0b079429fbe5d946180c5126ce49cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc05d219ba66e4aa62e1bec04b6761b523e109e0dadb8e63564568adacf47ff196c3983c74606c937757d7017ea453304c20d7c3f24884553fb335c32283ddf337ede;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b492757f889919602435a6bcd5e11c25d940cea8139c529574f96c125762ab5a268681bca4b9d1dd9d6dcbdf7ce2bf912e516226a8b4e21eb5a3891c20726ccf213;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cab587ac9e769480eb162440345efc1373624b3227b16d6befb85bd7efa0a4199132c9d08df9f985da09f2174759acaf907597910171e8f773c2531f6e838c5ab444;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h332595f097824cefa5ed8ca960d9997d6ba3f12ab26e319b5c93525417fc1f5e5687076f340050e172217b8c6bd9d94d1128a35d8a6fb3e89bfba74b26fdf20a8823;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73098616808fd9ab91f8f72af896935efb2833eced36151431d84c04a8891961908f51d5a03915c1be8160b65499ba14fa98cd7202f3d26e42b70026196b3aa37fc0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12d50075c7d4785623fa074d478577e3e65c519e1c9a3f0c1665d0e110bf4c8166cecbc517912a65103b4b6d85fd88d9e645a773049dba66683082fba3ab68caca135;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8be8cd38ba841bdcd5819ad5df8012396097e3a6e9ea44ff71a6c8e5655ed5eb15eef32e6aab1cab290f5f72fbdd7d0aaf47967ed54acc6e6d0ae31ff53bdb4249ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d069a2d9c631fa800deb7ca907c0c6b41cf92566793a9c93f8b7016ca6109e75b58d8bcd5735e6459215de2da0843c3896519805c648a36dc0cab9a86f2e6bee755;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e582d33454a7b903b79734feadcdc057487fb179f104895a04397acc02aaf8536d847613828e691e7295725ca83afb86f434a0e2cc06b410937fefdbbd144ff947ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h20f6da569b0d524d5c6e5bdda72c2d1f9b05442635a96829bf3e4d945770e1c732a097c2e76362b9140d9a1e947f0ab30e53d4d60c0e0bc4b4ec31ce535e48255425;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he60612a2e6a59e708f38420f256fb3aed62141747bed21e9766362c61cc821cffc769bb362d56e437f9976bb345685339057e5bcd822472dd2a5fcd99d037ba85bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5801b3e1b395acbefea2c97e17d103511e3ca6685669db2fa1343fece035cef9c1d3bbb2d88a47190feef499a9d59e1e81101e623e00e342244b540eeab7755abeb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a59534195b7d02bf8148f8fd2f06fc39d9e8b947ce19e99b85f0613b14f741a1ddfb94debd153bc2b96a836651db2f6735e439b9a3620612e1b5a752e59e436f956;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139c72bb21923a69c3784feddc18bbd6ea17939a9bef5e1334d85306417bd8373b0461a1ee17d31313e58761794301b85275e7ad2efe5ab30599988e13eee97e85692;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f52d0342413fb821414dc349c25235c387178ad33692ad02f2e6837c2b41cdeee71d254f87d124ebddb6cb5dad7200a6e08c8ac1c65ff97cbfa8f3254404c8b0ede7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf837b88e5b2e8b03eb4b8cd77c314fd58b1e40e2d7d3d379409925397050e26f57fc45f1ca50f7e292b781f8324cf6cc7da23c69666f6840592f66ba668e86d384cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11fc5e6475db1768a90edcbadbbe3e7eb6bd2c4bb0a4fa730551fb1ff28fb266cbbe0a635f64faf2b9c8bd69b40833f2dc28f059d36dab7388d4d4b11239e1da5aca8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c10f4b9b63cb7edd83e7e3aa8d2b0f3d575e412f81ee66dd1a44cf61479ca3dda903c6f852ba720d923d2cca73343299c8dc8b219b5b6580764b2ffc1f10c0c4f97;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2d9d74a924bb17145855319c061de993f81689e550185d05ae94342e367db461a9dc6fb37fba78a0a02f155809f33a56a3355c0df2a7b29368d7876f81df27eb163c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129dfa10cb2241d818db41960e8277879a7001df00c2eae19a95237d2a707a778e77b31e4cbf1f86736f3d8b0de3c1c5ced841554fc4ba41388b4ba2cb2e67e211569;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c5cc64e0bddaf0905090e7c8c854a2d8fd038781d617c14a96a7afa0f09ea79e4fda6c1b2b8f862077cc7714b882fff8ecf903a40d1d6cd6671092d2567b67a79e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he37e70363672b1079012bb44fa23537654003fcec617034e148ace3edda081c3e898365dc86a2d30c5a046c9952b0b4eaa1fc9f9b2d2b2336f350bf10c766d123bf7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1573d43dc915476b40969872f216e677faab31ede6eb6dfa64d1fa67478f3c161b843dabecabc384062f29c497485339a4e36743c34aaaec4e1b5ac5a8fe042f09dcd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e8d73dc7772e519802e72413dd502e4f4c5023021f765b3154fd207e40b677079592ef737e3263795433e8ad7267891497d31b846596d729196ceee84d1ff26f2e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185cc871cb7626409af35de7ced066e2c5e18b9cbab696810a714c96af8e8757ca647da431c7972155ccab992c8df7ea4658414832a2305ee36b4b8f93e2a26852eb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fabab7b677a05101bd31cd3288f3628bd3521072f06c137e840f834ed475d3acd70e5665fbcfa9989e8a82ce416aad6b732a1e0277c6564f16519127c410dfdc0f5a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a57913185dd9a3065a9dfa9ef2776d67bbef919d145c38c271e7ba8c72bf404ef186a56c075fb36e4c10c99c3874764640d86c664c518b40cc547706761856e1472;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2bfac7fd7ab3e6d05b8aee239d88d205019c9fbed027ee690bba7e777c8af1134d4883b180c7ef45296801406104fe4ce1700431d4cc8cab60bf655f57ab62afb7e5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haa2473814e98a9fb7dd042164d786a928e1190929ed6fbafd5268ff622ed75159b2371f9d471e70110048a152a3ce54a39da61e05b2e33c115ca70020691cfa7fae4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdbf4fb2a5da333fe0744aa86229186ce4582d0176e315b3aef3757708d57d51bea0aa69b86e136d0441880506ac029267fd94ca8c209ccf845bef0d3ec8995fb17a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4bd2924abf019a37b7d12344e2d39166145890ae708b4f01e41d0d6dca8324ada7fe5e975b1447e4f77588562248c397b086c9bcc2c8ad92f9f03e57aae177f9b1bd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a1158e34dd2bd2435c403aea87427526eda89013381f90dae0f5bf449846d8e1032007d5e8dfb799edae3fc23d6210fbaad58dfd225c13564938bca8cca70ec8200;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha263b99525262d909065b8e4262e5fd62c04a69c444733d7434abe26b6d41f3d95c62aecc1b4fe4c940801863213a696b1692f5dbf6a7535039b57421b52ae9d2ab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1569fba3b9f38420253d93bdb1f9a99aba7ce57251308d00c39deb9acc556a1d05f489051de5c2a3f226139d8414185f0c828dbc78dd1d27aecfce502606fea54aec6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf029c434490f19bbbef6189d065a633f4964be80cd75487fa418b9182657d8b4277c8e2146d99c20ede1ca4910e4613f11b4b94e828a67d33c5dd83089692bae781a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6c02bc930f3edfc797dc52983fed7faf782656af2100f0b024b4d99397d3006008334e3a99feefd32750d73347ac3a336aff01793240e40eb6fca83e856f9d1c0d4e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb8e17e960d79b6b7cfaae26e3f0d3fde4170b8e295e8fe0dd93e14b46cd80f95029c609121838f5700afcae6beec0a51da33da19bdf815bda2aa12ea70c1f8b20c42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93f47adb26314a314c6dbc4c2a04d7c00254ce8ae4032d76a7917c0b30ebe0f2b0c1f6a4246639cee98dcf50dcd7d16cbc834b98528dc0c8bc57b45bc0371d808b3b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa2537779d8b4ab815326659c841f7f497ce46ce22670af1b91d0debf3ce937dfbe9f2efd64077931db1aebfb5aaefc2c72f7d885cdf6e29d7a20c0ee6a00d21d4a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h97ea2757e6838c63c11f38d8bd38446cc393499915d6f4e257ae6f75874f1e5c21bdfc91e18609ae3567235ab2230a1c8a228df4c747cfd0c27db45bec004ac28ea5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7cd041c80b379515faf35ffbdcddb1c838562c1b426299393a2ab39fd7aff2eaccff39a66f7277031aa177fb54fc3d0557287d065ae235aa97478f613c4d19a7bd1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b88c731297ca1f9dedea6d4560cf4313de18b4af2f2a41b4bdc34709b36bbbe84158d49648d6eb6d86e22d1dcdff13fea9c88e7872d8983c656658bc366f24021a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7412f1bc561115cd51eac626e511edbf1bdad50bcfc94150af98f0885dd984f7cab3f4d14022731a9674546ba7cbcfa4bf63f2874346d3ee11614d8a897c518df87a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1168e47bbeb73c71a4f8569c5f9d39827d9dc394d589bb7a33e8ad1fe447360e8b4571416c3698b7e6edfcd4b645971e6788b17aae131ded33208aca38cbdd7c521eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h605a1c1d9f22a4649df1e5e79430d886c8d74a3cde6e6e8f730e5633933aa5df9218c91ba29f497a5e6763d147f751543e0d4b5c290a5e01e3bca8c747c1948b0ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cd55388f8272cf6c64fda484ad0260432c933ed768884bf7ad2cc7c4a47af61202001080f1da7b76613811efd6f22e8e185f9494431973822cdb2a5e60dba6c74bf1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h94a1d66f67729b246bc7f1ac23d75a5dd3b10d0477219460e8f64acdea6dcb380995a194a3e41cd01132d5b418e7981b6b2f8ce0c392f0429734e3fa2e56ed0c3308;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c835a2ce17b9f1415a31c3c9d033448e925810f1515e9d9c23a8f3d9333e7f07188c347ee28ea1a5fb6743a40aa30fca6301c9d316b3bc8447a7053e30046884647;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12bdfed80940e195b9a5096d0114fc7de56de33b1882f6e6045165cd5e8f07dfda9e9dafe0772705ad53d225de4f2839716d4ccceeffbde30f72449cb5841fe1ac30d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h160732a24c16178e942bd35e4946c304dbed4633aa6d6db6f45a22a956c8d13db0fa279ed62b043f6f25300f904afbec9425cd89ecd58b9259489edcd4592e831ee1f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a3d1a3b9fdd65cedf4ddba7cc5422c69f9127282160b07f273fc6b9d31ee47332a64c109702d3be3d1d006ce849c00c74755c66ce94abb451dcbd21a0497968694b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1831c6a1fc970f8f48486c0efc5f46ed9fc09b752525597882cd2200ef78373c5dbdb685a9032889cafc0248664c47560465f90e01e91a1c2e656d1c1082fca1ea4f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e28bcd8052a04e0dd398635ed3624598bf9b83dafa027f1fd87d9f7bf05232e045be34a7aad880e1021707899c6d0575d0194b90b5817ded8c88375e1183a5f643aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h883e544c3f5b473718531dd211c694525fa33cf6756b446659dbb189d3e6421a5326f5000737f9accb0272d8ed9a39c4379b25cceb2b049f3e7fc0b7bd59cacf93e8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h890f84a87e11a5781f1029915da508ee7adcaa707145e1274290d3b39c5d2c7047123ef2c58c23ac4475fb2736e791b21d64e968da7a248c942489bb3bad4df30d14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80befed3823cbad924eea191f940a3396b0c245171884b1291cbefeb8ec427c6c90449885b94d2688bd694ecfd2669b59aba888073cfe7da46c7044e8a37bb018d24;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3e499d4136a05bc3c0702ce88c0e2a8725744eafd08079ba093f15dc435237f7f6158eed45c2a9524a44bd86a542b9026323d06f2b7f7eee37e0faa2baf3943cf4f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h55a76b97be90589be976eda1c5d3fe782c4c67c9c0d30dd4c92e078cb13b08421b14f5e4f552ba3b1a5cf2409ac9c1e108cd856c3a61d625ea192c812eb15e5dbe50;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d49296c22293598f50af71cf1ad75b0f19cc39fce69a8c265f372653b9c8c60f13dfb7944488138899c5d7c9826243ef9f69ecf4dc926d0ae9a4eea0a67bc214504d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f57bb31746931d606e3ef921bfb418cd61de0302704b77375a18989f1ec99efedd7c1036a54830a903161ff9361af284c8731347680ceeee0b3557a8224ead80a68;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfdfed8bb664d6be5f66b4b06d5d1e962aa93fd2ff1fb45e7e927bb1e1421eb50cb5e182d7d146627018ca1122a3543a871320ccca375f81992f7907f4bce597067a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198e23b65bd0c31479ddef800943f3c3efab68085501ca475bc38033de6e05bacd790d9e1fb3e9d74299a0a6881de8b45cd1b8a44148fb023f4666b50a7b290a804fa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12802771c578ebe573f91d172036254d45537d45701d485c23fb8c97b37008da4b931c73a9320f50e221ede1a41f0c3caa68950b126c8d8b05099198cf210b9861f51;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17a5e193dda52e4cf66e9fd2faf218b6eaeb1003858669bb3b3cc0655ccbce58626ef377a68965515749024b027c5052ea3abcf4b4277a19a09707d01abd84349a98e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h56f683d5be52c05074d0dded8351f0208fcffe389560512f2004cda06ec6391a039367f642249c7a7f3748c3b182692e89480e413a03dc46652e823f37cb46f94505;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13ae42a93b485824b5f3bfb30193916e7a7e13771f041b7cda849d47ad3d2f06098cd3589b3f6772f29167031134325f0c7cc5a8447f4c7e9f887f19f8d912ab18f47;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f7e5cd352fe40830f704c67341795c641703bcf93f9496fa2e935e8a3bf8886ae09c5e50659dad67a26291ef40a1188e7367c26223877779595a2ac26354a0e4d718;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b26658a1cd7a1444f67ba6d3f277455eac2b9448844d0142b161ad48e2e3666c89db1821e570de409fa44db780dc841f30a628b0a1d5a1624b4fed6fa8463690224;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1613de17e670d2882dda5144a6751cad0fcb0dee817a462958115b8053bc657725060810d0208464a3e92ee52d1241bd6a8a8a8de7fe5d55bcabd9ca618e7e3d492f3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1836cb106311b84dfb24ec689772435479ef65c2ba8f17581200a759755c28d7f9d4f87fc12ad98a819b0d328c82d22fa5b3955b6a1dae38263a2b3d2ddb8e31c0837;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18a084e20dba22f08ec32e1476ffe1b8010d2fc9190a2c12174bac3d4f4cebe47312e9d9e2a682bb00548f447d41971d58ceefd602968285043669bdb3041028ec061;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he72f3aa7490811e34f25a8b037674ce2a775c315c133e89950df722ab7c529b82601da621eea03fab0f34da6ab9cfe93c78790273b09c499460f5ac925ffe79726ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177a051b3d3f6e7ce83f6a10f08fee8cf9ae3d959025aed74802cc72c5dcdd5089ab24967329d0b2e9f4abfe2e3636980143db4d381c9c364578752f81275307000e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h46e3ad8f37639991b8311396b85e47d2fecbf8bb90d9f7ff2350b0590871b141d1ec9265cf5e2101411193a1cb6c0b1601629c4c4c89cf86d12b07783f51ab2190bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h55f8c50b3bd5ecc5f36aeb766d53128a6e75eee671167fe5109d6892abb777e6a7f4bfc7f964b2c22cdb06eb5687e538a7b45d455e16ef70c506770ff33cee89cc01;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19105031d6a6397052cebabace4aa18528f795f4a88ea82dcae94b5fe39b881b249b4d92ec5d1f4cfa4e8207ad774f6e9f2aae05689fba38915918892af21052c03bc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81790f01562be703f8915b3455bf68eb35a881dd1f042956ab31a3d10f25da9991c992bd0cdc7a97d82052bbdf7c97973d61814b34bcc37d8495a72bf4195e714be6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8890ba8b127b18ca000f8f4993ac537eff53b7463df550ce51c3683506e4cf916f2acdd878ff6e0c78207b6896fbcc720cbdd5dba44239df6515a044f6fa483e65db;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4d99091b3207282b2e718436137b6d290f2c58d721591d3a217948c48d60e38a23dfa570c7da1b7dec3375a67e63a60880c78bade52e825bbe2c5709c836e83f6603;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6130fade38f5e709b809839bbe8a8183bef54396c0ac4ece1465ae7849c8041873403d0f70bfa54765387de818d52df2f5a1f3b114c3521384dc9d914c53fdbf3a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e30ab853afd1eae8d545f8c030cd0ab391be5cd479a2a6a6472cbeddedf26b4fa1cf3736304ec25f91723bce197034ccf1475a1610407ba6de4d77c41683111f24a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163fb90ff1f38e06e28bb11766665b1a9222d5e73d518503ae7e418bb9e09f05cd9978358df290a5889f982223696574224936ff7f02139bec64a852de004f286a468;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d8a1a1250113e392c7e4ebddbcde058f04bd1ef9a1f1050e022886c65a87c5d91d9ae3c82279c90aa9ace9a38181a70b38963775c2131fe4b971ae1664a2b677854;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a794c5caf829d9eb49b4655a3b84efd5a1d23cb087db27fcab084f1f73b057e276b91810bdc38a4bb4d27c1152b875d1f75692f9b97db2983738468ef1a874d1b21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1025b772ebc687e8f14f6395cedb62acb95fe214d7143e42d09a88bbac8f38b0763216ca1c422e86d2bcd76a543a22fa814bb4a22a651ea613648e91268db76d204d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c05a746f3c603bbfef17b643a928dd62d95898ae7758af9e9c314e20065eba8cb3ed0b98d35df72017423f8a326a00854a8ff076501535dcd10afe0d5e7850c14e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1828895c9663ef6f343f45ec2cd794128a19aeccd47019fb4d05deeb97f2820ea9434c7f38a51ce282bb72a92d4fd6231eab40adbd330d14a67d831036bc9453da432;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a532156d850c3a8af4a61d9cfaccbe11a1f8848fd62eaa66590d2e17ca876074afd7d8a08335654da932149e47947202be301108e917170a45e919db9f097e5ab29;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64e830518d56d6ae62e9104d9709c85a1a71f35a2993ea6fbc3e45e9a23df67cbdca660a12db69909c7fcdbf3d03cb0a9f2fb77bca815a8396b6232843f40cd89065;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h797875f477e9d4cee7fe4deab44c15a374a848cd6bf8cbf14370832d905e78492c5dedbf7df4471f4618d963dc52efd910ce7d672d9a316470f284e8149c69a32cb8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf751168b5cd8757d85012ccc9d9a7a6997ac61e47f40d4dbf56776027753a597ef907659273799cb1487330a53d1e5172f9eb08eb70ef1a7e3b2543bc2b01ac7edb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e956c1fd84c0d2e6e9f995da87aab0fa3777bf54f8c634fcce43d0e9c08949f96102024e80160a372437b16f87611b9b366904b5a5ee394c911ae58a103cd927771;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9bbb7212947f97e2229c101c5575457b3011dcac2b400ddcc2dcd7c4df4b611e2fbaae73bd9c623350054aa347bce8b514f7eb0b55794ef729e405555ff09c041b56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd0fd683abc15c9c0ac2456956df95f750e78e3b3761367b54ee15836ec744aaa17a569e1eb1283cbd13ec5c6046cc9d60881d63d7e9a55a3e481c1a6d34239c81198;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b91fa99912b8c8a0921789ff6f4ca10fa1695f0e50a3aebaa17cc5e8e42280c4f8191480212df20b0ec251266e65b62a2c8b0dd96a355f63a1d09649578c59d4683d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h475ab8c7e661329d622f7ec493503633f2abdfb6bb64674803e21797c51386d61cbf502e5c94ceb7237d571508bee9cc67ca5bfd535c26efe59f075a8148cb88c5a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a146fc825178eb8a9755ec06637d7c47456a52eefe75aa86eb0b04292aaa27c09cae1314acdf0796a998515eb122e9136e78707f278b2864dbecf93201006ad17494;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae9a3e7111f2b037d1aba9e7a3847be1a214d581885dd2e720dec7c44fe934d3bd50e1ce33f35d7ea237b46fd9f6ee2eca3da41eaaac4d22337c778bb2abc6ceb3be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hffc1ab61435a256c67124698378d2a1538d93853710c54fd1bf27818692ddab25972008c3b867c30fdf5d1fb0f3791828754639c0f0d4a26f429af83a2d425a76501;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbadc27af072cbe0cf3f3216d0764f5ca3003bf058e13383f959923b276e68d70019777842f5231f49a34d8fa964dceda4271c61a2ab115e1788b0c63a420911e9a26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ffb9f5497312152ec0f5f211eca4a8ccf4f44f0b99cdfd4497b95a18f546f8ef271ee2a1196ff5e82420e35576dc24ca6a6f5ecb0fd5dcbd684e725430be423a8d3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d850547934930495cba6595a55d85ab94881990ba14d96d0a531090d026141f213f4807e134f509ab2a1fcc3e51e4ec2f44eb51ad58cf4a0fca65e2d66c70cd7661;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca271d8c7933a7976e486fb1b53a0f50186cc5ea994fd0da3e059f3a3076b67328e8d0438dd6a320372561ca770edc1f2919c4511c89d75f6905f3e4782208f4df64;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf33aa4d48b5b704b41bf04bedf2c4fb1643c6e5a725d35db1af752497f3b7550c9c106e9a8dc8d14502552a0cd56225bbc4170f595cf26a93eb18540f4ff92c6b33f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35620ab3f76fcd9e25b08b35417620767d834f407f80f49df794a241b32a9af2f662a0aa7b9aab08366912e975fed5f4cbb472f0e14578b24be902fa208989a535cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h196ed6d04d662aaf9882475f739c0faf8d724b630bc688f218385592ea003b50787d4cf555d7afa02313f487b20b4116113cb117f87059edd1f3fac6cac5d9961aa25;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h421d5cb3016f4f0103a9c1cec3ea247f172859bcdec721bc755614e3da51670b7124725ec6bbfa44edfdddc45a6332df36bfc22b3c42daeb91416e2cafc244d6ef48;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d8e26ce05a577fa97ef798119d79dc21fef10ca49877bae941a34eb8ac4cfaf2b77fa27155fb2f57fe75efb272746b469810185c3ad351aa1d6f683eb2d1077da1f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b39e01de8823f7f98def162fe6e21ff74bd9637dea13bfe19be63893ca1e3b463a0f4d6702aa202c991e510b1abbfb3b6b4344076e793af8bbad77b042f990bae80d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4bbd9723bc253db6c26c9c7f7d1d904d37ac13e73cc0aab71b0358edf8759c55148a53fbe1fbba4bc018ce4db66afd9e2a16a16cac752e3ad99c080eb24e6c4991e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1074bb86886451a0703045ad9c06eec41ee0d9a50ec324d749528c8216d59a049d25cbfd6d349f4fac6a48d398d860e8aa3e0d977db3e973f3ded9fb27b26b543d940;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h36390c0430b1cd0c0b6c950ef5fd648fa59f75ecd269504a1d3c6ae276b1a451d32462d02378a8daf984349a5f0b44de995243d8594d1ad35940e853ec913fef5867;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e588d33b677cc7ebd6f1d88c825577baffbc2b1ed1374bb2599d3cd28b3f86abbba8b734bbcede9e68617af2cc0374877a464d126740700578c66512526bed305d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16dd7968f3d8714afbec9ded170340c8ab818c92d62699a0038f7c2cd3e3ce4df162f92e7dee0d0c0b55f7d486b6067a3b95e894948574c2d26104f8f672112aaa77f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a2927e1da03a11b14cbf126b1608201b71e14b2872d63d60ce16a246261b792670b8f34b00ce06531e5c279ac256cf9caa647e1edbd5ce385b3685d7424ff277a94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd9d6afb357b720eadf5c00d2a93108ccc94b907b090cf2e7ea6e26f0965bea550a8cbcdaf44809dfd475ae3484dc47e2ed4ff53bc673c9e0f3a1e3cf4d7235d0f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1865fe058091f2457fd01862690ce40804d295902ba85be8934f0df5fc55bf51707ad42ea3b9685d60c315c4ef45feef650c48876e24f6490f474fe157bbf2bf0c7aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf200f2c6838a06b78538b5ce61f7550478b68469cf0925a981830d87eedd0905556b38ec66668053f7eb2f9a054474e0f338f9c9bb668ca031a1828625798cc3d8d1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139deb45e9d6fbbd45694baf346fe3dd4f852a3d60f80349abe97074d7fd3ea90279d8e13aad3ae93563f15fbe8cb563bd52438378900ea37967d307de74f9718bf42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae12e84579da5160482aafd25951b80b894b32efd90e0628363c1e047c5527e78688a6c6ecc5b637eba29ebda98edc4a77365a51905b0bf8b997f8fa1428764ad3e9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d0b99113a1e8375cc7d1ed8dda0fb1efcc15a3c2690eef27a73559d5dd431f081a578d0262d2ae8d108756524a59935183463dc9b6e556f81ece8b36eeae1549fcf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14aa4ca49f5c8542ed293f124bee0c3839dd89c92e5c50dacfa237eea3655b582bf0a92f16f68a94e26370dd74521a7f3148cf9ea5ac6e0c7239af3d59349407bb6c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d0d600d16558c0c2cda467d6bd1d34051fd54b93ae0dad5c997a01a8be333c787b3e1ce22e4e3b39fc734dfa4b354bb7cc254c8e9731fcaecce229edccca9ce4889;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce36ea3a5e6c442361014c84b07263fd933a3e49c860f2b3ccec5a786ff29f4d61b5d4fa3c85c8111c15bb55876db7e26e53420926822ce54d4ee0692dc7d74d583f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h172941ce2f2311929327d5c389408a7cd760ac363140cdbadaa2a51d6f9e9bbf852cd1cce590fbc2d1f084fa8f6a83084a2906eca9e476ed9c9b70fc379e4d04472d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9185578c0e9ce5f082a4cfe7152a7594d496e36b5467ecc0021a33ca5078d47422ba47a378f9ef94520f21a66e5147372f879570903554162b644d208ea81966a86;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a32b3bcfc03720d2f009516a129fe25e3d147c130ba397ab14720db35fd5c810c0c19e2093afceaf4149f98bece752bbbe56abed825624687e9260f8c90b3b9f065;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59a6bc36676e9cc59a8682c6046f6d64f6b86d68fc0f8515bb7c761e03949f148e536014e0191685f6a24522aa2961065060bae0caa1c4bf62ae7db25adbe06e4df6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71f62eec95e1ff25a07c58f5eab103c9c30bd05df1a5beb16619d21b0c7169ccea818c86bf9f393dc86224cce8b95c68095d8a6ef4695d09700247b71226783916d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h188f45bdd2f3a2b8b17bc233850ad492222bc53d7960cfc2c3f9f7ab3d1ce7a6e0384abc3796df181cc4a60da426b64346bd5412178f825089c87bb169b4311b7f95c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3f9d59570c2286a1e34d49f6ca8e402364862fa333266461f51581e27541673141f3da3aa10c741f8dbd7710e8891b53ef59d3d8cae9cdb68c2d9063b9344651aef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e2c99b7946dbc760571097cac24c04d5041af41de2ee91cf5cf664ae46056670b4d14d34d41897757ee0c62517f0440ca91d1a45f1ab052673570e01e5d623ca297f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he752ac4b2f6ec3e2d43163c1e4ffc22cfe173fd43ccd634009124a8540c448441367a2fb20d7a7e6d0d3f02622c3adcc9ab58c2dcf58398ba6bd35da9f866cd94ef4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc4dd0b25ee8aeaa0e43d474255fbf02310a7635fb2875a8bb490e0c448ee9cce8e41f92ddfa91a2aadf9e2b01788a1071ebcb2e7b5991ec5b8ed7b5288da7bcb08e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc719e74a53bee4c33e51ff508007ddb42e8bfa5a7a38776248b35bdc24193dda474b0aa4309ffb22a84efe80f8763008fc7bef10c70c647e80521ba29524e8aa183;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b96bb98aff0c071330165126a4d3f598f62a750017b4f58273f48da9810b778cd3cd1b41b4ab1eaf97179f9d5ecc6b1b4b7afb20771e99305f228420aa72410c4ce2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34dacab2e8b58d97a4e7eee2a960f0d88824762f2e58173f85c2bc63ab7850503bd1310838852ca8ffa18c7063ee01f52eda82109e250f9ec734d1f95cfcc4855a80;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10550939ab6c9790edf052c46bcbb8366a778498f1e7ad16145ac6ff894737b3d6382a8c9c2bb81475d0af44058e71a239c5704a6549d76e22b6ac963e85fa0bab549;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3d707572e657bde67b4ba520a3359c7a35624adea2055d86e74601ca0d9a009510546129f59cdb47263b52a8c12a182c9a9fe4d566d626953b97aebfcf77c5fe08b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15285aef2bb61eb1c24ef3372c1a0cd84a5dc2f4007feb70ca7a273317d43238f8e016d09ed176d1ced5168b1575d590efc77499b808a529a077fe6f54caa7716339b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65e38e72e551bdbe16355a04febf12c19e11c6aeb94090ba721b44ff24e5dd6890fff3acdc85157f82a7a5ac97bac15c99e9bfdd26dd1b402e348bfda7fedebd5897;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15843921f140bdf38b67fbbf1e0ff486e20b9da25155c8de040fe6ae8216dfc3647dd3c8719028f8d150e43837b147012c6792d00fc5574ee7d064453d7d731c36323;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a4ec2b03a9db727c8ff824cdd14a2d6643447fcb66694fd3e36cd7252454c989af82e5893349f78d8dddc10982d8d8f343ed34f99b49f6740d5c3cebb8001695d72;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f98e2de409c54bc72eeb03ece19e2cf5fcdb9c6c5eb18f1122cdd928dce021419b244a503d9db1bffc9b2e3a3b0f01f1d10ce46c781e44cf447b7f2089c49bfe78a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e3d6f180d73467aa92a3bbf4d292c1d12672bb6d483a11508dfe5a3b8d22e8e9a1875c15fd3e48198f5c5d1ab7dd7415312a5382e34274a693f796f5a9145b968e33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90e6fa70df44113be585288118b5e26ff894ed00df32ece34b864eff2215d150222c8e9c1209d62b9383a95aea14014e6bf441c472068f15f00eb7388882569572a2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd9f301db75c54b0edf993df044481c2230daeaf76c085e239f10f5f4aa1c797bc7e288b2339559dbecf51e9349722eaf500d12492ed2baa371ca3aa5e4d8ae88665;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19061ecb0153959f115fa0b5a35ddea5081e30b0391e0d6a2312fc965c9ef6228e1b8f16fda9eb6e06c31bff3a933eb994ac180b45005a206236f13f7b95547f7924b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a218ade44dbbc88de021416168324c23f6f6ee9aff4d0fe6169a9d7806339ac8dfd8e038dc23fead34c23ca0b513c2b365bc26b6c8c510af48d99abe4573aa9f83f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e36551e8f03208f04c09064d871bae164368248388cfaeca04cc9eee917bcb1fb170be388b9eae38fb23a71fd0d041039721d60bb0dd2241100f74ae7bf18438c3c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68a946f86f01244d2216c2a9c2609119e288a09784741f7527e648e38e9620ee1f04e2e8894ce5f172e01333e22298620435456f5c50f672687879fdfac2ed2d53bd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1acdb118fb817f1ab05de8449abe03708e8258d107d24baeff233cb3d0df9769a29a2d3013a1727aac7a2ace23b56897319c17c8611fb8c83c34fb704d2e90e5c2bda;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3d0f9d0665a07becc23a7ba9b11402b53cf7c5f8d3591c24762f54b04366b8a67046d12db805b601eaeb46374f2df39f9f6f3691c54bcf21f4ebdea23fa4f8bf9ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2056cc8fea4809f97d60208f7ab2b7fd3244afacfabf9ccebe504180efa315de0e3fa9c4a1dcc73b546c107cebf004f17eaf36a6cb77d95ca8b38b45203b29284164;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf1d588e9c918b7abd7ea4e29f62c1362c9d5cf55b19cbdc2f5df2c0d5385274c571a350d9bc260521cdab1b5b290e0b0e2d596cc1faa9987291877358b2333891f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145e025a5144a7292baa39cd6dc05486b5b00e6f5baff51363cfee5eb816750414e77f587009a71fc6ae714986aff6d69cb74f7b1f48f3e4457e8f591e522c6b07949;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3eab8704a1b0d33f7be325a4726515af4b6da3f39fbdaccc7dbbc9a7de049769817ecdf2c70afc8a0c2382f2583862cb9a3a5cd4cb435948d2b0b517052c7a135f66;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb779df033edd1597a684abc3bb7c62c13f30e4cf569e220a51086cb470059e8ee00e9003fc91c1c93967b97d3ba598325a324dea49f4038c2d8c7e0908f8b7c8c14;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1513135d4b281aefc3166110ec6a5ffc213144f46c8012f2ebde5e461d39821790c37eb9231fc0a1bcbdbb33f9739a1df45d4236898c3f3a0cfe4e38ed9ab9792b7f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc107ca0346ff773a44c766c89e667a8169650e4119b91fed78b89bac84893196d6467bef488c393792f9c80603247ed6ac3fc17073ff9d354cdedef48dd5fbffb5f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f275c39966b969ea0d8e06dc82302e75edc51a0f0e8794ceee97a50470d685b76b4d6c054b92653a918fa041b5a3464c85a31268a2dc58ca2d1c146e15771c63a105;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c1a9c088aa579e6249ca5e5e696e8ffe022f620470013593ba6eb97682e43ec22e85dd02f130548696d9d619f68ceb509450f42f4b74912be0f65af89b68001940;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7d29dbfe361f1e66ae55c5593cb8949576c780c76d0b64813631034b73da6369423d37d1a2aafcb760014627576bd11a65c740444f2a954c7ff28a52c462e500e7f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h887e6d1850e5848871ef5f778c0c534dd222a121a3221faff67ec6f57c131fef16732be58eae4bc9ee9368b87b8142c3f01d49a8b550eefeb83b097299cc68b73bfd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a1805452d2752f0d9a6f79a0ab72829ede67a377834c89871b24b9d85d25ebf4757bac8dc056227a9d7efc2a22c61e25eff5845a0f27f2ee497ac56c9da8c93abe8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h943fd1a7b73b3b1012de15d424dec4dad45835090975eb62bb6043f358b571714330c2edf96a649b14fb367220dcb5560703b5bb124c77eb83cecd3fec8d0a89da29;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15dbc65ef3d967f114d34d9bb636112b336f0e3c8ec262141a166ce8e120cfd211f4731132508bd22b6a2a7fc94ffe110831368dc4f6b2ab2ca27c8fa772aa9881495;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17a3b1161bd86412e5549d4e7443b7fcd144fc75cd242d36d48233d443b88aa81b070dd51db27ea476e3078780782e843d6bfa6da37a27e92b3df866a426b6c0dac5e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13440ae2878fb1c915406f0c7df712a2d0e4f981154e8f594048dd63caf5b1f4f3ea101a99008e8c580d5579b5e6158f1e65d58d2552cfdf540178853e79c1b64463d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h147478df2df0ad3e4b7d9109599147e838cc04775c50acad23ebcd5240dc3939f9e6f55c9bd02ad105c9f8aa6e007175b243e858edbad8751dc32af4a48dc530620d2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67f82a19414ce4631641e75fc2a31c015de9d6843d308708b38f1fae560724455238b916d3575ac4b47db411fba05d166fd872b71e127afbdadcb8701d202b01197b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h84a90e86459e1c71b73ea1c60174874fb3a629fe1f790e0696b26816b1525d40736b12cc667930191790366d1fb34b47df9f6bf52d8f42ff724a9bc8cd884bd57b54;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f64bb83de0d6b47333272554a33582f0dd97b5645241732a3a404a2097fed2d6d80722a7c2d5444d2aa7962a00ee56a7478bc783d48f3af04d6e65ba3989a584bc4d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd69081dc35063d93b31a5fa0fb91a20e99837500483bd36caf6b3b3d252fb2ccd8fc8971325a7b68fab11d977224882f49a8c2c7c228dcd868661e4beb79ec2779ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14843791cdcfab833e5bac160646f8258905a73ca8516904d417f1452fd51f1b5379c22b75ac4ece66c6967ea7cfd6b05f3fca9cc5484c6472524a1090d6a0512cadc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7835c4c89e55b97aa1944f1010eddfaf046a276c86bd6c2b553c1da34532b23257c6debae067395722d50fd05e2af7c38902ffc0ff67d74edadd32025e138127e06;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h147d457c3ef5dc71948ecd09a6a0d8f422ab4b42f8d10cfd5c339f5af6e9461c2de49b814e4c435954abc5e1140f5747cd3c06de531100b8f0e5a946204e79cbe4ea0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb2c731d1b2a2170d7fbbe4cf793da94b741b05eaba5aac4e33d1c653533bb72f76e7b4b9338f3e4537e16f9c5ff98ac947d89d8287562757ddeea8e5775f687131;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h180820707db58b303c81c5cb4f2b11d7d326cf902ef99dada3fcc46f4c84310086affcab78454ca132c039aca8d160ab485f4b4a4f99c8e3e3e351ae89bff3b083a41;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha4d488e34f5d91faa48868af84dd854879986b96124b78890774d4f89e8298cb42dd17a05dde137d3b81b96e7e749b233adc1503db72a32fec4ba5a2aa800b91987a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc8d37b458cc08ebaeb3f44188471cc13f428e22574cd8a2a959c7959f2ca2b01d84bb02db6d4a1db5cefc7dfec2277cf608fb369bd13f3abd9bb63ebb25152b21ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6525ef378ad1b9cff41b0d48b8bcf9299fadf50bebc605cf2699f358008dfc36a2b55b204231d06fe07360e79bb47e24b1ac5ab058ee9e185c82b6707b1a90410d8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1986dbd0c5166582f4734980efd19d3fcaf2adb48ccefec2505ed039d564c1db7d19863865e5f385387170cec97ccedd6e71185a1d24281591ccca1d427c7d8a056d3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f9fc5bd1915a09b188fbd0dbafd2c259940698d3a1f090377b8b4e12d09e2c13d3bd7d9fb36dc7d96fdeb88a0fb5b3c9518ed3d4fa097ca30d31913946006d5fc43;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h165071874be8187b496406f13c93f2cebe8e75c7aead535dd98b0c43644a5593bc6435363882848e77d5ce985a633fc0e1c7f3119aaa46bb6e21b1775350e7a27ed46;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff862ea4fd45fed8b68d6028b06c98ed872945d7cfae4065c05e37934c782d67c92780fd3026020bca7fe1eaf4749714e96731f368abef4f2ce5a0c1dc866f78f142;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8e280271933d92f7c6673af232db53a357b262dfe4bb1bcb2529bb98c1680b2d2712e439380e80b97b17f8f6b130bc243e61436be8151448e69fcebd951b0524745;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfcd267339b2881211d9a26bdf6d04b7caaa0f3b3c9933c0cb0da50dd863634d4935b88c74c42203050d45d568c5998a9ef94b51ac552d5aa2596c878653585e2ba4c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bd7f36d5b6eaea9c6b4ca1ac4fc6ca760ab6095756f6acda503d7db7d34beaef21a105324340f4204de930fb48bf5bb3f7a28f27dd07817523a499035a6d0263794;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1344e1bf773796d1d4d5b890aa2bfd49f79a7a9832bd35c6c7b5aa660a67378d0871c4e560b9a17d9ff7be78fa0e704e684d2487f5c6ff66b0bab0a59db727d94b015;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f9764bf6e798a6f793d830b33e62a83f7f19a7534b6e30d9d2eb7b455f7c064cb3c916d91ea1f6b3fdf13e903a93fa6d8368943916b3d56ea2c4a63db06cfa94860;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h908d0ecb16f951ace26f9e050940dafc023aca64cb62517776270290d3e4322a0ecb0444c9c40ae7bb66a60477a705d82dea816551994d65d5f59ac20e78253a722f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he66b8220a8b4e5004b69813b3d413f701fb58f8e5c256b0938a5d6e5a50ddb609863379b7bf5e5192917a4ca5285a41ab833c3eef2c5c36cc98763ca9d1e0ff3da06;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c1efda094e76d820942ee0a1a232c835155e1bd54a7bbb23a4f9ce298794780030e762e49b6f56223beabb6aa9f87c2b569a6c32a182a0a569b5a6deee7319579e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49c620af4a97345fbd586951b98e080f3f23b23542d37758da142df8770dcf34397df338924de65af71495f6c8688f9ee2d6eb4700e8ee7f7f15de610b88da24a760;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15806bc3c1faabf48d02739e56b21395dbcc411d6acbced7e90a3d2692f6841c9d4166b6d3ac2941b4ffd94d7e678bbcf41521147a358bed6bc14324f5716f3a92c71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bde3fd82e049f5c573b509546123f0834b174a9e5b736fac2cee53fd687475ddabad87f50ec282aed4546567ab5a6e14a7677f37bdeeb847e1b07a18f26f5d75e142;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ccf16a2cbb5dddaffc8baec20d7164d7bcbbbc124adeb846743398e351e3539ef3b78c504f410e2138e1b092cdecacf4da937cbf80ca43cee26f9936393a1d9e068;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c25b419a00591ca10e328c4d5ed5931432eb7939b0d26da485a79ef53fea9fefef4640af34d92d0a98c1f5ced910f73c807b7d1671bab62b951f339c90c68edbf03;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h191550f7d04fe4f1bf45feb25906f30f31e9345fb6b7f7f8815f7de83ef25c544b5f68b4a55c5afaa3bbc82135ac5635701fc2f501047b90e7e7c38ecce6c30953ff1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f928811745cd8022b3ed4872281910a5c5c438a666443ab834a0d31e2d659118d5738e475a9573dc1a25adeac57f46e537b7ba7584ccfd1b48f6acf73bba987eef7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ac3eb368874761fae1e14c6703c9c4ad655d07ae64aeb457fca2808cc7259f7b2f36274006c8896850564cc3c546086040ab40238bec8fbd1df307e61e4f3f16f49;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6a33c2ba3f7775267a9a9618674fd83b9ce79f65b2a66e1ad33e703b575a185e8ed378da151b4d2a9271f13dd7d5c0cb71c355cfd7141c519917e78ee61448114bbd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2087f84c17c905d43ed891aaa0f7cb4be5addffe26e05dc6024dfc73cbfd4ca1677c8a0f404f46623f598b1352e577ac08b9bd33353ff6991925890b420422a4c6f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd25528fe53549eb3bb24abd2f3f056d039f59517465e9a87f3793b9575969bf33b6b3ed1a40562f6382ffe1b687c3361986ddea0212d191004f4d33ae37f282e0295;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d1162b6f64a8278b44db83d4a4b11b3d8c65993af3624c27a3bd8398e5bcabe55f0aae5212d82fa1ee16ef1c3816414ca3970ffa992109d5173a5de7636e64942e79;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16608344678bd01aa90fd803829991ecfc7dece259c9269d1333b12a282d229c70c79c0c97da759f666ef88fa6a3502f3660f0c50712ca4ec798540067d14ea448a94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hedd1c720590ff0cc8452b4ce1b38903fffacc32bde2a06325bf1b148f18269301462054a69996b4afba2e0094c462421bad55c62ee16b8056fecf9d449c75a623ef8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc80e37374f54b9c39fb8f1fa53e66fe82d39b3e83942f231f4fa3afd84fbdbe290a74af452ea1da3fc47b6ee4b231e3fa7ce19844b673cb6f8bf4dc7863d86fb833c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8ffdf5f579151cadd9da773de482c0f37c1fb542692edaafa6e1345b6e9c1464808128dd93f1e5c8227f413c2391cca3cf26357c3ea98441c0aa1d013d465baef41;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1184a27a4f9ab870dbd40785aea316bfe6278af44e5ad908bedd0239d114278ca2e3fb886ace824f4d6c4c2951002b99d4ff74b6dbe771c8c76bad6253c40c7851fb3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5841f6d4982292840d48ff2b6a55d7a9a7ef6f7cfcf3ea0117c034a910d4bdc49817e7ea69c71847eeb2484226ed916b999689ba9b17a651f3a103390f593f3b685b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ed70bb73724b270e0b9ecdb2bd473d5c2fd6cbc5dca4d2fbb8db5474deb783a7143f850186a7a5ce780a2f144ff7e063e1e21c3ad5802c83d9f8ee57ed231abe65e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7b96a5807a9191ee99b4342570931ff9dd37b48acd8f50dc8e5b3f8c29135f399dfe048ba4028ec8a4a5761c3a3e02d2bc20becaa98a622f65160a3d8021b3dbac2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a8510e9007b484518995d0ef8bed1564a25b514312ade2b6634a32d31bcac3c0d044f8a9966870a9692ea7686dcfd7f486282f64a834416fd2c8bc2308ac7f07d5d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde89beac667ef0795a35eee3d827c2e03d5e0aaa370e25b1cd36b00f8c1ab2d384beaa28f855ce781827df5a9271b411d3ada59eb57fdca8cd7bd5f6de8f07e63ff3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h56973248bc3c250dfc366305e7ef744044bea9e131ff7473f86138abbff9c12fbbafe7018b8e42e735b361d3dd9edb27e4d2a1a9ba73aa1cd6664e92c719bc0d3787;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e70000cd7f67f63e211ad23719d4e3755c59e04ac67aae571434a249fed548612302bc2151ecc53832a103398472caf7c4253c9ef77b47275dea09647cbd7e6152e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1935067fe8e247eb47286db0be308efeb48b3f34d1f61c8ea5caa9e236d2913f2aef140c1352942c5b83563007493ad89c12676eb85e0fe13a9324eaf3527463c908a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e900be153dfcef415f94a8de44baf4f872fb11979a614bbdc279cb52444fa1ec8eb5d178589a56b315f2d00ee762515cdc7662d2b7ef4dae31db55cb80f66420106;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d07dd800127d256b88c151630bc9dff64ab83e78e3ae445d07799b3f697a452dcc7516057e40a92f8d514d25d4190d4f5c1581fe3c284764ff9da509909beb4eaea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a20bd13a35ad3ba74cd605b59535dc8bc409849365dce7fdc51dc21b9f3e0c89e76c6aa566f6e85ac182043b0f21b813371ebd641009ceaa439c00b3c75c3ce6f5f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da0167419470aca179e6f91834707eccc60d6f2f99110f02b3fc7957d7266ad99f1821b3bff9d8f329ff3be29028b84e50f3d131c6f75406a6b485dd3e754aeab5b5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd025d2388ede85042239c1ac600b39e739cdd9d03fcac550c2ae47a2a037ad7387f027eb334c38441d06534f6a2ea2b070250ec244336a3390d425ebea563a80beb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h169ac79b3b05552b889108a9f57cde6864ca9f5ea1aeb25f896c8bf64ede9aa73bb1dddfd778066c9004ce52b50d45ed7d65d866a8a39dec1f26f23b4649f0e5e43fc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde78426686d6b335ed7c66ea5438e416c2499db5af30be761ea2b6ab8e90192bf3c49d965d762e2b516037103df35b9d22165dbaca82ba21c8da551be85adec5fd10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe728fae9f35cc485943c9303551316348d6a6bdcba08cd3fd229469ee96e80be13f454ba39cc5fa690de877243beecc0b1c1cbf60bf5dc9fd349e37347820c0e678;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd2997ba0912fbadce5dcef2450b366ed56e757bbfce83666453255427408142516f6aa61634d45d824b416cd5091cd08aabe5db0e0af08cb65f61f998e337d5e8790;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf195f5d8e0a10a8f0ea2fc75e979271a8bf13a70e68341b748800a6f1ce426eefff1b4d1b1af719db7692943671a5d91976c1ee15c209d11f632cb39fa5e85fce17;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc484b222e47a78ebb18b05c9ca6bf454233ba4f9e10e03a304e011b3661897cd21546a399a186421890a6c189b2032b39d9f24d607538566cf1494e77648c25524e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha630b1b1162e159a7e653701fd7018abeb06d17cbb398c3756a7acd242d5de3e6bad3fd48c88db2c4bab56584a96f7beb1a38e73a8d44906243d05ee5b5e0f64cbd3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h434d774debe6c8f5886ed876ee91fe8466778ae53fddcce64100e1797608e67c48b63a444ff7d3c9db4c0fef37eb4fff244bf2b67c071f83d99207b8c0da8797aae6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h993c2ac8004fe1fae46ce663b69445145329d77e40e8179ccfc581aad05b2bdf8102a99a612b88c828450cf1212e362a7e2631725130a87c217b73e43c43706b5845;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbed4ec44862920a2b0e8df68399dca2f71b23b367457dddba57672ab631b1852baeae281088ff281b8cf36b7f88188edac040580cd6688c0add6f62e73ca8b5136f6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c5e9f6ec4a8f038ae3d58e045d9eabc0486e5fec7a725e3216b0dcf020ba861b44416564fda217ea07702602e2971c3390439f9303faa9d44b3ef817bbc9bd93ff9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1105cee72271a3b605dd710437c68f3b9622943ce42111eafcf2963877c61efeb6d6eb912483434c6347c54fcb7a1960a95e3e3aa2ff5e4882ed8b8d5fa6c8a5253da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1339d6d77956de9d58e195334a208190ac9c4792bf16d4a6092a4f6ee731847f4acdefcc852f70d95fbfb737dbf43655ab1c9bd474263c73732c822ffb47b344ce26c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f0e3b274f172337dfeb43cda9e6f92053475845fcac7d6730a2fe72a9693a5cbc0c8fb1d7c2f988d65c5755b0a51f8cafd772f16326d1a87e3f127d024a3d8c0ea1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h124f32f402557cf9dc9223fe6822644755dfebac68d3a2d0b1ae33a31499d0e3f4d1798e7e05fa5d6c3c07ea98fcc0ababc74de88c82fa72866eb50af271bbb250b3f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12738bf38c506c0d8e1554be68d64de5eb0ce7c0b1f98cca1cd070a9da860761b4be04152f25462d6cbbc365691066b6848f8bec00d4359c80db1c0ecbdb186438147;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb2e0f89b8d293138fc2cba67e131dbe016b5c743cc3ca64d6ac53dc19a8cbe30792b0baa878c70a2367d0bf9e355cf81ec6b290ef185842c52fc9c0e4bef452067c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfb2079d77648d5c00b09323d5f249e3ce4746d671488df0a84d3dce46b3552a59df8f07e2c0132f123cbf16b077ef89c8d373a9d7ea584be983c3a723755ddbcc01;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h105c0176a4aefa41528c9687e15f6a4f5515fb68d65036818ed349809d5d9cc18a66538e3b126c92ba77e02c449d9c0f64b18f1831905c91be36268ff8b5f9fd22430;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155ea3242b0fb0e7983debf4821aeb8fd406fb5987cee72e12fb3fc5e4218936dec5d44e9d9445b373a9e6ad6f9381f9511b4b2a2c3a206bd0305386490ef656dc427;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1faf7a30c452ab2fc13170b2c3bbae496f80fc7fd6db74386185da0b74ea5789d3f6bc4e0ce8c774050f484903db17909baadf3c929d58ce75b69827cd9d0d8699054;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f9d747bacd5cf13a0c0b647cd07d437f222199833410378b296bd70be7217f25de914ff872d926a04a232664a3abc5090f8423b0555c5c3ea3f1f34fa87b36cb9f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha82a00b62f758231015ca96f94e99758ca02c3ae3b97c76b023a0c43f7b9935b03b505cb14f7d56ecce7f04d2a33c7bf0a34f67675f3e2d0e5bfc891d2bdd3fad863;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e020f6bd03dd0fda66c0a5c9cce5eb3e5c4583b960ae1a57d0322e731209194e997417e054b221bd7e84060c3a98be19a4caf6612806053ca6be01bae074d8823dfa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161511ce3e3c051580a67f659a26de003eaf8863d25639c278d7a888fa61709833a317bf34613fada417523ceb8f4b59ba21f1912121a10bfc6387065298cb50286a1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17321304a44ca250cba86a814d5b8ef97138dcf907ecdd00c61fc38420a5233bc77962d251e15d3b34b60320074c940ec3bba0f5024a83a628aa40786cf24944afce9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed69d1a21173c5548eb1fc07ec76def5e9c69dc5209677abab11789514efe4e7bd468cac3f85a0571726a870fa7e73063f3ba528ac0bb52665152aec434301ed3b21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f33bfc28883e96edd86426ec013ad59db4f91dc29d479a6c0e3d4feb47477f456e4532d469e532652b04fc306feedd00af994db5a96a58cc3dfc6450ec15a9f8162f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12e40d64449ea4fe4489cf726a53e1b95feef07b82575d961b154299666a36cbdfd50711abf87ee1bd87c906577fc8589353fcc7ebcf65e89c52a49c673d49547eb93;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6789bc0a93cf6d3c5c023b308cbb429e7f37b53cae94d34c39f56a60023a43347b12f5eb64c989288034e55346d0d4b43d44b0001a5d0333e3939ce127bc0ee003e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h737653b714359d85a7bc2ce6ba280e5e5c1709a25f3ffbff3e7c1d0f1642af176887c8ffc7db474cdba34ef20995de4a77f6db41d133c5e0ed74ba20aaabd707ed1c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1580f47064431df62739ea3658cdd1285116f78f3138e93b272be1fe42206170835aa477d410e4882d978e5445f593b745dbcf6aa55e4ac53d2c3e80dd7763356440a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a79ab1e4be0dd2f58fbea3a69f06184f2cafa00d4d01decb88e4bd15691e88e8e9db0a37d59c1fdb0916391e2e6e7e18c7564edee0e9ecc23926607051e2cb5ce65;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16250298a0c31adeafd3735a24a74bdec666874361d0664d504a937e885b818e32c71064e23715b0878cf066aefb358fe8e810d7a9507abe4e94a3e0d97997b95a13;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8097b83e92d7012e5aa4715fbd72fc1c0fbeb81deb3752a547d311e8cef7548dd7da09ba694506d4f89b6da889f9c21b51653b77e2e80738bbfc871304134a018173;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96ceff35e4a94b80ce59144f225556a6bc28bcaf78bb382f706ccb3491ff9f1dba81161d9b595a59cc496a30ced51415e6920312e1af5196816e92261cb2041082cd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf4cc253d5fcae2b4be0a9ad154d88720a152c177d3106b53f703fc2710b65dfc35faab5833dfec1db11cb408a0aed34d1a502d0a5d6aa2337a1ae43c3fc438f7f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e141a0aaa5423490ff592a4f34b5573c15ccf265827a42266976c15cefa369ce2ffe7394e45230feaced891d9675aa7862f6dc7278c78deacb99849b841b23b344e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1054529d692d4831d4e298fc37fcd2368829bdc35692f444dc65ffa062bdb345912399ac54818ee6393ccd5d3477c560aadb7565ccd88c6e0dc5dddc3ac830580aaa5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed328440132f27a9cd31b5639b59413eae3b43b13488939d5ddadeaa0a72e33507611b2cdb5d6126376d4717d6a9d4732f7392d0fc55994cf88251757b5ddae3a451;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he90a7221f2c09cb5f4168598d99f964036e6208679c7eb3158ecc5e6ea8b8bd0de4a2da6fc22eb3ed13853cc6914fde0fcfe86db7d7bc1d1392caacb72aefebbb382;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6c18b7d95053277660e423e08d007827a62f6d810e831af0176aec667791217a239c3874c86ec06d65c7cef635df77a417079061c0a392a6be8f565ef04e4405b30;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdff07dd8af967566324af9f1035e7ae46855c104d1adb04989a035b5fd64bf96f75c27062d8bb1dc0c94da9cf7f58115dd0fc86189f6ded3b8c94080ea4b122e278e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1adf14e7174197a42e8d02eb3df9df989e353a256d1db3b4afccfe635435d4e83983325e50a3e4a3d56df354ee28b439d5172fbf8b0c78a27f189570ddf992ae48e2e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17fe4956eeb422680aed0a173686f8d88567ab1afccce66fd0ab1cbf6bf457e4ee62a215513b76eee57a1a557dcc87d71dbe97df4217fcb2fca0019454153d74186a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91179a90ab3012bca936daf06e73ee1c2ca8d94c64eaf6699f270bd0d2de6d87c4a24986bbda8122e68a0003f54135d83febcc6a20b9d518ba68f3a420df703824bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19def2f1fb254945331b41a1200a294de37ef1fd2272f3f4a3bde8e262d8c366536bff24c8f13f2db5cee615400de31c70e7d8ee10d46e1ccba9482ca4db0e867a56b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b2efec8fd6a68970fc779f8057dfe465a3609da07fa264afd50da3b59d63e60a18b4ec390e2694d54199747fbc52fada6e0b6945badc8b167712beb6f9c299ff38a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef644ce16441e78af726b2a995bb932072a87803c5eed9085fc4aff5d0d6efe9a781b5fb848d2c147fca3704d072658a517699fb02f24b5c1740d250d288bc4b8f98;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108c8cb8e425fb59d70fc8f640e986247548ede0d8b825814df30ebfdef00c844d608aea67d06886f69f760f286a091279dce4895c6fd5b3cf580184d14c58ed00a66;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4f56c9e07555ef1b17d47c55abd142b9a71861fccb2e8298a3ff8781f9f6cdb13e4abf27925dfc7473c4b6a46da1290fc6d38aa9521ba4483a8c881a9bb75217ca9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67d3f3cba5aab5defcc7826226252efa55cc2423e1f4923b130d7208f39e1ae80094fccac9a027f617e38ee26753b958cb7e24e61ba393a2e8eba912df5a6c9483f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf6ab69d000f5498e1c75002f14c5ee7b4e423546ce77369e2baf3479d0d3c07627dd192120dac753c3907cfaa58b6a81889bd18efa5762b231c39dcaeb23fa555ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d2d888c4317a74e4cbf638ec61a5578b98fe2c1ed772c6552f25cb546308181412a383f7047eea68769c747f25815a4e120db070e672e563dc8cdd80f65faa2f424c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h740493c4083de662305934c60cc70189e4eb3f1c2850e87f864f9ac3effeab9f25917cdad08be0a4ea3302f94d66c03973a94efe78552fb653bb5a6bc6167ba45f00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199bc2e89350a6d7145a16d3d31366b64df69551bfafd7606583f4c1668acf3391232e044a51e78202abdcd2fd8ec422f6ba80e12d00fd8875bd82fbbdd8117111230;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa281d2792c3a42dfce55f5ebb029d026750746a58be23c859038312d1cdf48c0c7798316a617ae8521e8ccc34bde0f3df54890d60dfb2df6e237c7c57544865e9bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f767a886b69c62e7847fe6da9609a60d10ce2ab02fa7bf1bea2d9d845174aeb69ecea63d8ec85d27869ba5961b8e24aa213d20f8f5b1ab7078b84724488f56c28c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d5f3d3c0ed6f5c9a251c53a3c3e7d73f2a336563a98dd9935006d87cabb3a505e176c5e4ac1dd570e50306949ed384c72b7a52ba1a8ea04660101db327e8c883e7d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139af8e54aa7a9d8f181cfa67d0a30bc62502499a24f0a8186181d7d8c92ba371e38ec4c5c71ea647d0dd53adb6a7f04233fb07d28d09955d7421a04c3dc9583db568;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha152107f568c39e26bdd7279ba5034adf1d9776901197b56f7896f89e139e36992d461aa7654fc874079420612e034d35b1e80e4e9b50084a895c56f9ca15cc27bc9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h605c37e75cb7bf2b6e201208d755099a9142cc95b390a143fd951b933123048d2f83a10930a48d15f66e3d175f1e6de22747f43eade2161e2d2c6df892ae2e15c69;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8422dbace765080dd61bc14518e7724163f26788686720631f13f14af021829ae19cd863a091cc1cfb07c2aa869471fefef21472d5da1eaa4f60070cb7e819b66cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b156dec6f1de6c590cd9d8fd4bce70e02ddf4ec2737c532d95fb93c0ae3bdbe51004c3834cdb9a0296f7951c3de32bfceefe35b352a34d213cdd52f47391a7a7999;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde5dd924d1bfcf4c5b03b9629a98a9add5cbc745b837bbe668154897826a0cb691bed18ef9fb35f7690d5d0616db42e5197bc29d31a5cebeba9fdfa05be146db9e3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd66f3988125362d4e69556c98973f0a3d2b8b73708b26008ffd1049ebf06f74f1dedec1160b2eb47f796f38577df30b761bbb89af337c8fd386bfbbbf48ec92dc223;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61bb9ee7e2cd2b23512cb4600ae2445396d67af2ca686911154c554caf6d9f79b23589744c7320ba9630a8ce9423fe6a7c77590be5db10ec3dadd6094a1bde47f887;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83901a4c45251bc681baff21be63521e379b5aa6fc78fda09ac093112d5f03a3971848580c45d4b90f51cde3d33ee8a75650af534e73c4b8082d10da746bac776851;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b00b1ebacf0fe6c7ca96a62bf2c5a1ad5a360d8c370cdc31cfd8bf551d2bb086d0c2c8267e32800af7ae11fc39a556c16730d569d5367375dfb3a27f7c8870ac7c87;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1608ef0873bfe0af5d21fad6c98f87db14387c77cefd764c0f0e2260cb4230a898af6fa732ea95f3862da5317827e328b92b7045e4ece238a5a017038fef52ef55139;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139b6d0e6375a6bf51825cc049328d89ae937502ab96a0add82dd852fd26398865ae84c9742f183bcfb06887172f5133426e5cbbe5e40ad176b39a6e2dc73bbd4b636;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32ce5d4071b3af43ba64068509138b99206936f01ee968278928e3ff5f0f345421725ca4b92682e966231ecc290c0dd8bcbafb9f4d715e0fc3c76a9fd58c8cccc924;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5513a541a54bc1a796d11e612d05a8e2f852d4af235fa175b8bc004ce7d47b2fff420b44974a91c005137203b4ff77de7cecabe48a49bbf183ec32405bca6b9aed66;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32ff8fd13718fb15e4e61cee27876e4d8226f2e73aea03e4fe3fc4077a4fbcd8a2f59ed38ef07fe4ab9548b24ac4bde361c5e25aa284eef9e8e0fb1a5b5c5a9aade5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7239d468601edeee957826e41de0c7ce6ca9f6d1519a04f09ffcb3ed92356c39e18ad954f8bab6d8a25d59c8d9ab4a05c20fd705654a88ac74dd90321934f85bfbbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121239e0fba8b77b200f6a62a47e4d93bcd5d9b5737fb5ad819a73e7e0091064a278326ec8b75ae5a427ba3f02c13268a8ba6d53dcc6050f2834b3e5b3c7704a7585;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a02b80667843f234f6a84d5a3b54f848f731e85d3298ae4ee3b438a092e32ab5e4c778f875ed9298de0b27fde0de8b843d173e25ce1d8826148f8992fe771b9bab55;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185188bfa5d00ae177e8a62bc9d873c968f43893e71d8f895c06417bd9a8fb1b5a93dcd5f246ae8b17e88ea786759090be005db787c182262c4994005ac6b4c6623d3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h230b51c3249c21d01676e04bf54f6bcf10841790153c6484ecf0e0f0c91f8fa90630a966602b53412de29a9affdda52c83fefa8c888ac424c5460fabca60d0d7e2d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf107b8bef7f29a71e4feeaee381cc903fe8f8766b98990f800aa248edc34ca85a7f5c56021ba854418c635f15b84ae467c2e0997ef7c73c335705899ca50f7d4491;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f41b53c158a3f32789501c08e0d78bb26da2d3458c8db55a752d12d03512906ac1d9d1b679c02a241809c5641664492caa930bf7235426768512b97a9f35dcd2f2e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h356b0fc22e74b259837e7e472b8e3915a89c7ae67c98eb8f770b79ccc95d0872b78ea3f2f8374e1c229eb434e0341edac92e450f6b9b6c4c32b300e2b596ebb913e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h23daf8ccd0ca203192d7f3f822cf7664469c540157ad3f7ee8313431042e4d50b1faf646df49f469b058c7531efe85f2492ced897f7751cd095122e0a6c61c75235;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b10cdce2f363855f07f5568ec1b2969417c9b7152e71256149d0d7b4a0135007fe9a920ea2e30974c5e9ba1cfb484f77bd8f065ef9a8372e9e771f043f3f7d3f2314;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h120d03a02b0163c08e7a75001cddcb9dae9eae2817b971ee033a5849052732b386dc7e93dcd82602ef2e813a00a50677a72e9bca2ec47529328fea2c8a8441283b39b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc29a9f85ba0a83158e7d109309bfdb20e8eb88546b72848086c8bff03b2c1c48273e7ff6bd43fa27cf490b10f5bce774fe76b8ffa5b94830cac7cf9e73394da00aee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd129f8b3e275d7119151b2e7d8346bcc0d195f0f52602d77b2c397aed6760d2b180819b0e052a8865432d9facf61e0bc23e2335665e45e1e6059a1cd5f3d41094dbf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc87354fe1d3f7ddf1e7c54d550924df0b1fa3b6b75e177bcc40a394b6adbba6c5b1363e75b1e38aa9a2cc15d32f0214c30748ae0640871f1f07f63db140aa2ae7b8c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0d192da33a7d83c8851b430732506592ee7f56429218d04208a518c51f400bc7597b93dae4c1226e974040bbbe709b0e3a872107ea824346f89080761387de30e4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e3e930ea316ec1f1f5740fe47c5fd36271a60d3737d1f27c1e66ebb353159ab425a5f9b19fa4b74577cc3a4d33e66af9053b125768e9bc44dd6266b4e8aac26c200;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1438af947184308cab9e1a0dc3890bca80b8fb2b17dbefd43e0ab3aeb2cb5491e02c1bb617de440d7244b23f7e26fabbd368c4f1737c1c900df233f6231570941cb61;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c7f386203dc8ef3e94e31e013f8a41927aad8b09df5314bffc23a59533fd80a2e180cff87b905957b1f6eb04ab7c5bb5ad81114da30e2f5e5025276765b7700217d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h196153b70c67ed2806d886554a8051bf7376704ce3fc47aa2a108954d7d31f83a1f54b1bbc371d483e76751f9583d4dd61a1a5f2fd769155e3c1da6976f02516c2676;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e44a7d4bb628cce32c489daccae4e208ed05cba7b74cbd3bc64a31119b8def2ae9ce36f9d22913acd9919952dc88a6ee639056d0f2083e98ef9af939f4ee3b2ec57a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b4ab813add8bf136c8b702e48beb7772baf4501d9cb1ca33ab575b27cd6824f90b4a04c331709af83a3d2bc1d95a4f304c08a253d77bbe1a540cecf555357fd6183;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e3d5ed0a7aa9cd4bad3bc93abaafc5ab4a50297cece30abe0079fb7a592f9841056283374f78f330c6940bc29e5a5f4851afde7ae0d87af9435009e113a9bfb126da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a9a41a6e53511144736704ad2793a8641c4d4ffd7da554598dc6842be9964c4ec4d7ce16d50ff6f392b53b535d873fbaa95b5ce81592be64d794dd4290fe9b7dc347;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4706b214ab44f45b23d212b5d61bc77e876dfbf33a232dfe7d5cb95cbd04089e4f07ba57f52a6c5f55f5ebb891d4f0ba0ad63629ada922a5cbaf366c3f3be4aee59;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd41296181223c55ee07b9565e56c1b2821488334e2ba172672d4ad763823781e0ddfff996825133ae4d6a1ad4ca5262da672c65919cf83629b400ca11fdb03337ee7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c73672cd3b66eac15a12f97be27d30d45b77b4ee5cc246a1b7fb68f1e1daf958570096ae4e722b55dbd63788fca45727fcbbd3a1cdc2572a93c52a9ac8dd3a57019c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7749cbaa18d65dae2e4000d8335b7c74132be5f25a1975f264ebb1e16b5423588c14ff65c21a0360e0548a0beee90e65423999295d115a9967518fe175619440944d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a5fc573202284a388c2450b6f1c7f3e06b0c90f640511ce35a6ebe68abf8c95cf1188a5eb33dd9952525b2b207ff07de939493adf85963b5b04aeaa30f97c4d314ad;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5162b00ab6d41245fd779bda85d6aa55ce5129734c199a3e84e89775f71c44c8bca78a5e9522b1f0f8ce41a10b7620e2e69e13a7a5db2e09ef5e7e611d098eb9e11;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12086fc558b482c3880c7a2126f1ebcd98e60fb2087ade7473bb962f2276b2e1a711f5b79734912cc6e78d4263d688b0cb62b105a8233f37acba0660169be720f4ae0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ba654dec8cdf35cf236e4757c1810bab7cffadbefd17ade1572f64f24dd6807baf80b577eb508b55f6b3bcb10666b605c3b1c28ace2c29d4e55346ff8231d50250eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72993ed280d936fa1fcb22ae7086809c3823e80562c30ea13d14ebb873fdb4b61d44c8bbcfcf18be72651ff5cbedb4ff9f6adb412853f17dd53513db9db24531839c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126fee6ce7c3d93693e20d9068f2fadcaf9802771389b0030650432cadffb13de312d2750b16328513e4450d7f969f9ecd6e41535c544a2c38a879bcae22dccb2d9a7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1118f70e81b53c4bab4f6ab78e289f7782196cb18c1362646803127bcf126fbaaee8177697b1e172ac2cf95f32e3dcc03598459def86390a6841cf8eba2c805a7d7cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1391213834d89487fadb3068d2197607798fc3fe1f59d1f2f2dc64e4678b4dff67739cc9138933fc936086de2a07320eea6fa1c8198a448998b524b59a9627bbb470a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54851c8bdb50ed35602c9bf147c777ad7fe7e5b07692f7c6d11e40f5cf187895d3b7381a784dbd457e51c25f7fb49ca0c2a7b155ae6701832f4a9e2d6c224e736e2d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heccce025778d808fa15855bb37458586b61eab384e5da33a52af35a3a0892305b2157de0e879b4d703fd3adba610e5145aef8ec3b9e55102e412dd179dded7743f1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1021fceb2f5c3c3ba0ee093e334f4d7bbfc8927e031bee6c5abc6e2dd034db64dd4331368953ab7476954265597b45fb8bc2df915f24a9a53c7166d04ed5013350271;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha9ed9d18490191d4a99008b25019e948b393e407b7788912ff0456d34212faaa50030c7bbeb4f5eda23e33eca180397c2e938114ed53fe0aacd2e1ed7336c7a9c1ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13fc30a41d62242862404607599bc4a90c5ba98954007b28bde6ded466d68a9e2eb2c942ff960f2ee14e3cb271105d3de438a86a5011869641a53d468546f3977d320;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8574f84e5bdbbed77cb00b27fb49b9d62d5a9c12726b383bfa6e34d296458c0bf41a207a000c9abeb11328d0fc9e82526437ef016e4fb6da33fa9760fc17f481e126;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15da0ca065955ecd9d9cd22465f8a0cb87698d5ade526d1b1365c88c5a0f80568aa44f2522c91cecfc22a5536811daa03cad49135409b23b052e29af868e532794eba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17b342e862b33ad07a950f144f98aabf0ed1a8ac3efa6abcb0cff3cc71da2a8db091178d2fcf8886a37ded6ef34673c077c989ec30dd13530426645641cea3da5cc20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb4e10faad04d7c73cc078d2eee073eedfd01f83f3549f4fc77f4579428caecb1aee80e0c02be3d84f8d3a4a23113d6c9af13abac49a7bf243a5a72d6e33e64139e00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17272202b61ace9f77e4c8f6727fbda6c3212c12927e05e16295ee6bfe92a7f5bd010a6131734002ca855dd980d34f3edce95c59787277cfe39c2aba8149fcd2f0a9a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab6cf11f9f374d8ff8638595a742afb657df239ace401d6be484dfec28ea5e66452f51a2ea5e6cd6fe9abd6a0f8cc1af27ea5155544eba493cea2d79c792199395e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc8b3c8dde874d601dfca31e30b8f2039678f29fa264c9f8a81fcbc171687de38e07584a43f02740070210734951b11b55d19937d971effb509dddccef660236750d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e91498d15e591d633c6a7f38f9a5b9efb41bba6cfe722c0329d7ef27884983ae55947df8fbd143c1193c56f7c6bfcd0b0446866e775f951256600076c6d2f7650c89;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h179882fd4fd2cab5c7dd37a7c08b273bff24a66359465e69a2a39355551f08ad5f710b942bee319ea83daa022abca37ebbae9c8b279ba30451459fcd083386faedd18;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd52b18d0e8a2545cc44509e4a10a09e323d656708c36b61e31266294778a0e2e330fed0910c894a7dc6cc34be9442dbb6f4021149fc317fc00ee74409e885dfd2d4f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff2c9371834dce3a2af63d56857576763f7d025f4a9735bd724adc07e98ad9b44fc93972a1fd8f95595dc99006ca188bdcbc5e7ffb6ea69995208f3abee192ee3590;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9dc1071104876a60ac9981fba923ebb9e61f5fba48c944681fec1f7d095846382334a2214d9c8d1f0f5d7457aee02a517b56f29917000590f49194afe835b486796a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5152468b3cb845659c3db6dda0470e8fc53f83242b798d9a7eab3e599ba7f125df893872131242a8f8a0a0bb5942010f904dd093adfdfea51a6bc9a395e98035bb19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1e4682c56f9de1d8654038f3b1fb29d6089b323e85dc2425517a3581abf9882c788629627fb50b732a03bc2859d46244063682ac86fd3c4d76a710750c9cb71c81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1622c98a34cfc199b10f58b7f6d6b59ea4d6d998bdd2686f37d3fd982b1b67a8a804277c8dbc5080146d43d90cba26cd422f1917945ac80b68a158afea6a3c077b995;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h142c227008ef36f1937593dad2a7181c726b5921e4aaecc957b4987c617b49a8eec4a0c96e7126c4029b1a6b9fdf4db6e0a819b8938c30ea6585a35755d45036d7aed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17eff9ee344b2c47fd8c1eb6d7cd763e156fafe724e718ad9d09dfa167cff3fb5068e8352dd1e8c31fc0a126fc829eb83293095d5105d3fade0055f2767964b332c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aec95c1bb47b5e24292bfea4b13c6809a285338eb5eb640487bc9fdeaab848a719735175f588bf9bc71a054b9c4068646f93e185a22441cb25e2689afebe8c1cb685;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d217fec8bc78dc5234f2ddda9ae8e5ca4645c6501efa2280b6713b3fc8342412bf910f5a7b433caab0801735b7e165710db5f0148fb04bc5ab50f64cd3bfe5604727;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7539023b6aba84262adfb5caf015273a7c01b2e9bf03e5f11e8e2b0efc08c531ef181afecbe8d539b76c79891346dc17a168d8151b0f23573786305749b93b0c9f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h28bf2b525b718ab764ced9bf8bac895fd226542d3c0f7441dd1d17950e50de454f29d71c1a3633b48d7bd38839b6b27dbeab0ca36d07cf88d769adfab1094d469b41;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h579a189ab40e5ba943ab3585102198ca409c5336cdea4120620e4ea7ff2e3a46e29111dba044eaba384626b856b334ae42f3b228715b3fd81557b416c13da4de5169;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha06d12a558a4a8739d371ed0be2cec8e5f7812db8d6a7f4feec52c7d98925c737ed59227efbea5c5606e71f807f7d8d18204af5dd446358e01fdd155dc1aa665463b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h130cc27b45ef783b6f3a0ed21ab494796515b2de10ffbf0e5eadf30e868380874a0170fb2ea54da2a2c3177c6a45cd030c2115f9bb4475f69cf50c02df1c4ba6234bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2869e4ab22f6a7c4cea41e89515593c103c0343cc5ca864836c1f651eb6380dd8fa15e0b1b04be62b36f9376bfab63165509c30b130c6a3d3c63b5b47d0bda3f78bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1132b3aacdbfe737a2afb7ac172bec364f2f449639d4c8036014a543b2579bf303f7a4deb5f94e35abf8f9a297ef6edd7b3d871fa5ec48a481b5a5e1509e27f63f9a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h783eeee2c8279a724790f17967930ad0aeff15b808bad89d26082a171e802d69b10e881ddd587858f392a604b60eb6d62fcecc573ad1dedf8c483ccdd1c4e4686d62;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha445973b557a1cebe9fad7bb2ab02e703492a40eedb5ba1aec241bd9e6a99b10e7d9cfce42b141fd8bdf55cabb03539805712827a7ae10a4d2de78b1c5e14dd5377d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd15186579bcd26b9764266ad0201424bffd6a477e2c6295a703dc043d6e3325275842282bf4e45dc5081109a56b7713a3200b712274f51c9999b7be5d97f146471af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1959c82511cd95ef87b83c812aa2cc8acf0ff61c2b14db3a686c41c82b6e16fc4311a2b41a6141e96f78fc690720ab0cd51b623e7619d827c9a5c1d00c463b22f348c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef8fa1ac462857e2f334e3dec8296f97a2ec9ddf1c678e9abb9c6d67e8c7ae16221650464b623837c11e51a2d2ea1241dc361ee7dc1bd55d1ef975b4d7e8e59f9014;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1ee731f6b479dce625c09c51c7eb1ba605d3f6837412962ee555cf6dac283ebfcfbb97342f50e937727f15363ce4c77168a7d6720641019289873beb7173ab97a5e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c3db773d5cafb07d224693e711be66dc884643d8edf84f5220fecd93b4d3b4cb2eed21467f207e8cefb94f3adf87e97383946a18f41c0d03c3a8fe1a1d5888c6c6a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f65b6da1807d3a4cbc70545adf08c69f6fb78ad83a38e5196d63d135394e8d4addf53ef911bc709616487a0d810823927ac1f7481faac6212ccd6d8ca1058d9ee7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11bb8e5a0d15b85ea157e5811d04b6c6b397db02878ee44458184ba7dd4e4ddb5fc1492983948f4348abcc99fbc47101407f2e010090b1b172ca12bd8904ebac8c43e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2abf500a136e18b58a1348556f7d18d3c851d535c83b36b1d857d72fa9b9c9d791dd022080f2bcf96a47b1e2202ac59f65550e8245ff32583cc3e9957223a1554531;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e7fda586fd0aa5146e4eb8ce04316d6beecc86d2af17f502456eb496ff9fa17c28b6275fb362c63aa48da96f650a76d204e3c3e317c97ebae2897508d814150ce9d3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a71d7f6dc10da31aa57bd773d37ca3f9338340c4fb01e21b6b741d500c1597d525e73d3e20cf78714b2007a2a24fc0d2a0a4a377542d3a744d3f95569f75a307d2b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9b6e198ad1f5438439e08cc92a0b23ad69c5b282c7570b61d761e5bec7c3508f11a3614d8ec01cba2a39334e495ccaf2fe2209b46810f63763509cf309d89a6beeeb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12ff75b1c81af4717961a867f6e642a0f2eb82900e6c8020b00afa1282c375e3ad5ac8ee34d7739b602c55985661e4c722a4c7a7defa923ad26aa01526fbaf42d5ad9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91cc4113b81c543231a3a153c10a82c542316c8387fd31f3e7382db88a6ef06c118fba32498286dc4ab7e8c3adc3dc4cd203f1c58d8a97dde00719b6713b3f222c83;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h135857acf097ec09325c0b2c1e2fc1e3c9998c7f9331bf6de82a34682976f5c4cc23ccc5144126d294eea4c800df6484141e448f1f061f6111743471ba4e44142f330;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80ed6f02355c6735fb3b7a06f910ef2e926fdfbd22689d20cfcb421239f201850455c33a84ddd009b15157432c05dd865aa99b4d376c43fcf8a77b4059ccd1625326;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h619e5bc78ca7e8377b526570c935ffaf7e70ce811ee53c3d02a98f09fc1d8a7dd952b2315f61da7fd0de603d79a3697a625b035faf1b9afb3cd4242560af85c38fbd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12c5314cf388c9c07303b75bd718efcc93524df83fc77747e1290cbbf538c1935e66d52d3351c3321448895add57e6346701b6ebdd93b0082a98200134381db0cde05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h363c2c38cd5978cc13fc26b79f809f20c407fcbf53f0375d2fecb730ad52eb32823c39696d941fe5fe155df24b4af13d2ebd6b5338fd21fbe82c3eed32b9d9a03349;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf5c0e11f22334603afcce34b6d23b96004eef8ed1ae7073e78be8af1e83115ec2fe33628fa3e66edb4dc9928b21aa9e3dab9be145fd01dbccab0d8874ed2a6abf714;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1318022d771f8ab2412544d2529eeab5ea36f95449644d5384a2d5e7c3cee076eedea833f70b803dc453589968b3629eb729e9a5038cbd1e4a5af5cc2828ef108fde4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49dcdc05c2a2d160ce9418961901880664e08ce150e92263781af6e9562a1810204b6174ce1cc2a6d6f4ffa8a08aaca740b2785203504641d2697410b138944a5762;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bdb3d0da29011737f8b97a404a2fd3cf616d950fde238dd666a545cf84a2aab15e636e5870f28f78d03c311557d25694bcf9bb66933696a2658f3002e283da2245f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcf9deb1e1ca5a9738fcb4fa4636ec7582db57b7b5717b5530cafb5ee6bfdf10763dcd334a6dd93e44dac53a8149d30c1469d275fe03b2d286b0cb958b0627c828890;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9571c5fafc77ba03cb696e4de0b8d0a8b29dcd1143968e5397069b88bf109e993b0bf109ec6d20e6c73e65f1afac648c8359eba2c69bc42550158de0ea33eeb691b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb531e25f8a86762b6460018b43ef4614790101cc4496fb94a46bd8045d3546ba7a0fbda7259644e51c5ff40d4b32ac01689e8c8ede1fd6ed934b04721b403991a349;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a71ba279702b108c52c9665a96328b63c083257a5f8f18379c67432541610d6031b40ac850c9d6e45e131c93aa340785e13d1e06dc5ad7ab800bda27711b053928b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1138c55515b4346758bb44edd41d288866a07b9d7493e5c3d3e641bceb38e04dab64b50cac84994a2eaba600c739c2f88041e1bea4b974708f4614e14887dcacedf2f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf24c999aab93efc59305eca2a842df931065cca0cd4b7c2b391585adbc5a707498dcb99e34e5cf362e0cfed430659fef6653945522e00431e26e1f9921aad6ab27dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d55433060c048ada41aed0d336fdea5cd0200d776f0d7f2343e9b4f6c9c2d470fc0ee3179b51029dd584339dafe019050c6bf005e11d0e7ea75c77b43e8c7ec1b57;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e43b0db146e321aa998f4ed1dfc6222a2159a56403e4c498c7a5db4552a0da72d3495a552c960f324b0e753bbc1f8c53c59b67f14ee23d32287308a255e597c94b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b87df4160d9ec00d8e92aa2c86370c0380e8e2798e0e55c64eab46d67f0fc9803d683e1cb6f043cf16c54f1ee2e8c437d3c67fbde9e9ef7dbcd8f671293cfa2e7d33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193652b3d6eff935107a3c40a7df26a58d1b3a039af55cdc4ce785e28eb83e40bf3b51ea59704016589af4a1aa820ec97538a492ea8bcb49ad2468d5d98512609691a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d3f739e89a85a26d8466dda866dde6587301f2e063c6489820820b38c7b173cb18ab6e43ceaf8620c4901dc7ab3d0a3c7e2f02f16a468d22829235380957db9289a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe87231b351b4d69e708ecbcd9ead79f014ee5bca38a8c68d8ce448d7602488f1bb184bdad908dba2e3931089179f31a18f552aca9d83295c83802535cd40a63055e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7b6dd4d0834363dd684e93155bd6b97e71493350aeb9a592b42bd380dbbbad6080999ba2f485406c8c3840fff7a02ef71acce6f56f69a6c13cece66dc46108dc057;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6fe53ef05ef3b5f94d47f99d93caef34aadaf1705b3beceb319abb407e1d9165dedf4d644a62c1a68ed9d7d3e48b26e4b5defb8b16b3e60ef7a7d6e08f6d98ed465;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c1fb74dcb2d5d183ecf5234c40a75847c5ac6a5c498bcd0a59841844dc268ff1c4f3d8a6c6e699c73a8c8beca2611c55b6801cf2e0b7c979dd533049ce41b0f678f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1718ad331e0227899c1e19f9250b5cf7f5e2c5d56c9c5048a39bea7b9f18f55967a7bdd5443ecbd7a72fe5f4b90354d788766b16acc52cfc1c43e15e28df33f462c9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h414db9134b536b085f6fc365d39aaeb1c9a08a485b0d2a1ff46000e353f952103420dc49f7fc48f9527ee495e141b7428b9048367ef9334039be56f5df7e986e83f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27e35f58278e66c762baebc79b7b4dac7621650afe220d6f2fb7d17aa7f2a5fe138d865360110a3705fe2a74ee5e935b3741450741d2da9960a63e09f6ec97b26bc5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f9ed3f1316c730991ebcaf4ff76c9b9a3b4fff1e9b2ac40b739ad43caf52601562b7bac343d8c58aa99387f2e9ad0b386f5ac86d40f957dfe37d03e68a69ca4894e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9c3a5fe1bfcd29baa793f1cbea67e14d21249437c424a12999c54600781da77bd878d54aadc615096e6e67dcd9748e1197b3bab04e7f79479d8c9e05bb7e7137ce19;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h686978d99a23bb644200289d5b178fdcd058e61963282a59e717f91c008d0ed7ca589974b5c898bb60e4428ef27a72a4842121832d0b41b10fe720a095de96200ffa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a9495a866ec495ef5e57b3f50eab87e5285460e1782536e74140043d845c34d4d354a860649cbf21461b9589fe13d372a5b5d35ea746b31cde799d2bcd68f258dc40;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefb48212c27a907043f8e19a1be0bc369c5c77851d44e93edf63fbda50903b8d3572b3a8248c062a9ca6087494b0144c6f6d1099115d9eafcd4aeebc8d325c31aea5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h71877623b641afd9af9c79f9d2f3d6b520fe7f853832f684e075253560f237764267830705cac27aae1dbe4f98a6207ff827bcb7519c2593d3664866ea15f7e7597;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ba5b33b97ee70751c1a54694f2633137a96e8f505f8249af7df08becfa44ae716a937981b3e480bbe340791fa4e6251dfbe462049886022141a5f3d4d8608a153115;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21c31f7989423ad55efc060912aa27fd883af7cbb7c8732e018aa4c62940b7ed23c3ab15a78bcdcf152632d8102736c2b1cc62ddad28d192072336dd4986adbf97dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f1d122cd72734d476b37bf241e9cd87c7d6ec9cc38d3f5ccbd1fd818794d3d83b0586b941e1b4fb19a896bc1d256465d96dc033085a8daff15a92e0f03bf4b8aa0d1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9848b5041623ccbe30e514bc4137dc53e6288607d501d85fdc4b43af3c500ba6f88b3a6aa6edba73d26f4cb9679c1229198885675e8e55da471fdd68162e1161de6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd855c4c82b1bcd54c9ede49bb52bb5875ccad3d9e5d059123eddab37ad1d66572dcc15967cca5d49314c1cc6dff3074c45ead9ac5e090cef75204636af9abc5e83c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h172f6753bc431efbfac50c59443af0da54b9365f7f1bf304124017c9e37108a60aa3bff53e7fbb87782c2ecace04366a1ca8a9d7175447be8ae803770e73f8623257c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e236b1a7c5efeec53f09cfe0bc6ca8c1f12f307cc5285e2272bed5c6783d7fc48743947911331383f005de281b71b43f0536b5dc74f983cdbc8e65c36cb48c4c6e66;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h494d98f2d2d00924f976942306a9209b5d2f5b779776d9aa51e8cecef2d4490ecd1d3cd35e344f997dd7b2b6a52046391a05e7026f22f3afcef4680ddeac5fc69135;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea8a54c45ed10b3e5f92dbd01fa8e9f70c308e20bf3b01147c0caf955d1b94de4a928f25028abd0bbeeee7276449518e8bc020da272856fbf30718372bde8edaf9a5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edaa02600ff3895f7306c77ceb7975b8df9ecc03a344d68a2d8850acd55b91450c08cbbc36963654c72cbfc8bb981ea464fbb0200c5ecf6655854515f68fb43d40b6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c7d2a51f8892e9d7e7729cf9e213f4948cf0dda35bb96c2907865754099c949a4acd362727b34b8b9014fcea7d627b7ce3ac6d0117a146b241d04baf0cf458982d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h571a16395f35d4dcf7456e60434644f782401f6d462c49f94fc32080e262393f50b54f62f8f51163d198d0eee9c120408c3336f885294bbbdb82d59bff40832b07b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcce6740d613edc5b366a1eca00dc08784b05b5027441fc20e195137ec8dc2ffc2b351776afa4a3c07214d51b5725671e401c6307eb368d4a5646c5ac6779f539571b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c17f74cf41d7e0decda074b913aa396f6d53ab46350f84892b895ce08a3f09bc5ec9b1b81b6eb6080cf29b1bdca81f335f27a37d41306db64f720e4aecf52074b6a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15869e15089d47021edf13cc33150ad49404eed961d89c46580445c5c7d15771b9859b1efe27f1edb4e106b851d1d395d6ca46d8c24ecf2da10eca46ef8f916d42453;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha70557010a0c80565bde69eb674097cc1f559876665597c19f20f88b875a6a7a716bb01978ed44b97a3d89b07027561bd10ff55d65df8796624a4686bc67f32b5e00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd288a15215ef833054459525e526204170ff86d458617a74607cbc56dccfd10ae845056b9998b6b2f84847b802e3e4f5f69ead73fa1ad8a158d2ed8baca5bce4d83;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd436d9c74901a13114549317e2f2489c97cae77c3998db122807d0aaf22b9dca4f2dd538de5ca4ee8a3d78ec456b149a1c6187058b73caa8d081a3c0211414af716e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefe4481209e77d36e2404fa77fd709e0783adb85b10a346cf9900923d2f66dcb77ad118b76e73b8ca52f6dcb17d3253e548d4d0814abc78d88c9246743f2150635c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5de9b9b963c5f2fa4ab7f0b187a5164bb2c6267f4e9348dd42bc1ecaa81e1d90896e21a1861ab087b23dbbe4fcb86e7f607f788476bf83d6267848edc3c535ca4deb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3eed52ee987a05a880e5c91c04c36782ce468882ffb5b084656431a9fc03a0bf94b1ffc036b31620749cd0e755aaa8f5993eacc7ab9a6fbff032d05cbf64fd5128e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d3ef4f96d7dc96cf664a61ac33367b8909eabb31867486fb1b13d1cbadf20fd60a072d6ca2628b2f17703a3fd2b4eedbf740a95c827c539ed37a243e63ee5409702;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b90b748bbb1e0313e52ceaea29b6a13b7f422ac42cffc5fd27e6ffa750a9bf8b0a3e962638c592b75e5db466929ab13c2320a5c9547779206a9b077db1a7c02eba49;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h119377c443c2954458233a7a8e974db92cb451c3e509045954a9ffe9a1bfb57f9ab0d8ed894689141d3235ec32444306e14b9dbcdac1b9e914196c2dd30a48c904f5d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f35cca2b162e49bd42600c1abd10b0465bca61f60aa11a3b3a0c756701d2856a088d96fd21826002ffb8273708ab6bd351d14428c6be47fc1aed7ccfcdd5ec126a8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75cc8a19ab2407e38004de70313452979c0981c8a1f87a082c59fb6517d5ba62da36b9d410de9cc2c633f6af8ad94093f1cee3ee75ebb4c9b0c03726a2b40a3ec610;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe14d1f7b85b5aea3d5fab28a3c97f8e848198565fd922bceeb94fa0c9ea6784a23b1fa0ca4fa50560a6d54c5008f52934a4548f2624e7f61f478f4a141b783804d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15869f5e2d4899a516ab47a8dacc91215da781a1e036c3b6dac803f6b5afa2df974edb58a29aea433e9b49fa37dc66a3dd43af2d5d6161bea585bd5915759ffd7968d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0c7411a13f546e458c1423a375ecc77e8f6eba4b73a6e79fbf4bae87e778a486936256c39c24b92c328ef94dfb13bfd35d8f7cf1d23745e53b538c1ab93864ba20e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d291fcd5e5c7975b07b8bf5bacf935399d93c696b7f207d93a0ae509e59d9b9f118b1a7bfa318cd234f6d2e56a86ab84a998a023366b72815246468fd50f6cb98996;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca8d4b3ba5fbc2d81f277a67041eb1f600d71cbdaf06a9236488107e4ec31093fd212f446700acacc1ae7ebdf968963aa88dd7c2cbf7da1eb223f40e6a3b40e98f6a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcfbf80a04a773bb071a44f53e3555f49d27c68ad51c6bc581d7ea130455d3ba5d703f005e8a6248b90fa6e4d6495ad66218ad4fa0363eea51e92a9849f6af176c7f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154dc60c5a0b17aa734fdca360e2f24ff95aab65617fd7c73300319948b5bc37cf5887f1b40cf37dc7f39013fdbb8c24b1944705546b498460195e42dd1ce7447f9be;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15f3ae63396b62f6a863752940187779c2df92adec1830850598eaccc1616a787a0543c426f7782abcea8f6444890d22c075741a715136c56caac7c6c043f045c8554;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12016ca2e1f5bd8cbc2ef1c29016b4dccc3bab7b81eb3987e463ba9f6ab1e67e317e10a2eac73a2ceca27787ba9c4564fc6de85f1a1dd90cf33b7d3096a44e4544501;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91c91df18a538cdb0ea46fced2499849a5ada0ed7720cd68ff17ddbf2ad0f817f5e412ff481518a682cfc3d03c469fa72556eb8c1fe77763e7a92c3d0720113da19d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa8cbed71a5f58e250eb17289b67a3d0fe83d2cd63816b636c2d9a316860a09911f73dc79817a686c50917b3b13068e32cdba4d2b2affc06deb8a992f18a3522be33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1939dfda975f3427c1009c1a1bd1dcea95afaa4f9b160d8598c2bd7a8396b29d32cf7270d0e0dd9d805c39cf4092c8017df6867e16697f30ae1ae4b0afb6a8b182d26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6f62e92c93ec747333c44399dce87b46f90dcf4a0ec49c9287ecaa884d28df57f18a87235fe9daa2ff6f8fc2311e9e361649096b56a871ac93e21cf2a093fdc4e060;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f61f0033a7d5813045fb978075df8b851040b1f24ccd371f70081eb35a445e345de89066c8970599a6d036905322eaf042f53c3c211f22585aab9616628d0a92082;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h396aab3b333e4c4eea49d08943efe6415f35f03ef23564d2a8714b47bf224c8e8f50f01bf9e1223ef9878a320e9381dbc932cf7accae0b14aa1d75c4c3e412331600;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13da0633eee8f2ae423651d474e95f8ad6c66b017c0733ff4c1704aec7f6338ecaeb8bfd4fff0dfc44b595fce91cf47b4c687fd05203abf21d4d5424619c1ab10f4a7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1234ead73dbe567baa1b539b82a6b691b501ed3aac1377220943bd1fa6f46fa19c6bf76389a0e416e1ef6463118e25918935b907342a6f5b3eb9d4509ce5a4c11aa21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfdc61fad24eaaa09bd902de7d140235d9e7165a739992e38e9d469c2240b5e29276d7c57ef094d60e7e42d9b7ac85a9b5b7bbf02fd7a9992e391821dc60bd3e4a8c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c3eb20f9cc872901903426b8cb3071523bed6b3842766a05d3744e2d7115ad08e096c146bd88256ed6da83253f4c156249011391c246998e22095539902f9a76272;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2bf8d7af445407a9c5aae7808996abdc8f485df62b1d99c27b071aca52ba70d0b13f5b7ce9709a9055a707ad3bebb2ac1c03d1acfaaed30f1905c3d8657aeebb2f1a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e29b4a9a3f3d53889609b35ff181956759b43e44854ebd285184ec866cf6b9305d30f42c1516f3921473cf4c649a331ddcc01f5076defea25a0c983b1656ffcf71d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha32cde2c86c06436d641531b591e9137f5d94a5c8c3b81b05e4d8b3c125ac58323659c67f00700a0d5992da0aff25c88daafe7d892646411fabc9f1aa2f05ce561ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb30e2e88bdcef08d33bd7b0b76d0bae38db36187c84ef2cec0e1b34f45999e6357acd45fcecb198c10b0ea4a5bbbae6d42546e668e571db0bdc338f2b7ce649da1e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hda28e15e47d956c75331163484850a638bf2316c0742abab102191de151468d3b71168ba90a9695f8d4635d8bdc025dc0d70393b470aa134e51fa85a73742e20239f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h876299af2ed3125639538c8479df7337d5887320e2ecb98aa982ff166bef618019cfeb7eb6bb46736f0ab904bf0190cc0257294d53b48b4b08e8a18186592e6ce795;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfccf689e55ffebc8717aa6100617c979ae5145a870edcf8362d34899f09dabd2dd939908722dea1090f1b31ae05b8f2f3aa0a9dfb39c49843fa0e711f3fe9746164;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48577d4120e228c4730802c8c7f261861ac5adb8ba7354f524651876cd4b77e2e85843d32393f4bb72cd552da288a19f4c5f83609dbc39a502ce5891dfaa8c24854d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81b6174a051970ba3e053f191024a5d22dd15c374966bdff9f6617899159f795620e361a71a4ad7b249bde66b8c6b71be8d933b69d05a2f65d4ea37eccaefd4eb128;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f69dd6e5392d61aac0b0e9226f547a1209326b541d9dc62a4e4fd4602508577c9c4e5bddbf742f50d4b74fc43b8590b390cf4507baa3f53cbc2149ae6df09a0dccb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h346fb6f11186b0688893fe99faf68417e7609c8c7deed8d287414b588babc315520b5083018c21b66cd7cf7936de9ad44f3a235f111343869213b12e43dac31af386;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c1d8d20507c9ce53e3a277ac6fb4216c9a9abf1bc6c15397032d09b37263b057d40643f29829ce89b9b3c6e544bb84d47cb5e505eda0c65eabe08385ad54c330e4b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e47631c08d61e947376bb0ffd39d8e5a2a7d7f27a780433f29000459bf5acc7acaf38b70b50c1b1970707e5070f71d940935ce46121f3cf6c8013aa2e1f93ff89234;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h883200e798fc9af3d4e1b5fa43d042128ac4ddf71a8a63d8591e4e12cae2848c4626337907feb7e7f4081e74328716272a78ea918fcf9a99afab6640bbae603a06d3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bcd0c7a75145cb60b6730ddd7d09f48c7d41940a381975619a60eabaa810084ac46986e63db1f3b42afb9286ab662ead723ff723548cd52c465c4226c61a251707a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60d940d71b2815adffb3b900995e358728a60d08646dac5ae0c815b17cf7468fcd3f6cf135304235a6de8233f9e339bb2816d262c70fcc7450ee0e1829a6c5f040b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86f96587372aefb86d2558afc22f607e1c3ac852f7c4b0cfabe0640899cab2846b151589fff1f565e3a9c1d4b53dcc47c4034817124357b5708c3589455709563586;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa6677e662c042556e5a1c3ac560705bc34715b74e991b70068936ce521cfdfae5427c25122d2a04d3d3408ffd109b50c41ef0c67c3949c5e7b16db305d448e8b8a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51735f2731f87b61c24b937ac555fad9483e7610e32ab637d34f01c754f64545e890837f93ddff44971d2794c7e72af31ad716b4488643fae72bc2d4474c9ef7551;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a32a1aae34feaecd84da7a682749b1652def917c14a8ec878eb544099aec360ab15c3bf79747a2284d5fb0d4b9141832d8041b7fa0f8d32a37df01c13f4df6b3a27;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2415a41abfb2b66320b815b5a481126ef615b3a2b1812dced8d9213a9c621c0acece10436ada2a0eba26f841ed0501b164e4303ce9a6c8ccac333ebf04e3afa721ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19f79b7ae763b6ab7fcba496f1e51148a896c055ee062686a38252a8790f9b956ec1820420a8f4f70c6c5730233dcdee81a3b2f49c8d4dd9357a5cfce9731d85d397f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8d13357f19675389842bdfab0f6aee30250ac7db95431589ae10db687e9dafa6410be76b4908f3bb7ab0d39b1bf545986617f062a40066db51e4c23228fe749ee945;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha7138aff552651a0e974aae2b76ef684de870a5d9439fd5dd935a6221217eff24a5f806868f5f73f1c99d47c1ab7f5f8d16fc5f65a30e414209121482e795fb0a170;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h123c88c76b3db75ea17bd7c4a435fe4ef2c8dff1b42dab24d03b0e2baa3bc0272187611c012f9d5c7083af58120937c3e150ab11d4cc976ee039657b3082903a80258;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hebae140e5f5bdf16cbb2388ac74ebdc2ed129a74ce39affb535bb0336ef76f21ef008aaffc64624fcbb912e4a9e7bbd979451b6ecf067d541b6735324c2db83d016b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163ff7a484d97b6e1f8332287f6927c82acacc12319d15a19528bf1d830bc3ef6e7581b3094c0d10d72ff183a3f1a195d77004849d59868bb4b129cadb8c9619cb5ea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h162a616f5d0b4ad6ee89872ff61f812af2b0b371c88c356b1fe2028fe84b2871e8d388f570fd90a851c2fa002fa935c67fbcd93b47b02ebe41246fe043af991fe933a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7269fdd46357e9f50a2c9c83c3f686bd79a4888666ce48a03ca6a1632991edb1c3fdce2f224de1590d377a29ee3e3bf0b3723e50d6f8f1ef53f51aea4d9b51d2d645;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12b0f761b57a836035d030fb5b40028543c21556a52dacaf2e3ee7efb44171428fc3a44acf4c8ead3ab1fcd3ead1510684427bdc3b13785b142612d9349067e463dea;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a2dac79ae9d1b6970cb30461e247f3cbbded74f585958ded08950c9c738542d6d96ecf032e81c383296448183070f3bc04a0d4679ea317a204c461b75fa728c5620;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h705b724dd587d9aecb3c0dd8a68f47dc62c46e4fa8d4168604979a5c6009f71da67f8678dab29e45d83822ba2fc56e1e75fb7364d1ee6993956227bc0abae76d850d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcbdb4bd5ecbaeafdf435583bf60fbc3b2229d43ce7aedc414366680277c4e95c3f1db7cc2a5f7008e5d18b31f0ba51a27ace21b05f92e1af010b3987cc06abeee46d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c24092b4910fdfb1d1a6858eb22e018682dceec4aa1512ea2f4a4977474a0118d6379fdd0ebd02a1a21e93704c0f29f75de1268b6176d6f61334cc51fbf6ac5209e0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1c0c6944b1b15737877979705272e1f439c75ead43951bcdc240a40b3d60c12dec1fe6ed21a4633401c8fc453750dcf49e2ecc9cc4cd7455300d1048dc2cd951c9e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1774f9ff47b32f6d2709316469f5bce89226ba22482df2b59f25ead5e6174ff1f36ed08965727d8994bc3ec1b667a17fefd4522b0fee77a2e43eb6922c876ab8d99fb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1794478a938124bdc0f42be066190e1cfda54006302d00a8a62db7336ea90965ad3a511a9dbaee72918e689ee38f6672b5b8b516ba33a0ce0a1657278dd07b3f8cd9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa0ca58990283defe6450abd14c291fb98bcdf513f935a1e4a88e42576357caafa5473f6668eddaebecb0497ab386839ea60333d2160567297c3f0c7552533a3131b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1598da47c7e4218d49de4b7e87707aff041356dc04dffc183a7c747811502161f5d56b5df6d1e05b34ef0fc8aa0f9a4a6b1f40464a2ecea646558196dbf6d0e92a991;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e920b1bac695c75e5dc56627c63375be2e6e1a44ec09e1fdb57046dd1f26a67ee1a32ed278d5ddb22ffc2570053fe8942da85085736f7c8d929a44c6d71fd86e6385;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e4ecbe7eebfbf08a02eed327d4ff2786982660cc4a9c8edd915901b2c44f500aee0365403d099f549b008e24fb814cc9138d2aba8723077f96e4afd0b6d486243d70;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha68fdffcbc420abb52404234e107dadeed35d6f9b3b20ef0b27df36f37d6f5e1533b7a805253865837ea36ada5f34e4b952d0e276ac675b2253c5b533cf540f1b6e1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7cb43ab96163e1f24d5f67c7cc00ddc310df14d287d3d260effd5c3bd6c46f16da612ea68a425d25a442175b7f2d1aba857b6bf46c01cd546d5a47da6b99ac1dce2f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1650aaf9e8c5e845316f2df9a3a2fb6cf0d468d7c9a3b3d06303541a663e67c83687746ae1c60ad5c02921a4c2b70d6743769bb2fd25157a258d56583d8f394408124;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffc3b32cb660ee5494158547c0eff4bb1461b88dcabd3cb7689af9bca4413c26c295c2c0303f48b047b2ab357f5c3b3ff7d79fee01d5f92cfe3ad932c23346028636;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha712e0d21ad02f3d966e398dcb41f7fafb271ae2c3e35494fe83aa3bbbac135170a5d5e3395c51a11e1a13a54e07c4bb502199b36c8d9a411140ddbc60c2f2402499;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138364abdfc43210c65248854617297dbf2f310c7d6b27e59a64a6936337cfd9c84cefe4e9c8fff776a382b3c3e3e0aef0341371cee923d2995584caa3ebf600dbe04;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a06c0620efc2accdb394930ef5fedbf6a8b25ad0709acfb75d0d2768f82ed918dffe129f9df582ef7e6d870d11dd8d3a779a65433f05e364329bb9995acfbb599f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d86ccde430b6d9f3d5ea2f9c7d0915aba44b4a87333fc7353bc918c5fa5e2732abbad7031df0e496863f764837c19d5ca3ac5ae4fc1da459019ff54289add495873e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da6b5d753e073adea5d05f1a2e1c0a167d4d3af83a2c7c30fc1ba0169b1bb7017ab65a29f0198c2eaad26655659e06a802318a99ab20af9a118db6b8349eb07293d8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c330d6000ad3fb5e691cf0dbb51dfb2a1169eda45804ff7aba2dfc9ecfb3f95d20c1ac2945a7bed89818dd585776fd01e0a2eae8eddac54792ccafe6c077ab238da;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h91d12fed30dd91a89a8044c963dca4efb5edc20e7b6604d95ca15173d56ac384133509db1ba65244cf394b3189697fc204f8412de8e6f9adb1930a6be64a2aee9a4d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h160d638d4b688ef22440ca75b289ff663688f965471a10ac97508f596675b06ad356779183c43b489b5e654782f92c090fe6a23827b0ad64a3ec77116038a41afed74;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35ba287ae2fd1c06d8002bbaaf1847bd63902a23c7ba3bce4f1bfe8a5963fe86e8162f5fde4460d24a4f26892727e4626cea744844111f59e2f889dc0a69ed723e26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bc61c98ce07360eef6626a8556df41622d071a38390e00249648cd5573f474c40eaf7a8fdc417203b3fba7b7d795e0a36f047aaa0dff619951c2fd360c950f4871a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163e0705fbf6a965491d89ef537dfceb364fa8c3ac5d63e5956808e6df698426ca2080b241e984ef97901f7631020f3530b3d4636189fa9e2ce379a241d6c94451988;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h106c1877c6dafe8500c101fe3ce0dfd07a5a7e28635b88cf482ed70cad77ada3376550b75298ab26c29698966f47858d594c843859c84c57e66963fc34be98e1c4708;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd9dbbf388852b66c645c894f918206a3b036631573bc4649a7be3916a806d9c9a02249a0c686ed2c8e993cc6ef2231f8332c6d4e82d6a0cc8ed4b8c69638ecaef87c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h22ceb8e1027fe69d0c3758889c647ad7f310f85b5fdc95828d9917005719ca6cd7c5221df6965833006f72daf74ff79d9c5f0fb0ed66f263a328604b4f7b72ff7814;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1916ffe4b810d087e11a8fea0df71ae7f9fb6789ee59af9e526705e36b82c8ae8599769e3aafd2298d65b61dd230b9560bfb53b4652d8bb3ae22630543f9ad54cd029;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1439b91fba9ab9b254695fc6f8417283b662111c8eeffa958481f23fcc924f27fb1c3cb62b3289781357a1394e7136580e06d3394bbc343d2e569180ef0a562a2d217;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13144f090c3979e498adaaad3352870ba70f1b8de2789153503c56e655bcf8f35017df7df58b38a5a4ba20078eb1031684fd07efa346b6b5257f62f0f7af9439fbd15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3b91bd5128f9ce7de698d596030352d201254557cad08e1f4dae3dc91313847340c8ac6c136a0ec811ce021035781eb6a3277804eb49e4aa7a228d3a9358f96e727;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171693fd7d0e7c1b577999665863abe7f1180dc2e2b3acea40d4253b270b8f2fb1032309bd67dba8c9340ccc70f1a8ba12c5a8e9e9a7f53a184938d9e78ca8f6357fe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b55d6247c15781e7346ef4e60e60fc928d00a3411d72d0410759698fcb7d393bd31096acdeab66832fa1ef24454c74daaf5dad7a8c84a277e2a6679957ce592c8154;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef9ecbd940f8a4cbfd7c454ac62bc0903e47ff05b82d5d7c5b9e891375b7c009d99617a5e593c3ea796fd688a5e0b5de3a834ea4ed33ddf24c9be242232b40403727;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc49ac06c1adf8ffe0513cfc9a4f665d52bb60e0d8efd78576394b42cbb7a90672e21f64e3e88db6ab8e699a903021e775755103336ecffcf502a64789655d69b8d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d860feb512dd6fe264a58a73025b0fee35f1562179abd7bb0f82796373097a0ac82ebd62c9a2c386305a98328925d543a39bb52c8c6470af8c6d76c7a57ff8efb9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ca4294d0398940e53ba1ea59895a563d6971b3b59d5da673ee05e6949d286e5391cd3393fd5008229ae059f455c2987434befaaca86b9763316d43acfd5599909f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4092353fb6eba109fdb6555e17bd6102c988f45e6cebcf1a07d95523db827edd8de9630ff53e8faffc9f1396924d4338575c7b66fc211bf5abb2863710ab2054bc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a007c395c0338cba4a30522b375b7bbb5b2c8c87a26355f8bbee7807193d9f0f804f117be202add5e0bf0fcb7c25f4ae40a6c57068670fdbe08428a1ffd2c9f5c307;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dc61e3ade69676bc884a93f358f43df0f5e8850d8bac300ebcf377ee3973b86729f9f5632c59107e4f011d41733ff219c6aea065792096f90aea07dd74f83d893e9c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6285dfb7559e4c63163dcd6cfff25f79e976b62f2a489a9983be923d4db80779812aa418bd08f56427331fff9c725e47190a5664f4589d166a33f4906a0b641ed1c7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9e390cd3b651e95e7a60c6421c38f752cce46ba67bd83840ef51cb4ba0f9a55b5d713bddef7ec94444d0871f77a05a6f874d9c7fa1689fad6b3b06820f6452e43d70;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9dbcb6a2482f67ce75941ec3e8d95463331a3a4402ea6c61d267b95e59a526b0c7571762678423feed7888d050520a84c304b1bb4802b1762f712a2f953e0cd8201;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb4f90ef77e4b3cebdd7a61881307bf551136e169af20c9ef03404d511b5a4f91b847d8b7acfcc4f6c3f50d007e31b0ee0411d077ae345c7a7157c8f868081b1f2b95;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171c5a38f1124b610b4b39497942878b9acdb8581984b99531bacb1c21748e411c7e1362095c851092b8d29bc5cd480ac978b1ba8a99609fc261594964faa2a0e950c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e3683d5543145fbed8c577300a0caaaae3f9967707e1237933ab726cae883bbfd7d573aefac17812d161e72bd25a461e5105d78a400bfd4c577ac5f99f99c45c916;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f812b335a6a66ba29ad2d4d10c2ddd478f27d725ea047d5aeaca22acd3885dae1ec02c0d0315f4d4f0d276445c3adca8ec357c38f14eec328df2a34a16579569d66;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b9887fac725f9cdde5dd3da3f1f1398622444983fb4657ece85bc540e584d9e707dcfb849074192687243d0696475d9c51ff9ebb3a11fba44d4135d95a8ed04781c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h202a21450aa7ec04305534855df572ec636f6579b733c7e07d87d9d6b78ba8c2cbddb7c5a8b88cd4bbbf08014ab413e5a72ea8fbe8ab3a6f76cf98e14b9898e0d2de;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hced7c7538237bfd988ce5d7242348a52a24941c875286a81e40e7653493dfaae961e87421b4b0b32a024bfd38cb26c74f9cd9b998b431e0c78e9a65ed95a085ffb84;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed3ba69bcdefed3072c4da8e531c612b4b331d305543212a0ac5077a4f5dfaaf662ce1ff53a9514a7a6cde8dbc256cd842b7c43ecc54d7d02ac5b69e2309382edacc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17564c8d06e6bca667321f202e98653d9d6aac89873202494adcf9fd0f14ce02662896e7825141e572d45ad1baa5b3681cb18b73042dc802c6e2ec70e9454d3dc101c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5414d9207abab1154a088c66aacf4df24bad1c3efe01ea20ebae9ca5ad1a10701886bf4770c424ccf5bcd8385902a47663c04be354ac8bba5a9f558b9560cddf9e99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf3dcb597dab7fb34a62d94e9ea212c60f5bdb750bb3bedc0d5cf98f45da0d99398a8a765034ccc86289196e71e17587c4df0b20157db8ba015bad25b103f84a5893;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ba5da1fd296f3ba8a92c71c3a433ea3599dc16fe4c1934f3b9e6760384021b6fdbca212b212e2e408c949b5ad2c85d7502ed05db9e33fcc36da1b613b6e58fd8a9ef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126dbb11bd30ce435c97f6f4e0567e7243241f1e896d1ed36760040a11e9ba3845681f8ad446a180518573bc1506f0fe6bd54882c04aa059d80f9fb1a9ee2d7045c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hada556337c98f5f93673e0f8dc7a048f83b45884711743e11a2361151296b43f132fd72f62ff4aa841794edb4c9dc29ece39e24c0f2ad23d16750a6adaa858ecfc81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e339e497402007b29f0aeaaa3e63f1268d4f0fb7838f1e0080f16705d8cebdbe02196c38aaa35bf8f69298a835193ded6583ef6af3efe2b3cd9713562335e5c8f918;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb0192ded69a4fb7e02576abaf4184d88c513238ddb1dd29f5a08fed5d05a9c0df4c121ddc6442dca00e1b22881f4d905241daa0baa999b5a747824bd8d134ad7a8e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17e9a191890e0136e285cd6fa69cfc5e7ed6dcfe64b95aec86eb54f4d9fe21650f44f899d5dd76063738f04c7a4934872ac50c776ed87b75fc0eba9b46736fe37dde5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170ddb5b1f0b0e56d3bbbe1c36cd67ed8804941eb05384fd9de21633c9eecd1f4ef9857a98f950ba21e031ecec14eded22c8f0aedd52f5bfff77b0064849ff40e2cbc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182fc6c59500008c2ff8566565ca20d6612272f4fe22c48000955716482beeea14419450e630bd6e73e240ebeb7652142ec33e4aa879750f32407c2972939e1db4659;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haf9f6cdf8265c4b739f3b31c2b9e625c7ab2fb5a74f3f073319bf4d9ed69decce3d3c93b79214d991736bd5f5a6521cc5107d38b66275ddd93b6aaf25bde199effe3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101fb43b430f2573c531bee1c0e585f5b65c1dd016f58da51860cf6e7d11d44cb3dbe998a1b42731c0a34a57b7001da23e528379b151ed7f91b4356095c30815e2a26;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8cbfbaa798912cbf29fbe663f5c9886eb301c80e7d478c2eb39ac91a3e4324d0c27d93cb29ca4a6ad426ddc0b943a95822d4af12a64e18ace44ad373b63f86ea382;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa1ab6afdec4ad266010e66eebc83c26eafd45718623dd247d518c449b2571ef5e7c9ac7d3588b49429b08951ccd16e47b9fee23e64a0e28878bb86e9894bf16e8e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h691a4202d3cb9bacb7d5d1621c5b728bbc26e03f46fb6575a4beb77b112b0b19f8fd31d86eb90a90b0f24d40509ac49382b0f1c1785ac99aea2fd1da925e8bfc1c15;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f68be700fd0d0934f0c56e29607487d0b7c3696efafd02e423a014a1077789ad8763b5f18fd93408d5cbbe6019e4a438c055b7ceece53af8a169d2bf09f60966474b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha54153b1451930c1b817642a6412e11fa1dbcb273eacf34985456639e328ba3d40e5921a8fe451b552a6202c42eb271043ac2dbaf766710dcfeb5ccd4ad442249e9f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73aeb95dce260f3fb4cc99686d4de5bcfdbec0fc3f33a7bf5f76585bdf140024d6d3745f05b97f26f524577ffe2db418b483e226797b1533725fbd1a5f870115e3eb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f80624445e651b5c7358dca2f986c48ccda34ec1c787b3fe1d30d265369821ed71e980728d8c3e113ddde29420f429b6b22c8a9bc3a1c5c5c9aca7e7545fb06719bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f7055679365a3a4f8e9d72aa5841f8fe6e98e539faa23eeacfac85b446b22272a209355c44111c2b04d753e561939001fddeebde74fdbf35d25c2ba092c728eecab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e18ac023ceaca4f2c7c645667e268d3d00b3c2969dc42e5e247e329bc87929f9abcd96e88a676d5e73b1f041fd9c0250a2dec2eee01ccf68f2e332038c2119aea50;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c261bc8bb2056a6b9092c5df8e5afcfde4fde139f43b0dadf3a9fd0471dfbead73c1d081701d87ecc7e3f91ca301d39658c3d5500ec4c6c8311262c0ae58a51c8c2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80fd32ddf221c65832fbd217328bbfb46d061c4e55c0820cef1f05b067a1abf8dde6d0b79790f74ddbc2f4f33d8eb0f14822118244b1af4d2c416309131879cd4510;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h30ca2fc1d8d6a8e9e5d538d77cee3d8775c9af22cb8e45307f8cb31c4832048e67719422940725740390759917667aa330d4b0488a946ca6fea50acd8512bf3c7316;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e204c6f7526d65f3dbdb8a00d5fafed74981543bd22af02a4fa456d279db4b6ab5d0a6bb455de52b3574df057699109abc7203b65e551b80b82f3742389e2d89d67;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f24bd11a855277e245102f00ff08d80c21098e42ede6bcee7663e54df61b82e19b79ff935bd172ac1d0056f094dbf493113ee58e927641a6d674d58a74211600860e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161b567ec2d9b5c16617681e41b05471e30b0d27d790cd0bea29c5da5908d6fa2a80392589c329eef0ec3f9242f2376b1b96d0036a07af0bf766a0f70391c1f85a2cb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd1906c10202fb0f7df61ccb6804fe281acd115d6a0bd0c5c5ad6cfa25ddadfcd905efa5a766b9ba696a9cc0418d0ec8d2447b7b7a63222441591c0d8e3cbcc72c32;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h171c30b4b67623fb862f6c50c7b6c630486a0eaafe0cfe21444e384de3b45e14137682dd557db4facbeb4b1377771675432b1b7475b9339144c4e2594a9d2e7f223fc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had0d87abb6669f6245c14eb69ec09106dda7bdcffb147fd194353d5f134503ec038e3df29484ea95e251edf9d7d97bf43905249b0df592136bb844bf026c63f39e34;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfebc629aa4fe3da5d1b7c0af80cc048da781b43551f3ac8f98ab123a125099cdea8321f5cfc47b828f4883bc5b1cbf51d97778ed8176e9e0b73e457c064cfc0c40f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f3e769b8ed8eb12e7ad03bb3cd0bdacfaeb0e007a54f497586e74b289745300c8d460cbd0a014f1874593ce3810afc18e30b88b2d1779f6f3e28fa01e4f024e76971;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdcc5ea80c5fff4904ac72ca53c247a1b2bf07c8b66a8366adc6e6d6d830a6d99e0d780870f6fc5dd423f98bb1ef2a301c17d3f64433734d84a43129a1e7ce3465b5b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h693bbb0b06411e04975db858ea0837c5fce7365bc281c223040ee84af19bd6d31c507a508f10ea7f0c0ba4df757037518dd30a042814cc9b71018f45cfec09192207;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37489d26c5e870358d31fe9a2371c9c4c4b0e67654c1fc15dadaa2484cc9990c6919008cdb6b42ce91921d38dcbdd6f983d67ef6ac56d2f2ca5e46bc7d0c54c3049c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6151ba2b6df308bde6550c82008f4c28b8ee66f3a1c48f89a34a957ea89646a76f929650c1f57d4709fe00dfb385172979ce0d9689cb6e61c1328753a4835a0ed06d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4bc552be6fa0a0634fa07ff6fb5ea3a4ea65aba291a112bbfea2cb51c3c8f407fc7c94059754d2e949949da9edd6bfe37143d0f1d1e121294edbd7007fb8eadc504e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ba7eaa0686750310465763dd1a5169c4336e701818326eb57f76da333e40fea2b3a9529df066e69601a783e0bf15ac03e3014b5c335787719d416458ce9fb5053cc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc1eeed347c3cd9a87c4ae74b4d30e70fde89d373cff550f3b93646031a9a15fb802d2f56ba1b3a479cc2da78aea1b5be71737895aac95f80fd5af5045980248512b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc4103cc4e03ec4d27b27a48a2a0af4b5daefa8e499b38567816ee317371f5a50bd73bd8cfc9a1a6a6504896d0ee831d467d4d70029123b3a6d54b075379d465ef196;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf96701e66c3bf66f3f7e85098b5d8ae5c1f4ebf57dc917bfa9faf5d0c420d32bf0ab3e6d3d2892e49b2236fa974ba2302d3727e12099a3b7185a5d26cf6b5ab667c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1af68eb64da05b0079101858feb9f9cdf3773064c0a2e52cc6a574d6f8a9824ab30511355c57c4a9703fdac24cc1b607d9bc73345e746912f98a57fc26a9e49d45a06;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b2036c785550a591a1c849916e7c11645be7aa39b96575d7ec4405aee0faa7595ba38f0ae3104516e80ccc11bd1a9679216a954974ecb2a0ebd82cc2ffb64f2ce92;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heef75a1f13696f895c2a7d23928241a95d4f3dbf1dcacb1ac28fbeff64bba464eaed3d4466ab7d8bb9175497ea2c4dcac8e185eb8e1b435677bdcb94d2a1c96c26b7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ffe84676d6af1b9215d859c3bb6ec4c9b4a3d20e2e5818b53b43228ec36a76f09a274cff95d0703e902cb9b38a177d1072644303cc2ec375e36c807c258adb32c25;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h143d2a6b66ac578b4cb224fd1148195ed1b7eed1e1af4a0f810b7e39da9a91e9ac15b232406ee513e7daf10db67f12aa13552f95da1c8378fabe67ae419bc98b6f52c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75cab481a88371b5b4a33dc3f8584e6e6cffcf71769ef7919596f055249151885acdab33116129c91232207f0515230a15375e734c362424c1bd4da3a6342e4d9b76;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6ff1831dfc743670a6adc76ee56a320f0402ee2791915343d4ba3784a4cb4ff89ab03a446bfc0182bd90063fa60e5055a1a1edfbacde43024dcf9d1e8f4f8f266af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf12a8f1850f27f5b94d2535d7514c9288613036e122fed0b0d85f062aefcf44a0b2cccafe6fcede424c4a92c7f092f0b8a56dbbc447a1f86e74812c5221804e126f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139b66cea142cc62efc9f3474a01098997432e218b8c7509b7fd074fa7ef7fd7ecf6b9816a4179eda5699038d90e670268af44e12a51127a15a460005a574cb709646;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa7f8fc84b23151895287a90769da2aebfe859d560f120f1302f2873bd6811125b02401030c3393a1edb132969e3dd8e035aedb1981de561792810093bfb1a7f6a41;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175410c91083e5eaefeec8d48060f09053c6f2a7656f401a66631c4b9d2b1dd4e487257a0bd6bc70dc6e094e925d4d90db99ef10d53dedfd53d92d4a15bf01cc91fd2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2562bb2f6dea429d4239e46f7a7d4a0a163569cb39099f0ff6bb9c3e02747e159403fdaf87253ebc2414aab5296c24d17809204f75b2d2894af2b08e6d573b0e7183;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf236eed2df3c486bd97c7ba98a164998be405df6148539405c90455a104355dee5f44c0783fc5a7a43fad6791c1dc6725e92462e612a3ceb01a6ddfd6cf2f0ad7827;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1620be85248eb878e28579f3b3e8f460ce0b08a073e5474f347164375289a6f8cb36403f936b9c51cecb98617c47751812c647826c3307bd0693bcc1759de19f0b88b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he43028d9c95f5980b33c6f448f51316c5f805268dc0d48ecf66299d0f8ea810ba99e9699a3071cff8a4132c1c08e9b5586afe0297c27bb0de5e88c632df2aedaa612;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b8a53d65c95291122a59cbf3354f89c87e82b9bf2bfbc457454add995d9cdb199bc474b19321a832fc827726be013dff23690db3e1cc32319a67bd71567deae3f8d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1afea6600ddaf2a8ba2f3ea8de632d8fa12b809a8db87173baab4b019a706adae6941a3300675dd233ee8f228ac2d40c39c361c3ea3e073e9faedf43e429e3e291f00;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1868875b43ced710d1946e7c66f31e31c8b1c54d3bb20d41370001148a87858ea51f1cb738a22ceae97cd1008587221d8a9cf2ccda3e3bdc4d38d49197ed43ddd2653;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h59533986b80f0979fb8cf29b836d953d68def9ff5162a6225661c06a359c0d63274e85336eac8904c36f453e163dd67772931a1cd21304af4b599f9fb6e4266908f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6a2d4acd385670d9d399b589265bac080420eb7629e1f6425dd81ce843f4e5a187ee08e70a711da8aa5c7a330ae9e68a64d4135db528f8ffc0bfdb867fa0e01fc84;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146c7fea23f413ccf48b023b31d50bb70a48605a7e6cc13e33d4a36d190ac143ef4a117257502fe0f47b6033dd68792e83058ea801da3f58b27292e5616f25bb5cf23;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164354ce3e4af48d3e151af3d1393680cf65f1c4ef85bf048b4bb8b4e4ec5c0c482963e07cacbe8add1b240364a0fd12d42b4539a9357cce54962834da0a6099f1931;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cc32406b5a4dadbcf265566391c9f97ae53ea996fcce9ed386cd37cc8739f54f538bbfa32baf653ec65b3072b7f4a26b76dee46c78c58073a866a437e7e21487f685;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbee330968122e4e907da08cd5563bce46e3d06ca24000908640ab9c5434f1895eafbf401e22a5cd69480441107d748fd8d15363d8fcc5fa77b33a32da1f7f86d2495;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6448431480c0b797718b86f6abebc90050f523f2603ef06055eb6b8fb40842df6d1748e25ef9e490a9f5e6636ecd6e2c792f925009fa01d2536cba969721cbe64e66;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3105ee5e6cb3799b8904ceecfd75d9f186952619d37a98b50b4c0546cc78f237bcff2676124805d6e953ff9d9b6413e751696d9f4b8d4a97fd00ef3983de667d7de6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce58ffd724a8c4a1b4bdc568cb68da5669325a661b997486d6b486eac05a051ed35141f7cb2d6b075d137670369490bace0530ff57c4fe26b5fa5ebedef64dd2f3b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89d7ee154588fc45b60e931e3d7db8ba40eea572a9b26e5277f92d326e4458bcfaa7f7c8c21ac1e445bd380b05969b0e0816105f340012c51051752ff630ee130be0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110c90d33694a372d6b1358662f86f4688590ce0b436ded44012e0bda6f5821b15da0654a5d3cb8d27f654391dace0d38274a3982b15fdc60a1852d767dbc87e714c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0da2465d1f56a78572e2cbf30e97b5d6280cc24c75ab21fe9d1dba3b965a7923f6b830b9e3831945936257a3b8187dba73837e39f1fec8486454600745b8dadd5b9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdfa2d6f7b625d21b39209647ac662a727e60444a0c7199923c9ebc9d74658c9ad80fe2fcd580784db4ecd336af3c46357567e4793b24ee3dd7ff041eb2a7779732a6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha4a31252b965ceaa0bd7067e6edaca6a4767726f4dbeee78bd4647dace27a203524f0ad69f97c02ddd7a411e399671f9d73af11537ab05a8a3ef861ed2e2f5091064;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h799356d333e738c73987a6089a718415395e02ce27c0a9806667ab89d4fd5c401d19c3fc6fda4a18eb26c2b7ddd5fbeabe97bd4f38eaf9936bc5b2ebaa18fead863f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha23984f17ff17d5f29713b78c482dc55a42c041f1026c2fdd9e914c6a04b9b7992768fe9da38090c771bba292a7d90973640fb8aae82f95f67eb7b8b54619d2c1f28;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1866092fae150070510789da9a662083903a3225770716cb7e9b299a895d7d82c691260c5deb833e59e7dcc814492dbf6619ec95fae2eeffc1ec27ed51857b65b825b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85819e3c383c35f6f7fda29322723dd6eb4e03b242f6c0711cfc1c8066fd076e37d0db957d7eb0a3306b7026bbb059ae2ac59eb46c272bb4b27a2c3b114407cbf251;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4d90a47c1712bd9f93c162439f1e060dabd5f1fce44ae5eed9b3a9caa71cdda038f29209935574a3b5f2e920d16efe764727a273868eb77eea27b88e5e9c33440e5d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he245c7da1399f188ac6267dc62d8812a09c5fdf342053c423a5a80da5f6127fe1de06424d39fd4278de39470425f1d53dcbff213cbcdcd952b491b3d9316864020a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc2c5d0069e6234718ff7f2f6187903d8b49b485611cb2e2cc0d35efb641e02d6f0f6f3036cfb3a737ef811f3b28136d79320ce2ce01307505aeacb0ca49f56ef5a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1688cbe14afe51d1927e693fe5af2f47e7d354b333b0f47fae561aa8e5c4e243a84d6c66e15a76ae5f9dddb14f7219bbc8b38199f0d22f8f3bcad75fa2af3481b36ca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49ce3cb6fe26064b283e1b8c7de2bdc1b90c987e0c5cb6f1897a1c97c6de5372e0840898585af2e710f4043847682d92f2e2d9d5521af0a27d42e554d18f9a4000dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1383efd7a99ef9b2a6d932c16159b1926672103cedf595a424a9d085c1e40382c862d5edc452675eb50ffda8972a46451a319972971de10c10b45874cc7a1411cd275;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee7f5dddaf7fde059ff2e11471a26b6a47761a23a449bd934a16d9ca2f998a5920477964677a5062d5ebc5edb560c6291225652c81740329ab29c78b9cbab13676d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47c78dbbd908eabc11699bb0f7d5a6a41b2b2c5b4460993bac09c023798cf88540d8cf754ffda80a130419d55abaa0b50b547d291876e134aac63b77b5cf3590a40e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1715aed857cab9bd8d0cd9e3a1e524e11bc4a24fa4e1ede81afee2575eb83be131e507f96a2d5a1b83364f7a49164366d7292400bf74b070d83b5bc2af2ffb8f37f0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c9f5bf8e2a48dff3a7ee1e1659adabdea5c3e438ce23900dddd566b7ee9efda913e44b6c8512d64a9230e0c7a596b49fee0929eea85811ff18db57455b6e62faa5c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fde002088d58c1e96a35a412bf82938b18d0e516baa928fa274aa04a1dbc0df470d6cde263cf1f1f951ef6cc6c006100dcfdbaf3bbd0b3ed798828f75f77e519eb7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h177b6528a80648ea24d0de5d9e1490a5883ed94d7ae429981544162bd552ae276c94d8864621f90cfcebf3b6c9e0050d6de649bb31fc066c9788a11e58a1a76cb0694;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11c922711bbb3c8567b336a57b2f7a30aa556598b2448988a7f209034144fba0c7c4738d27d6b2cf5f1851a966766951028d5f52045b81340bbd753b23208658d2027;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1749439db47abcd82619e83cedf0bb3db51ddba122f4b6182afa484334d659bf0bc70235a4f76e455d823bf179674eb5ebfe21e886c4f4154a4d4e9f6851881bf6795;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b17427b5b8108527a1eed34693e0ce2fb590cc1dcc1b171a3f228390174047e1c1f5756ce3b096d78357eeaa86f3dfac6f3c48a72c33f077b0a05664de2ef94fcf8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6dcdc772af9bcc959fa9972f40c6b1e7e4addf2996cd7b9a0ded8add860b80d3fd7560849834e5f807c5936765d34ed84fd816a06a9d7d0be1c3890dd24e1817c584;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3d39f9b8f13bfd55ba4c20932113fda97c837d943aa2f28506adec6c6694c3ff32960a867630780c4acf51b3ac3ea81fa56dec03674a763470d994f7e39671ffb3b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5fa9f57b83f33a4031393ac0394dbf04d5f1032897640cc05c048b8bb865e0e3b2a558a828d91f29efa794b147d5875af00b43516025417b772eaca74c50d5f6602f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1468f8d881a38ae61b5e57dd1cc0145f8009aeba79b7ad2bf1249a7cc37f4bc071b5f2dfadc4d00a495c8339a49cfca8d4226bb156881fa6b53aa88898f32c91d8db0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10bd0bb978a108ff7b529fb7cd0aba85bf83d0e743f8a7ee248cdf1f5a64ab800bc632755ef0107e1c7dceead49d5fb6675e913515b543e14326141d8f468b4e652e8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf8d34bc5c6d862b71ba9eb9ceb4e5a9896856f27a5f88e0df7a86f23720372813b31123c795dad7300663ee760c24ff64e3341f978e016fef015c0b08210d4ae4bef;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6025f59900e2d55da7fbfa1c162477dfcd2e36ee16fb12df262602d3f6299ee049ccb45ea8c7cf8cde8d6f25ff4beb90dbe1d0abccae889ffaacfdce465fc6f3daa3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a459804280772c7e607f3670af70fecdae24d711b5406069c2cb273598c79811aad9df3a113f28d1af9ad8599d89362c9fcef20d0edd93343d8cc607e84c3f328709;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1befd69e2dc77e2079de2d7a2c66323c0855032b96f733f6e51097d9d7e33981163dadb510be81f9a8da89a817a8783d5278b1b57b540857c60a63b40f72dcdd9cf8f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6f255c94a612a345399b99b0f694f93ce16892a60f5d609462bc2b6d60c7f9df09e6211cf1683f92b7122f1e4ddc206e34d52a805555d6e2e0d4bf9be846052e8a9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c874aa03011e89d307f58be42265a3a827b64d7073ba5d320166797385e910f60a93b11fd26ea8c8be7afa53929f2bcc8e822b907db6fc50cdb33df8eb49fcfca81;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h443ca801de39b5337c0a787300baea3567f235c39d7264b4c6051a24b160baac0cd1a34ede32c050e302af792447554c652be440f802e43a9159ff2977d797454726;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h64a98439d4d217934ca2a61f74fe3b134deb36c53b6ab6c2f6c7376046d370bd2eda2a53662d1483c1ea942ff37ec518bcb0c2887a384b6fc19a94c699ae8bd92a84;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfc1a9ec83c485886321f9e8510e098c3ec41e64757af8412b9185c9cf283c40fea8e669482d82b33af6c3cfe4f2d063e35e751473c567526afb00cf778d76661af4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd538cfe0b5635955366e8aa960d17f2b916a9d766977d8f11d3d2ee0722991f31da4f51257052534f25491647774170019e407d46f10f93e408dc8bbce259315b489;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e7328c51d6f6a88582afff4063dd4567bfb26fdb32ea05ab41232b6fcd6c6fc846f8c3e193f764fe1360dbd74c66b16dbdf55224cbc5855dde9671ea6d58f377f99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdebbeff8edd1e5026fa5d893157893512e7aa37f711e18eca7fea827f1b68f048747b982be15644d9b5d005e62de1e2af398a86ee427ae925df9af10143d3b0e9b1b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d106eb41fe6965c6f5c57bfc2608b06579afffd84ca560cba58b5bcd8f23eee5c66576d92b80aa9f8a1f52e72ab6d7b9f3eb109535fa304b96bb17ce0c7182046c4d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd60e2a3369a0c67ed2c1d9437292892aa9052a4d40e04aa46d05230a34fef9ce540ce04364b3ed3de7305ba2e68df7a0c708e184001903b0184881ba1fc3557c6d1b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110f26b12789005542f4f21f3a0893930724af6a2ea1eb1ea4da25e7b8d8de6a61c9c0d3809e727a747cfac7187682c75843a75f6404f4ec6439782cabcf3b226183c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb98b4fa6e8777ec5eec6a5dd40493fe54809bb2e9ae406400344455f025743e39085b4facc33332009d321a7cac9b5ddeaae7f4adeedf4fe746cb13d290bfbaee60;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e23f3748c0469160b8231e7be44bea90ffa22ba2ec566e30fe32bd75268f6b05a3985d228ee9613b179ecad1f010348fbd2f4c7456b79df98394bf45231a8c342670;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1675aadc3c087424c2f80d0127b9e286ab8adbe29fb53161ec660f3d90f30440be2ac05a0b215d8854f1d7de7ee062fd5ddf0f8aa87e3632ef8103f9d3419a336489e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea4678979ea9ecdda8f83c0e4533fcff8549690a98cd636bdca93a3df36f3487f45a6c4b2b096ad9ecfecc63d1fe24199801f4a12c7fc9c5a7821053c0dd37019af7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h136e746a8e4bcd39cd935870323e7666fe9db07a63e1e1575a2ecae9b214fae7fd40550b79ffed97029aaf0428ae8c89448d306cd93ca6b853e6e9f90273789acc20c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h760700322cce879fdb5b19f0bdafd8362be5905009b13199f9052deb6e028eda5207832669e5ae74a3bf01b7f8193d0b985f0cca2573dcb9afa008a1437c97043958;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1c9dfdd7e12fa1536392348948d1cf5eaf761c093c2173cac48339ba6d49a6accad4757936a42db3c066b1d8bf5022682f005f60dd00a35b3eeb59bbc5d3f4842b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d627b2cb1b8a9ded8ee1aeb05de555a833a3d0f41822d2c2d9470589e866307f196ac672b0b3d3a087c7f2fe6a3a4718889390210f95eb2e0d2d1ab34d96f5e0ce05;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ae2d6293771f5822c14c086d230e12705b8a51169593eefc4ae2cf67b7fa28058f67e5164dbe46e85e33befd964b37410dd7fa3f88352937c8d01439f56083d20b6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118124a018d39f0b3572370662681de8b78ba6e8726652966df806068980a18608228d11d8beeaf354717559ed67333f451d779fb4ba7258503a11055ae16076d9c56;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10341033a4f8c48368ba92bf3268011fe3dc7cdcbec9b49cc27e0ea9840baae53b72edde0b26ce10c7844fd5c1bfb8cd2770f6d6a28609caaff35cc3ebdc797db2636;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9b9d3eb6f43100bc0ef5675df3eff2eba2025402da0a9a0676244058d98dc4cb227851c5cf9afe5ce79bf3205f5de361163c371a64e4f4522324a4b7d0874a3f61c8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8662a489bdb3b48e5284f48088d81775762b5bf24e4080d5723509186f14dfd66faa8a2eec4d4f4e5bcb5ea57fd1ee74615c9fd3af27a42fa6acb9ec351de47d739;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da343dd6891b82df22825812c77c6b227fb8f35410a64e96e3ece7977ead882b4e285e235e3f0f51783198116bb396bd261d1e6c1f121c6c9d0cda6c53d7d4907a7e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3abb9b006c29f1842339ff3e86ceba643a45ff67718eebd5862a6ba66a4a6b1d09a98c94d1c89dc8eadeccd1afad04cb07fe589f417bc973dda56507ade11b07cd0f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1388e504a2b7e6708500d8d038306a5e5eaa157f91c700addcf22b34924bdc859641ab1a7a31ab88ceab8dface72d16ea089f8ddc25d9088c661c873d2d05dfcb2323;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he2b4637c3db336f02640c4ced9ee9704144eb3a2a68a56ab016bdd9aa6d28907cd1794fe4e7460515f3465270730cf4b2a46ebab6519ae4cda5970258320e23a3498;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b41e687bf432b7b1192ea07c62e27c83c59f7619351635aaafb6ee9371de3a6cf9e9ee81f36271303a64757813f0e409240bab64156abfcfcd133d4488f0f29df62;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc15d1e7eb9cf2018c38539a6f19d41ade1272303d277a8df414c4a58dc9c743d20acdb5b227951a9783312c44946272bcc77265df243ac289dd6d2a45c3641c74600;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4529fd452b71d30b49baaa1578103184e82a99cfee89d2d1afd733829556215bf5d727fe31a3ca905dcf4aa72ad464164bdbb95551bc6c92b1e439b62bb93404174;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2400aa9b3ea7bcd7946bfbe72529ea892b38e8d0a7969252f906937a74510e14f9097ea1225a4210eb4c5d1b3b14bd2092c1050fbcade3014bcfd34507cb23859ed;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e96dbcb730195ad6e7c4d90f85e8026a327fd82d52547a89cb825bbe18d2a9fad83fbfa08044ff15e4c17d01b80ce03a871b04cdcdc5b8944993b589ce6c8efaf83;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e1ec44de6a1d74e580c38bbca6e4c923bd846952ecbda1487cef6b07df02c2f0d69d39d9fba59c154b15b8cd78a781728b0b9103ace932e35d6567a8aa79b82be6f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129a8ac14e398b403942e596ba0f4c6c02a27c546e790062a116197faacb7ef7e2e33039dcd903e6c321556dc2d8f99f1dbbfd02ca94f3d17d3babba9e42eaaf0f41;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11edf872ab2a79b2dd70bb0b4ed14792025f4ccaec9fc65db5a00fc7e9d5ec279680a416921d5e79566dfa50274f89f08d8e4cfbc76f0b5460085b814f40b47bd7770;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf58849e8c2704293733be890b2dfa6e3cbe248f6c2d6de0e0cbd2f4caf79db5e3af163cd38a90f2d1b05180ac48d68219e1e71872a4c7c90bceea4fdaabff4cf899f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f20666d96be18c0b16b890f9485a532db7ccb1234440fbddf8218a5a6c4bccea7d4662d54e7b244ecdde3aabf91947caf5b53fca337ca60d7bef23383f45c0c351a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce3a30a3a6d0a3dc6e538a4b1108a8056685c05d5cc7e661851a0bd6efef2af9789c53225978e9db3989fbeb541148f7e49dc7347c1f5981de4c1d2a9a8378884c4a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he74865edf0e265192821066e4a85fcff9d08b3f1156d393b9391e900ef341b4d88c2645e1a4d7ff1b5855915b60bf5b36c917b6617a8ba4481246fe722a7f12c061d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a92fad7cf5f8444cc94edebbf8735c10c21788a0015fb1339b863a86511a433d8ec5f7860f6a9cb9ab289957aa5b7676f13bd4caa634a0ac602d86d0dab6faf0851;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f30eb9df260a915051b53f53edf4bfe3920f343a3328c2168d52d2f814b60938f5007390820088f11fa920d4d04b797857094bef8537921b5f8da08074f7e2cb8a72;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f5a9cdc198472dbcf17e1d01dbb6841a5041ebe085af85dc0e5daed759cee045fec91b10a902958fb8a806e3b3a6785e135c397d83c98bdef39e8348813103d04cf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4d86458488676c3ff7582b84b3c4d1ad9dedc7b8c5a62279db524767e5cae49037d8477fc3eb4c1b2f791fea6373ec85b71292130ada5c26eab553d0cdd03f274cab;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h882f1eebd64ab63e6cc22fa67ff9a0c1219454df9b675015e37ebc14fc28dc59428d6ed2e7534d6b18356515547c0951a31354284aa3f2d1e393f1727ae41d6ae5c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14921023ce913597726384d4ea7d790d065b95c8b7138442301d5abfd48600913c12b1ca50d342bd59304e5f5d77ee5081a69417b1df2ba5673547ae5d094cbd500d0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h298ad368b4ee702b043fc2fc3974729c03f5b5bce5d7f4add532eb409158a33c20e91a2a1fe4a9bcbe894a68f1b2cbf9ab31db0e9837facfa69f05274b7155256420;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha164ea9e7a0805a4b15fb8a82b6e3ccce79d7a3d9acc57ec763f12add8686f8d1ff9867aa751d9545bd92a47c43537fcebe34d5102ea6b636cfb10a6bfde5a76141a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h700c53082b955a2c4b40e7ac31d00e7d205f9b7e3dd11872a183baa29455973d25374e1ebe82d9ae257a8f36f0bbda150817175f7aefe7326c7312b6164c656b0016;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14bc674e879c33bd84556798fc033bbe6833ddfa298034a81cd36aa9b35caae577b4d2077e21d3c3c564a6007e9c52ca613d44f9c510d60bce4e30bf0f3871cb54f33;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h547d5a57ccb76fe5af009f6101a1acbcc5dc31ecf635a08e141d8cc1401b0019bc94c657228edee05df13033192f27d5e0dbaf7954aa5c9ef92c05daa08b5fee91a3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0a9e1497abbf8311d096580aaac34d8a5590db3218a390860204855791c13c2e6446c03d504e35b76d2c3d5465ac29ba8b5c20bc7fa1e01745dd0c62938a1e61243;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc02f582f8d4840bf55df971c806fcc0a55026da5a03af1ab72f4179b959467e8f0c153d2e4b49d9786a981b820d6d2ba4e16bd68d33bc9bdc9a3b26b0be1f75532c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4865d616dc148dd44ffca1cb07ebe4cf8ac5e2e41f015ed0b645469babb0a0d8aab8639b87cb9bcdb4b75ac2c2f661eabb69089571fa78e65e582e369d0dc4248a69;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1abc1673932c5c1e90ecba44a32662652f78bb7217e9788dfb1a12318069a54b83b3aeb37abba023ae6d05b5c1fbd6d3a706f01444f23d35cc40ffdae860d4a752f08;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170c020d0137c25406a5537fd7f1cac32e7409ab11b5e0fb20e705aba0e0456ca2e895a67696871fe653d8432a19254220e0c871effffadc44728384420ec891ebf71;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ed71befc88d1f9cfd52cd94496af9438e9babaa0622aa590423c275a3abe324762f4eeb4a55b419d7df89faad21a905662e38ba9004e02e07723222162f0c061465;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be6dfda44fe55e3cc7a74b62769b6b0a0e4153e2f973a9d02d1ee1d2b25fd9c561ac38a580f6569a6eb7d5847e7a38f24a2e3c615785b4b00bc33e9728dba882f38;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b56c2173cbd638595eec70c86e91743c1d57738bd7221b43bf84da4715b9f5c725296d3db22fece65ddf0d97f9c0737ff2e32a1eecd5dcc2a5b270f7cc85c74d6b10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138d722e5ef0e113b7c0f75710eea920b896e22139849231ff479406efd2bcec69835c7f83fbf02ac3ed32bae9bcc9f028e92ed0642518736697d00a5fbcf6e556eca;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7bf13bd524de338200a0cf1115226cd87a19482625987bafdf4ac14fbc177fabc7b9b6d7da9971ce9efbf6babc24da7b091d25ea90dc7c552b276590ee4135d0efce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1019fc2066257ebb7e091c718b9c9f14129b7d14c0a015dead12d218e60ae57dea903456f510f8ba5f3ac076ab459a87ee7d1a1eb115c9241766a8aac91f73f334a95;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16d323f0480f5cf5e11108eacf46ba82057f1356447ae4512db8a1de775d387c337ddbab0c01c8e8941faf0d4de41587b3e7d5b3e0faa3e9637baa3ebeeb85bb6aaec;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1361e58fe7b7f5db2eba3f5d5523f02606b53bcbfc987e3eab435ac73a7fe1f6f6dd96c1a9b23135f5f075ac2a8dc1ac75815cb4d03efb53712d0bd718f4a88677961;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f52686a4af7c302a27c90a82b0c60d382ce34d4e55ef1e3058aaad305ad148b6a673076084a9f561cace586ee9faca531196c68637323b710fa766b9ba5e9d76961;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc1b236cd9e9b39b3dddd7b8f9a7f5f4b6d797d74013f8a9e33ce4346c6e10b2a2dd0a3f0fac0091d42f1fe4227e2d34c913f9fc0cd944ba2fbbcd5f7dc61d954d42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ae259dea0a57c25c6195b0dc5b1865b10d1ff713e70c5a71cccb1a6a145ce6db8941dc1d1f54c86cfb391c5823f7f44deda3ea634016c19b30f6699125fec5fbb10;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h75814160256b868ec0d3bd7ab850337131eb4a90513b26609a193c48d596a1836d7d70a22ef85751564971fa797c1d043462fca589403d8ca451bf565697e8f9be74;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb20828148689dde54679e1ac88acfc3e7a6afe52449bbea055b367d9a39c7553918279c14baf6aa2b35673cd9dcac5227a6b492e1bf6a04f4431af155cd8b857e767;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1323bbcf328587a933cd6c73f6200844c469bbb37a1de4ff2ae6fc11bb614a4d2668c759fb994c359f86c707a7011215b505342746a18d0a623ae497fa53c2b79f538;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e17d542240f5431c58946253b235e73bde4cb2556f0878b1e821465ae97ad123423bff387df5f929ce3f5cbfd6da81be45b963de3c54b56321b0150fdb749d1087bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34d41dc294facba74c70d1e9eec05f3ef85fe355de8ec8c955d5cb4b2425faaaffa8e31bc5561734f3837d678abc7bb051ccbf8e99316dd20fa442b7312b7c8278f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ed10318b29167e7a716f12ccc29c0fed926ab3e7fa81c5d66a2a5389ec097b1f85e71907a4d2cee07de06cf94f2efbd45b9bd0ef3c161508aa6851f8c21e5574187;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb48eb76486e25e8413c3f794c1a4b55dc9db86f4ac22f4a6f2a195c62f6a1e31fea41268dc018eed8558b9f63955833eb185bf0951f472a4e28e847d2a817e7e69f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87f918ec78184c037cc5e6f5ba966cc3771c4df66b5ca516ccaa74727a6fb0c40e2196609f2be801eb3795d3fb6ac809b0cff86f4220d0b1ee2061d1f6024b6ffbb4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d7fe8a641d022f2dcfce81fefc757af969c9a524b30cfb123e1d6face0e94db1ab933f1b8fe7040d30a57d2bc097289a7399cbb2df36acf775f98315afef3fc379c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e2b969c213f1245c904b6c0451cb739ea4dcf53f42da7a1450df6c1e4bfdb1060828ba54c137d5c91a83fd8636bd3b240c24b91a05e5e2df1575738d75602d18b8d5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc16ecc79438fb0f2aa05188d2991ab42b9d2542aca7d4f95b617394f03374c53ad88080cd2520446a68b8d23b60a6f1224decd68b14f664e8ae46d645b14c30df137;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5a3799e32d5ae1748936d0a68c5dc595a5934e9e64041a3dad7ad844b4276b9bbeb17edaba552b336c418f9ab8ad9664346a9ed842b21bb2030d139f246c285f4d9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10830cb15fa7752297117b231b3f881dd4609fd0ccc34adbc58da87a1ffa6470ec67a0dd15d48e3af066921e806774c65ee74f918a137466063d02e7e8bc20c2a21d3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2eee3202bba002371726a1e0c6953d48ab66d3f689b8b8162c4743c29b6645e57d6f2fb2739aae8afa7096a65a6d415d65bbab2aaad69a627ebe6c19fc4a84352fb0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a20b5a240b9026e74bd993ba80a83974f6db2cfe340d7d4281260d81492117d97f63cdb0be12f9b9db726426c0f7e460cc4eebda9313b69ef5ebda943ef07ff359f4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eae50c0d4c4c795a1b6a8877d32a49f49b3325ab215076cea97a503264b4b213f3cf3d9a28cb873cf28cc4c860edc93e7c863392fe2111d11756d441818c18f8df2f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he43e32e33c2e781193ead0e7d0a309459e829a75b7f0c583a522f7c72eee4ced2b633a15b6daa607ba145e45678c92b860ddd2b918d70a365284f3bf2ba2b5a3a21f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha93035e0521d8cb9d2326471dd1e4e6b246a8f547e9ea12e0f70abf283c80e988cf668fecdff93009fa92726e775832ccda7cc2dce06329f1c999955e1379aa09682;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a84fe82607c6098413ed1e47b9c23a2fd05a80cf8d7170690b1260e571664aa6d1b7d6f106c441d3b79b1436df0f04ad71204a93f1a1f6c46fac5341a3020d15971;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17e91de9f04fc104ead9082a069b2598d93ee4f2f6aa0592d5a037dba7949ae819a084d52eb5a8ba3570f8a9eb67ffa1980fbc9efbbe92fbc29141f6fc9a89f78ff51;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1908f75baca2979e7214cf27dd30335c7f0e36496a5cc53f2b0f9ea6f291bb63c7b837a3c6d449ab47bc5824257a61856ee993af21b8e0a545057754a4bfad92dcc8d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd8f49947e5d5ab3b47a7fb7707e75437fe3e8608df8ca0a9ab2a12a9d6721160ffbd51eb314275f854ba4d6419f2291428e623dbd709716df897786224513c934dc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h760a8a59f44ccde0709e4209d86628a41f978d54669464fbb867a109d4428f78f4a5938922870f5bfc00388c1adf47a2826e4ce28f0f91acc7db1f8e768c83a13915;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cdcd14d491fc510ac3b63e3eabc646d538f5b1d192c431322884ce4add244f69e69397d6fe09f4f598f56408b139cae346898447a1acb307e50a2af56fa688518977;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17eac39791d3613eb0e538a61174655bf347b41b5623362759a3acade425aa1265d20c1863b0aae8f818905dcd83cd15fbe8b5ecf74d19b33b662a8b4828625aa7532;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc0d2ae9ccfefa4051e439731375d651a015bdd5489335b41483d1a24aadb206b9c2b87c07b7982440aac8c81796a6560fa29ceaeca5e212330014ce36b62a1ae5ba;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118755204468fdecf88e502e87062eaeba48aeed95d91685b70cfe27e82fb5bd92b36708101383ea9b6e7ab8bde49f0fb368f95656c6300edcd2aba389da029980d2c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c4933d505979a83ef9bf14b3574383d8c8a2c212db366ad6c13efd624cf4d0d0491ea4df5a87d25e45ef1fcaeec7a52a268deddabd8cae0adc073aae25ab296e5aa4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9fab659e32e2383d929ae5e1b2c79a5f3fbee4fa28d52a0139acfca83c28a0b1d1852f54a9957a4fe1a586fcacbbf728bef24b963d93b2a02837b7c8275823c39ce;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b8858cf4a105977fbe9b41549b10c3aa8862b7340fd50fa8ed2ad103b76e8a2333a3f5962ed6b9201d4c725a8f19117bb9dc0312ea7f3d30493ea8a328f5b261ab4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f114352fd241d5bad0de3e489a1082f86e4d17796132dbbfc528ff79f8ae790a0130c6f9153fc83b8275a39871b7804a4eb958f8f95f0572ea9c097fe7ba41630a2a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133a3bfe53a55d691e59e58fff2ce432f112074a7de734b4803ac59303305d74a9d0028611c8b3d64e6b8aa5789e811e200a1cf7698c39f79b7d294929ca72a247442;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108e6be7a75037af73646f92cfa18e43f716225e14cb378abd56b2d697952a62a9fa2115979a61f2c965c5afb27ef84f7c688895b4cc2c1fd03ac838e9ec7a987a7af;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12df30ff9722a70938b989d85e7749170b2be18a548f930bd5f785c768b74f0744f7a32e0363ce4fb1890a7903bd23ef02fd51d54e88d4954679585fa3adc736ac62f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbfd0dab2349e8a3c3af952df7a0aeeedf882a2fb13c2d83c91a75ab06aef8c708483b63848b9fc018adc331efe573a25862651f147657398e412f2964b7a0857e8b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcfb236f95ff0b0bd66b5d34767482c6aee590780b0b716c090b1335f3ccec7e7807529b5e875f674076a14b85397dd7f77ca07192d3584fdb041f52fea0dddcc8137;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8fb1949d4dc96bf99cd35df6c32928e267da6b17c723a02bd60bf892efa5cb202d3c90246ba3879c629a483f39309b1e9bf44bc3e290257435cc0c1635b8ec014062;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73543a42c0b6c288d6d1a397ca44cd227145536cf38611e069a4f9783d7d5449eba1166fad8e9001fc5bbffe554eb587eef44e4e972d9cd07500563728c7d0b91eae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6eef91f679969015f2f824935fa87d8d0d3b9e3e00e48d8cb990c0d3738a73f14b8509c16eadadd531cdeb0852f33908a0d86a45156b20e547724a07a8f52564feee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha7d434bb26c676e9e48a4a7ae9fe037ee9e5963d4b1c0910624fa88690d92617c674b051d993ce89118f7455f08b153384c60e05f34505109e23123c5d1888b6ca2b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d2b6bece8fca4693aeac1cd0d55dc101dee5e4969679258fe3587270ad470dc48a6d5c1e7fcc71b67faac37ae6002a932c079192494bea2d880ef1646ccbdc54c42b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1070c5cf798f24d25801cb5d962b678c4cc2a98a3d36dccbedc3cf87d8d8d5454223212496c9ca0e99de53d5c0140188517df030f9df1040ec0d5853917ce3cb5fb52;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e62ddcdb8d167ce525c6f331c58ec66890a98c0b03440a69095c9e48a2d739fdbebe0b03ae1dcb406e15f540dc2a71a643e82874c934f9ce7daf25edc9aa902f719;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5bc6c106b2ca5c69a6a2fac0f7dac80b5653c5d1d1ed10035e3a8b0cab67208b7acfe58b8e73585a21b4de26d8ec65d3a03b0d3a4f4dab3263461753c5b8f715f2ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc1a6456021db2e1c9246c3728501d91d1efe665d81842e057ccc3fa3722fe481e88d7eb8e429fd8211607cc6b2ff185fc5f63a03919eec64dae4f4a3326f44e79240;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cccc999b27726cfa8613e2f4bd803f5f00ac1451d3f42ced46102b1f7432301322fad9733409eab74c2e18bcaa620b53f4029aa1e7afd98329dd133b50643ec51fc3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198affd18c2aa1a368328a526dae71021a3a795ee67783d46c5e57756ca7035b96266c3f94b917dfed546ae30100d72c814e8ad84fe98f70c69da12caad5effe8a112;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h39eec80588a5ea976a951bc72e5c45b1988045de61f2ed64ab4b94972419079feb0013b584e7df8df1fadad235baa57bbeeaa8042eab69caec4793c7837e2dbd4697;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef39a4a8fb4f161cf08341814aeec359fbba058700fbedec10589898b27f1fa972167265d1b4de85559d3b948824dbfee35e3bd28c185ceac35acd148dd456348f3f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hededa7fca25e43d4fede570951f57896db742985c304e651982f0a3c559c3ffc8b0c35240c622da9a8d495639a4963b80b53263c6ce4b88541e9a64c0ea3fbf6edb0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15a8701897e0f965fcfd3b3ad347fa6cceaf9486dfeca23496db1d6b9c75ef55c5d671323334a74329c142c328e147a77729d908fda9a53ea43e6c1263c58db8f3816;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c96ca6e7e37efdd207003e718a432116c19e571a5694dc380e5cebafc2356ea70b6f5145a59f8f8f6dd85e938380bed261be3934f1371db1376bac02bea1dd9e84b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14f7c6873199d9f38c79a82e0e2fcbc4966cb89ba0a5ba251d67bb3ac6313c946f22f6494153439658e2606edff6598eec629288e56bb2ad2cfa3e6d76bf546e055ff;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h186aea2f6e20fe6844952298aebe1d65f749a0b9617f41d88b509d8d52c02c1eae2dfa0d46037f2fd8053b7077a4aee0fa315735b47bf871745ff8d5fe83cfcdea9bf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37d669f6e5d247998aa763be536bd705d7f11d95b97c18765dff97031657c4617fc3f55f8c10eab42db6502e5d2a2b2f2f4bafdd656ad434c69f9c4072be962682f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h609023f647f3fdb4e4594fedcbdc235c9a7beba66cfac17c4f0806be47f986a7cc9772d5ab5099fa574411de1892879e2381d84b286903b895492195c7a2f37837ae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc456906726a299fb1aa468b2565fc255f0682ccbd6b956c8ce0dd5ca592249e14f6826e7dfe4e8b360cf8ef75ac003a771e0e56261394337156cbf11a7927d1ff80;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed57ae3cbdb9c94875d1eb18c50268b13b1144a63aee70e2ed5cf31fd2b30bde054ceaccdeab77196b8a30a85eb2cb63f595be9cdae715483f93fed706063b1799ee;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h142ccccb5a6f95fe09edebf834600e4f131138a3854547a159f29ea609b1fe6a0b6959120deb63a16d1040ef95f3a91cc3dc60b97a4c2c5d9d2387c692a2d4739c5dd;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f6c9c135dd9f6c1ae568f858c934b674fcba1e3abc5ce02c511c6984c19153f6a584795b3163d5df9dee774364f652ec86f243f4836992c509ea3098febe55c19d4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12faaf9ee462f4b2ed79e948d845fa1aec09519d884a96df42a4285ffd7da618ce67c51b41b186287c25bf4ca2cd98bc3e53ae085c81737f1f519d420a40f3c593ed2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13161d50623d99acd80ba7acb86a90a600ba7fc6eb9c81b4faa607838541474b8e015c247d6afbb142000442dee91b0e15254c54e742da305969735a7f7518c8f5314;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79063ef04ded04ad766e2ea7e1ed91936a4b55e07d4db8c447196ddfb920d13d478fbb2ad65a18334a04c8725e5cd2155e868e570dd3b94a772ee6be2e36f1548447;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a77977b4a37f4ce029285b4967e1b9cf201f6b795366ece7cae4d6318df962673d463d8a7487d1e8c549680598397fafd1ef450c2f776c153ac6841a025a78a73f54;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c4c8267dde543cf0a2295a683f99a5e66102e9f0376fae9406c7d9a9c3385af1b1026eb86f35b11fced93168b56e37e0732a33d0ffdef2361a1ebe06da5501d615c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc5d7f1409386638976daef2a349660a922fced6c2f175652519b00bf7f37de17840a4dac92fed961e219fd558b02455eda6ec36d73faf48caa9a1297e10a73e2c57;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f671d3decbf254d988a07faa286089818574fdcbc161e0912db6a213da326bda2ba57e1ae32b48461f2dba265ad59db5d2559d3a6b5818da103c05057070c10a318f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60a85840114d9e4d57322968a6fea5abb1a5b309aaba290f5dd2dc1fcda9ddfa392bfe021e640070294481a544c67402a60399c6c716871f31d516c779e333620189;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c7878de4120381b5e5fcbae76fc54a797f2eee2ecbe0efd2cd93d267419481cee314728b016231c68103417b23de2828d8cfcf2e0b089fe39a3d6be11d75d2bc0b0c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137135260b4a17a182c25ead70ba3f22355ecf188940337632ee3b752a1d620539b5fedacfb6e4b5cf895a2b1fb13b1fd73b312003889d4e626d2cc3d872caf78c41b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1873934afa95852d40f6d5fa4fd6378af2e490260a18b3b0af0936173ad6fca4235afc88fd8d87cffe3e275e4cb0078adeb5dd29db98a6acd0a9d824b9b5d0b25130d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d387ab16a3e3979faf094bdba5cf558b1850e14a6ab92ea47b362352ea0fccd124b87da1b8bf50b8dd4880328973e9cab18b896c73b6bdd1aa8dec101b94fb1678c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h805b3da9491a01fb5629c857f9417adf82eead0e6a1bbbecb961a0259f851a00d2e06b31656ceba23af87ac6beef38135123a3e18bb4e6c06efe7efb563ce0e5f009;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a26dac1e05343c7f38539b34180429057af65137bedca8eaeb26b93e107798915adbd6c2b1d089420492e9955e3bc15c600f48201e2270381f08669014a46a8b31b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hff1f81f4e73e5ee8e41ee5e1c35d903f56be9c5eb54b6582b4714469c6dbfbe6595c64a66ef829dfcd8170c56bca54b3dd73aba499f62249cc4a21b6563b17ab600;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13994b93597ba396ad388562e959588021034ca44377b76e4aff980172256e2eae5b75084ecee381cb9fcb5cdcafefde14d67e857b1c748d94237b9914b01bd5a60b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h52dca10bbe5c000ccdf6649a48ac698974efbd974af3a5a7b8410631c863fe5365c9429895d4fe518f3aefa9d451cf3d3bc29e9f174307d2b4597b87d2cd4f1a4c21;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d269111ad57e1058da4789db05377c54e5ace352e17f59c02ba861e6c09349f030eb484408d282f30261c8d3542971b41510942e8321fc238e31c85fc7cea62d214c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83278c6e40022f72b7f9792a531b8ed147f79187118c5a461c123933ab03257b0e4bde49c940b0be77bb0e0612551196f61a0b99d78aac3a090132e6ab40fe21f0e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h40c46a07a3a7a7efbe02fc1b36aa7db104521b8f7e16de5c5bdced6f9ae4aca7b97b3e18bb00794ff725ef8faea6fcba02835f66777e246ae0dd1d515644402cb30a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fcf9920b6067d83034183f9f625ce0e1d12d9510d9ed212c83038fdbd3ed73af55e27879af227c3ecedb3ef147e6046e0988c9c96432471f24031eea756aed5dfe2b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16637d4b61bcdb954a989923ca4133a36564a809404187e1837d5adf910330b5e0cf3c0a50e8a24c7d0a9830b354a83cd01530b2a07b05661d6a52538c2b56014d466;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190291ecccd567afb9ff690c88dcd82a1899a84e5bc642747e66489aa6460295bdaa2d8b7501aff9368eda88acc1cbdcfb74c29acdc5eb52d857bc445ca6771524def;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h921ebb9306bb62e93368f430c0f5f0909915ee6a175688539b4dfec9280f10a9f75713287d5c1780dcc2751cda5690ed067378f0285d677efd74d31085a3655fc3e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h172a2ef68f6b2334749e12f6992f2dea90e95a669ff1b3de22e66242a1811bfba8d0290b5e550530d59c23695277df829745a5fc09f325a9d7c4956161dfe22416994;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc4e1497bd8954c3db307882998e54994ccc042a5e4480ff2f625e9cd87304a886e9a1cbb668bdba00ae5c0430b6c5c6d155cc0bd9fc619e750562cad03375cf9d226;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa28e04c3e9764d224b0e7a0d9b0d8a153796bb3a302e71008fb776f4319a4cbb256eb4d042e0ca9726845c93dabe3521ca4ac4c90c062509f2b5ef9d272a8e6dfa5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha92ada442f2191fed998135772ec2380d297872a1b04aff563c50dc54fdcff19f152aa0d857085cd6a74ef750575a42cdb45eda21ac8ecef5cc824b72ee7f267af42;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8322bfc8f8006431a1b2cfcd234e80042158cdbefe41048fbb58fa3b7029f4f2d593a39bf7ac8b8af76abbdfaa48a6e1f5748fbc4c1eb32b892a98e19bd653815f5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbc06003bfd10d5106e8fa20bb94f96cfed23b347d141f2b76242c0897ed85594058fc718494497f6bb3762e2c36148a1d30677d578f42c9f32eb1fbea1a9bcd5c4db;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18cdb48b8218e8fa9b41ef8c91372384eb49234bb3eff009462dd68be6f1b8b36c1105e81f3360e63e241b79e8f97ef1c3a6a2dc8e321c704c36d228487b6b3c90cc7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1747529a1aba8659ac251b84501356c2858d2099d1a0405849942c6f432cba1fdd621b2bd84c3c20929d1f0e2ca5ce13852c757cd2ed3d99ec27295aed9359b10f710;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9f69cf39712428df18380452fe894414121692cf1fad9598a1a1bd31ac506a804bceb9fef0ac174703d993bd3d1b93d8ee2d47fc42fecf093ad7dc970aa42ae85c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5452d14cba32bd62a44bb4b6fbf498b500fea5ded499adc665e5abb4dc2154e80687fac853a76121a7482e2493361edd3b5262a67cc08c23bfaf6c690f4af2a0e31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc529cee93c3fdf2ef551e52ce4b16b3d62939e845a7b18c05adebcfa8890d88db3819f375501576df077725c7c98dcce596fc920e06bad6b6f516b35134140f65ba0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156a8a404c2bd37fd692e13e7baa40311a451940b5da1e4e1715e7145da0220d30809180f3645644a55132ee3f2920778685bdd36ba449c55559c88c95e9207197eaf;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb4023c31efcd1ebd3c32865d2c4e566f24b2658669dbe12c18e2baa00874578209bf4bb600f677a95e9020b8b299f648401802c43304af3af724ddefe1d2c53e3d08;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcad4ca16574a40574e9684a59551295031d12ad1bfc17c2200e64a1b25c1097493220054b83b96d14925a212578d2b0091d4b42ca1bde83aa1d2ad2e0380761da032;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e8f464dac0855f9b7e075e42a862a23116bd375b80d4ebd609b4c89109aef85fa5c6f3d5c358ac028c1a4c1a29cf79deb6ed2f54adb96ed990afe54d252d6730a094;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9251a4de5b7a56a99b171267a92815aece9a87303256933572b57f709505fc4a38e237ceb4daaaa4efa71eb60ab7bfe73cb389334aab20f494f93441e1f7f40d43e6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had4484c2d3f59fb7b4c3b628109da017c43f1b214eb609f1ca4181b3004e16afa4d98aa79cb8ce90f72be01cdc30e6eaa40b90708b93a72672f5a4d13723b89315aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h821e14a2153d7e920edf64b5ac04969a52d8c66fac533c20814e11b14beb17709cdb73c4c367939f65f090787a02cf3062ea20f84f6a1fc76cd64c10fc03a2dd4e99;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e55c23d36167184f4170dffcfd81176c7b036226ff90eb0bcec476ae7f6b821c2f5913a64d7b5ee91c49fe5902d9fdde36b7aeb5ffee8858e06c25cc4659dfc80d9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h558bbd4eff841f31dabdc92feada1a7d8d348bc043d35661b513dbd86793c04a89a7c5da643d90298d29328d1a146d93e99ecec058544dcec85be0daa8deae15cb20;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13452972bc531cc37a1f5992f02b03c773be1e4ec1c3c7740b01e9533768506e75aa48d8d2ee3f97e345ce62675f2830c529edd71973cf878d56eb87916cc884f3f31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ca8bd1fcd398ebc89c6ccdab06f3298ff84f5de7809677d7acebe2c652e47b127a394adade0d4c65875ff37b4f882905901065122dd738437a112b8b8a1455f7474;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7682860309257bc314f9d1aff53933c4fe83e890cf2c86e66ad0b762490ec85108b65e0abc4044346df93ea7f802c7cd2182277daabbb8c6cbf60e7f94c4d79cb94;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd740a77943845e6fec67b4c8a1b155934cca23195304ab319e9846a0cf878469c9f7f97e93823caf754a09a7522f7bfb7fde2ecbc613e635f5b60cce922fd1b9c11e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3eec4525eed8b19a463bb4ab537ffa30125035b568d7e7fef56d0a2fd8ada00c736482f0e0395d3cac64d3029abde6078366bdcbc017ab957de05db0320e9b2a95e7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1127812500643685eb10bd0ea6b7470f118f5a1fb04c7ebf7082993e4616374fb11892b50259a5bd02f0ac49853a12c2dd4381a7a60f487a4d3cbc9ccf6bb535a6467;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bfabaaf23af77e1355dbddd6db12256652d196fc7d352d572d998d31fae5a16b0bd371d46eb4382b0f091b3d57d1ab279724b5e0488946d354ece4d3c6ccd8f394d7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b23e44d37d91866f5fb6c7c9031843c9699295fcbb42c54e8cce4cd8d2504c80ee503a609a832730e04daff01185b429a4efd1253d6429a301f243edaf615ea19677;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1859de593bc350851915de0bec8d67e24c32643d8d063e924049fbb74ff7bbd8bcc1ef685a8c12249296ba227764f2b735bfd56318a8c23f0fec93858df62a0668392;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f687e774e2e717c37b193dfe26376c61db7057cc26368738bfc033df6b63c4d78ff49d0209508bdb31995dccdb98b15138f423d68ae7d1dcf7a769d0cf36b1c2e83;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9486c44b099d442540a1a67f9cdc6c77a77206dfbf6391b51885d5ad3eb20976aa276eae61a6633e1f87a0bc034c084e019839e673b2cb41507864274a5f244d7c5a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87d5ecc0ece6eb507664980217dacbf6d3cb766f42be47a28e135f8812aff17561fe49ba109ae8d11607783588be13c4e417d527f2b5f07586fc7a8b1c87b516266d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1959f829f5c8ada778a6b4819144213c2964c7214907e03f00fbd6d12832019d07e88191656ef6a8508ea34551a6b515ae9ec651b97bc4fcebc3a59dc23381762cf82;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8eef3d3b3776c7aaaa70c0da0da397b71408d9f0220f3f73b52987cb20b92e6f1f56e2581d9444777c339b2d7d8cc0761a632b6ecb326fec5ed7348e42a2b697ad88;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2e52577c0b8eaad3db7959e27bb80dec4c9beb9397e229673e6c0dcc39ed7fc8971cef71a5095020da566dd8efb322d170bd4c0aa7dbccba03742358d6dd8218dbb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6c59c45638405ca11f36d600c2d5caa6f781347b032d506578d5f77028667b8b4c24a6fe37cbefd3e6e6dedb00640732df4fb245e90c4933b9891aeb30a818697d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10106075608946905a43c3035c3d79a9e5e6d860ef6a77536328041dd5a6e4f3de7acc17f555c99e0fdb60e32b78465a6baf44047870f21db002beafc4564dcd8dc31;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9d6ab6367660e88ddc5132991fa780ea40225fa9e14bcf3ac662712614e2e6f1fe9c1e79e706ecde3a56111189ca35fefe273dd2a025eff1351f1e4134fee40fe13;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18a88a9a2e8506e4a47c9557fedf4f6a22416f92fc00d836d803712125173249d3de3c111c510cf73fbea2e9f86e95641bfc4bf7bf9a0f0b67eb1ed6ebbcf10a87ee6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed54980cc941e93fdfd3cb1206274711327aed1662c0e9a84b4633939641802abffe0de4d945c09fda8a6ae83f0c32ce905f6d538ec7220968e8a654e06cf002dda2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd96b7e0d770f848c1d6142da2d7545b228b67a3e5a80ddeaa827ef6f8552c030efbe9430a5309dcd385b4dea990170b8e72359990eecd3028ad4d38f0208ab675650;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60215c8a4cc10eecac6399235cc0517085a31289553526aa131d93a5125a41fc4d9577d224aed6fa1beefbbddc198c71ac7fb367db06e4f1d97d0cf293174de1cd46;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166d6e172fb6d47de88b1224d60db82026228e4e9230d49c0253373eb764f5f7cd5a5f8f6b916e26bbfe226fe6f4a3d71e084d2959b1f12ab9557ad4b6d3a61a0ba0a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea94788b6016cd1186fdd5f433455053c3bda1c7324b72c3a022235d9bc7ff461f1cb001808cae23ffbc83fc95a96482c0961ec8b7933a9601ffbeee58c8fd3a20c1;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha747e0fbf10a05921a4f2e038c51c16a76156fbb26181bcc1adbac46fddf8064b97a03fdf74a8266a4e2967c1bd0bb96e2595c812bc43c0aace7f39cef9365f904bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6dcb4ee2b3f4725714c58c315afee099b7a1fe86d934f67c9c90cfca6fe38fef07d85fe69c03c5b65f7def12e950d894aee4253415cada09daa0de89f4546961018b;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h170c01d54018ee14e9fbd977c96fa10bc78cb12acbf3ab8b87b12dad63a74e3f53d01615135b67986a6f7a0f512d0f41c11a76117a801e6363746d421c3a4654a32a4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bac6acd9b4fedb88fdb4f83777e2fd7d7986f976558494d9502f3df676cbe9d50c103c2d337f7b427b1d54a56d743f871829cd83610e83acaaa1fbe4a15a486c736d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133f120fb383d7f24f054b52f7bfebd38c6c7c12feb9dfaf1b472741ba037c2e9011a56fda9e1cb5c9c612ff30d9852e57e105c360d907e3b7c30fe801ca513ff30f7;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h31bed7427e39a60474f6172bbc8fb7c8cccc289e5f9853580c1e8c511bf8c3d097bbc74ee599efd4fdc959e3f7d93fe09724bf81001893dd7d2ca24153af75b26de4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb76db811eee4fcfc1c35470452a97ecf85b869f65f99c80c112eeb5d203d0d48794051604152c8852185c7a382b28c828730ece049f530a86eb8ca6b744f7d62dcc3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14fdece8642878d97b652f6e4ee2bf18e415d70bff7bb71d007bc3644f8e56f9d3df0752c31b20740dfed4ab8708ed3a4e9dfd7211cbf823f7af9cab713d7f76adaac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc004d2882cedcda46dd3d7bc7c2a3b8edd589b65dd3edc5ec1bc41fdb05f00a7c32f49024ade95b1d3511a246e6116519bcef329e370b5d8a96d0a37b30537d47eae;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hba791bbb6dff2a90778fd6bf160ab7ce61f5e95d4587166576f125b1d78a12b1a67d12af8b5dd6b0a9f668863f452cfb9e0a7a39ed65191da2da5bcbb8571e80751f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1055b0303022b32d29fd3bee99d6a02784da63eb7b42d72334ebc5a134da88f1c41f88487fa7f83288eb0c8ef048f3d119ff5af60fde26d9886c00d113fab557454b0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b8841f1a9e0450a04d1f844d3624c60139fdcda430d47e35a8edfabedca3ab469ed41a5a4d00e0bacf68e88c7be9808f8f683b12040721c71ff25389993f6f67650;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4c727dee0f7b9f35c144123697f0a0c56c9d2a48b8f95b3abec995b51d77d4fb3494be5c5699a5173c37c4aa52ee9764ce3fc74837045d726b1e9c0d3035b38948c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cac7b4c12754893826616495904e8edec2b536c53ba0a1d0823f9edd8d671f1478d5a18afe1d06641e24cc52b886b0fc3415ee62b2772454a151607041242692c816;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1816c51454f64dbd9dd1d462a82b6221f51a49f9766ee7ee4c16d0f4afb3da5b4aeda95c7db9db1f81ef2696e3c67025fca5c93aa9182af5dbdda7078d72a4a86c2db;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3e2522371920491620107882d41ed010876aa9bbd7c9549bd5706827dd745971551556a28d41b98d88988be69546f810e0752264a76845901b9077b3e3aca890aaa0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he82f9cc2045945ab2f41db2dac2d196f6cdd6436a38ec7ea2979cb310c4f11ab5d4caa6252f4a048e387b0d0cb48326e2662326909991a4dd17de743bdbcb76d489a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h616b4228da92975e9db77f5a8728023096643eab85ddc6325098c30c7a3f89437da38eb8dc07a5f3324a3118d215a4e37ae1fa1d1aab6b6bd7a58f66eca5c329adfe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198e941cb91b4b2458053fd99b504791ae41c4ddb7b6a868bda8f411143d781e2724099f8159f67eaab331f38e5fdaea5e634df12fee7b2bfe65674a186be6196e0aa;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a6d5971ba73d3607b963c556e0bb88bee1ca452420fce083b54a982a07a5d0f3cff54d4e0c17c8954102c748991e5d3ad8c598411ffc1e49f1f51569afc9a1d5e40;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h369fc899906b7f70b26e6635cc243c1b1ad6ee8b70fd20416fa2b527c3f5bdd011ac60199b6bc5bc8600b61c4c8b6dfeddffa1e602d044b6bc754e1fb08bd7086dfe;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5210e334070b8b03dad0b324dab98e533dec399d426ab95d592ccd1f658458df60ec41828ba88ee2498714a1cc25a43257f16820e36cfd9c24ea2b384c73b51839a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ddfdc39d41615bda4b8b1b2ed3ff4a66692774b8e23bfc976e3e80683ce84946e109ddfd6be3e5fafbe3d1b6948abb3625973afbed4dda2a729f55dfa03fb96a92ac;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h116aaa8db903babb36a8dec8bb66d3989cf8f030d90e2d67d5cf82fd6212cb9075079c3ade9907237a9d5ef82b2489050da47dcf95d56170ef81e4e1d79840c3ac04a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcae2dce724a7dbb50357d0748ff558a619c201a0e1f75bb13104386e06ef03d5d0c538e779b3a4be5b39bc4eeebd0718dcd6203bba453d9e0f3b857ae4338a7d9bb;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89101ab32548ba5d036febed6b4294594c704aa3102c05630c48ebdeb39eb4dc8f70fdef5c164dbe4fe629c70b2317914c96aec488310a0f9dca0cb86c0689d7301;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd556b266882e6217838e60f76d252539456d55802f9e8f49a92bef2fa7f48395b1680f55b8d65fdca17153cb30737765bc42b2cf1e9d2e2a4b3926e34bac44ada7b2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf5814291b8a485eb3302e7555272277205219e7fa6857897cd1fe2e8e2fb3a7379a073bbb4b788abbd23ad9e098cfc194de54de3d82459aed507580d804e52d5c941;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194581b415dacb2cea18719abf213c9dfc6e4da6035e702337c07b1bba610a8c6a43b38d6fe815c9a4f1723b408ef4c2bf349039bb1115aaac746669bf9d31232819d;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h255b147f902b147759b1834f43639d7e9b7e4673baed09ef6a9d89c03be244f9272302272834f0bc9d5efc2bdf5900735feded1abc74336ef6dd4465b9328b492b48;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ccdeb5f18454caefe3e2e4f4a37c54da842dc8752c31bc2cc0ca8aa918a7a04b5099ce395a9150ee184edc6d92bc369ba238bfc634dc5c1a5a3a7d7d2961636a88a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h154e3ea24f4cc2bebe768ffd23b02d645de39930b7cf539f2e4f305953d2b4a6ed489eca6d7f646543ccd3cab31daebe1df715b49ce61da1fb2df3cb10fe06fe7c223;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68764cb6dfb3abedeff8b6e16f0367b25bd54e6a60d0a1b53cf57f9bb83d0dc78e147ed656c80e1b0ab852fc83da3c40539ca4e7826b48bd0497dbe7acc6cbbd57e2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1653d8462c8b1276918eaf9009e2e99f7e6b1482a4347c60c3445834709bbe7dd09b182492e41b6f667a5fbb334ddda929c7f0394f4492211ef0d34b98f176a61a940;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113d99c5a2fd42a2bde787fde89c8ba73ea9fb3a95cc9e56902709aa11d829e45b8d2f17df59a107e762b459475eb5975498ea3096e8ae09c41b8e301ef50162fc5b8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14662233d033c27c85ecf15fe5a46c455bb4a9d012c8afaef8d26f66ec201edc5320368530f3eb09dec80cfe9246cc973509b8dc3f8ec59bad0cbf9195c1378ad387a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c0207836a63d1cb73f02714560e94ae66258a97a7e35f585ecb178c30092d5167214c449cc8db4f6f3fe0ce2786f9af0f372e30b2f5e821e5bd04ea7fd1f3e0448;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h37ae6a1c907ee9b3684ae19ef89c151394481c84463c78c414ed6f852c362d614c072a40c64fbcae5ca488237858c9a0335d3018cb23a9c6d66e03f59a31ba48df7e;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a03c3125f91589a2c6aee713f547bbb17d435a455d49e6fbeefe2af0bdc6e6ba5ac49881eff6ddeb4d05ff23c41a4e9bc83114605aee202934d43cd4c6dce15dbc2;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h77887bdded607a15c967333a39c940f17d5d3fcda7040ae69e917307bb94f5b263c037c39eefcdac73ae114bd519d52c2632601661d43f77b6a7dc22a9e36b024372;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h809d6d628c1f02cc1846e0021c47f8a7c16bb71674a3fa2a61a0ab95eed3a569953255a7181b66badde94eb2cc6bd3a098dca894e331ee8da09e1a1682426a76a20a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha1302c9d74f943ed08c595c95b55e47b6f6d8803a84a44787710628c486e558bd4975070add586f81be882ab9daa69304b6f09d4e9a50116d21e3b758427dc6bee63;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h294dd7a9554600221fff90283164ebebad8c3c25a41827a2866db6b858656788758abd27c3be639b2219c88683ffce126269ed88c2d6fb61d14564e9658103f02c5;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h122317a15f6c6483fb4079fc5d83b325c1d9b479fdd471f9d8a59126d4ad1c8fadc2742e7abe7e4aa63c0f8d328ef1b9c2d3ca1c904cf33df62a65490b732aefb96b3;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2ba82a15156b8b3b1dfc643838a34f84d6182a0cdf1d32c3d63c5aa78ff4b09a0d971707b8f4b12208661bb1e7bb03f37d9498d7f6d44ea21c603eefd7b0156c30f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f0aaa99b3f1b17e4607b0fc1c16da97bca9f7e83a42a1881f15d9b325cff3240860f8c3b7660fb10a0ab55dab7d2029ab45f83ec676e713a0f8f3e8927cddc3067;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11639998ef4f95a89b0af24035cf0f9b3dfdf06875f8541a82ac9fe61f7c58f6bf89217c77d253568aef3dcae45f5b56a7bd03cd450fefb0128103d9a826b5b2a11f9;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfba8d440d4b72500d5d3847d26220e22cf035d7f6f790c1297128f84894b6cf304b3a5f9a53edf0e8fd794a49088a0919f873c1e68be8eafb9f04b714a38644eb330;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13fce69eaa788d893d72497a3e23527757aabe79e1a38e8d6fc84b41fdd636a82b871788ef8066087cacde73d5d13344db72e8fa14a50503838e5a26ce68b649c929c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h87ccebec780c43c88f21ee2fd5321d0d6bf25bf7abbb2cb5e141dfbf4569e52aab598916721aa0b84f3afd0d945ed8f96f4306583e3a818fdd4ee754b8c6e4cc02c0;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf7763ce32634891bb75074afda10ec47d9e4141e89cda92948d80575ac6eef1549e14e74efbdd6249d67dcb6a1e0ea83ffb2a00990496553749622badee8cb52d403;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h590bb20e2bb8181556d244155c20d8204a12e80dc10bb3e79dff9345a0416f8cbed4d80538bcac3d321c4c96f4fd5e46360d44d01258af8d1dace95763799e9bb802;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h50fca71e5fc95e8b8318d5907f15227b58f38607d0b762950025aa9e794931d185c8d5df4f2066d8961afcc1508377ed21ed90993a3e5b4330edaec7b988c8a63004;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ae02f9f09dcdb45b07b1439b272c2c91874e9454842ac6aa83c4df36d20074389176187fb4b249bc1052d1ca776a85631af6d6666284cafcf61c60d463ba40a0e1fc;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66f67ada3924acccae1bcea2cc8c0153644bdeae2db08f5ccf7d489c5295182e16bd13b6f196a472fa1c761093c891806796bc64e51137bbba6a033b4bc6c05dae8;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eb7625f8eee069515ce6afeef300cec37810c501dfe8e1b93083ce10364bcccedf24ad135cfd54f254a7b64363fa7bf83bd1475e98ae582d58a31942db1d34f60c11;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e6252a006b009d66ce80bd591b51ccde95ef3744c37b7cbf96d9528576e51e2f8259d8ab2beb5ab5c4413872c027816bb3c7eb7b958aa7f799c533774d80bc4b71c;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h90717a6c04d0c011fc5b08565539e74a29dbc3e37b7a3c7fd18f5d3595a9bca4b1530008064aa91ec8e9ced493b40c0a51ca817630eac151f13f438fa537e3610020;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11b63c8710f60d85c250a87d640c303a39adce360053bf1eefb3a1dfa41c63a3fa65559ea4b7163406922add31b9a9d4dac90be7c4711668937f573bea9fb9d4abb87;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb1298876899894d38ec6f21763ac653a5d6bac01a4d710d318b33df9d58731fcf94668f0d2295f1e89252fa3db7d3820424561a38e72d3a90c84cf97def52153e221;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1286b81f1d52e3545e1a2ae629b2900ebe9305e09b8de590de897858b83ee326d180b8196aef35335eff42349304a3bba1434e77619a4c1f752881220e685e146c0c6;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c04088a3e156d591149717fc188f01a6eceab31c76c3d2df7ba3c0dd926f8761e4f537884c46d62097a762b06a9250a055353f3917c16a69c17679fb618e59711a;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d96b50f04a72b7e9c66404f24d7bce6628abb0547ab350d4fb4e545c456cb44277c686a4c7d9e0def55aabcf9438c07d5c87d6d4eed74689c4d4258155081d5b45f;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81654e0822488887ef85760fceffb6c32db56e2e441f86bd4669dfbc7187ca6bc5f128194fbc4e530832617914b9153b16b29fcb368d21085288954968edad72a232;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14923833abe0bc7725c28a414759be074a9dba60a87df4f3e940dca1753af0350883aafd3704aef2be0cd43ef0811f4525f62e7d7975304b03bef1861470454e508b4;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c90c95053e6c2f49995e146218cafe81f341dce551f55b47202c2dca2954b253aa2e1e31298e77d08cff243a9e5274942162ee4c8c4ba3d301315e518c3ff3ccb64;
        #1
        {src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e29e76a64f169d5da92beae0a86fdfb350c49fd391d83c02921250cc80655c06d4fef2eba04d5dee451f43b3a9d3de6110df6f6241566ac91ad48c75edf6ed3b7e7;
        #1
        $finish();
    end
endmodule
