module testbench();
    reg [17:0] src0;
    reg [17:0] src1;
    reg [17:0] src2;
    reg [17:0] src3;
    reg [17:0] src4;
    reg [17:0] src5;
    reg [17:0] src6;
    reg [17:0] src7;
    reg [17:0] src8;
    reg [17:0] src9;
    reg [17:0] src10;
    reg [17:0] src11;
    reg [17:0] src12;
    reg [17:0] src13;
    reg [17:0] src14;
    reg [17:0] src15;
    reg [17:0] src16;
    reg [17:0] src17;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [22:0] srcsum;
    wire [22:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55b9e0371ec17ba843c3cfd75bf037450968ba41f4d56bb9fc028d1dfaebc4ef2778eb2df9f2646c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13083c64146785df5cfcb2690ca8ed2f4a04e500a883edb8c0b225bf420c93e4aaf163a13198ff41b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f0f7501eccbc0b3461e25f79744ff89544f3c8dad041c22842214a9f7a0fae6583529cde70c614a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h444aafe095e175867c2e88ad4e2a77bc3c7905ea193e0baf3ba5accf98702163f7ad574df3f3ae53c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha759b67d24c0ccb5027b8d3ee4b052aa36ca28b16c4a67a54b87bb720433fb0d6a944d5fef424562c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9cc686938a38329e297892dd54cba3b5f7458f6f6e82526625578359d4a7fb7c997fa7e9afd8eed09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70d7e217ab8f2704b9a47216df7de6d854d7c3e71b09d88c042cde25707e6901e7576f13c53319a01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e7fff129ff171501c4e4ac415b709b818685ea4166f39173963338518bb8fdbfd5d9c97f16a038ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h356e9fa519bdb8aa70e50529a696214543e4529fe630733d9b6f5702144f924de0fc5a215ce83f37f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf13d58bbc48b66302142588f644ffceed1f6033e5dc6212c0eb5f4bb666a1f509c78e5226eb028;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a9215a69d3811f11823a29be2bbe20e549e17d0bfb5913d73f7c8aa95421ba582d13ba4646a441ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc331c747f4b3e313212c499064e17aa9a812e533e04fb16423c166880fe8add8a020080f51f9414cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81c27f73b96b2744b758d5eb3a0c6970fe7fc0d8888694fea281e46d84ba20672c48b37b2f6613401;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd142a643a161aba6c642fe4b988de32e40f569b9179b946d3d305312154a9b686b91dfe68bc657152;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4895d94de07a81ec529b9b85df732dfbf87fb0f7e586bf15e0b8b0f349a1d57a72506b8f99d2f2243;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cce0399c2546ba3d0a0207e3c718b9242f809f9e8db0909c2e6b263a9af16cf23c4f957d6ce8a7cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6445132ec99cb3ef142ee2841c4e40a120c94dcb10b96cd84350e10ae5c0337d9513a63378b8d6b02;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6870386d213685ecf6aff03afb6f768b597a0385f02c10b55b1d2829bb8fa0c3001ef53a1cca017d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f641aa2e4d0f7eff2b5ed5ca7921678ec8002a6457bf86b57a4a5bb262e60a2fa5adf67e4e8fe74b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7df13c2b71ccf2f2567bd9e1b96b7f616fbc069e95f713ea4085c412214600fcedaac348e5ea7dc5e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8af77e21c056bee242486e528251b3314fe23d2db79df3c6db47d7c1eff8d2cd0297b1393716804fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h387e4600b2414fae8cc506bcab83a735b6aa2a4cf7852114422a5d03d4201879acdf21e74434564ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9aca475d5cd1791d93852b740c9f9cfe0bd375357b0c799f25d9a33f80a1797c430b226b0960d5170;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd35ee9a57a5086228dc4d5efc96d456aa0c728983d5a0f7ba8fb10daa21bc5120046f25bac0a357c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb45c27c064bf9f60095358607b9f0964602b75b9baa88695bddd757ff6378e42cb10a4524eae8297;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d13303d85b589602ca9abee011ed34b89908a1a6cac68c914d756e497bc482e0c3ac7e9af16842a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3941b4e367955cad026d2548cc9ff91e1be92656752b7dd49a3db7b0b56d9397cddd2543822685bac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fbe36f89837109b5c4bc8a7c549ac6d669f1e4cbbcc88f7309df38618bd28948d11a12c61a47a9f0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf646b7d01c82c972c3c4cf1447eb008a573d5cb9f42765cf0001dd29bbc1c276184ab8503eddc94a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc7421fab99c75bbcb429ede4039c401af7aaa511930528ac42661abf8eae6858f75c64fcf7b47ba0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28ef1dc7b4c095a01474d5eb3a13c7003535c871b86e455713d599334e8acd3dc9093bc723d385133;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82f9f53448a45889686dc0f7cbe2dfbae7ffe3ddf7c7dd8dabbc6a37ed19b2bbba30fd29c2864d7c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcacbb8cb0fbc01284cf1563e2a550e891cf82f3dcd26d0e30407818dd88275399efebda3492bd27a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b472b1c4b03a8f398d7d1995114384d6039b1c16ad9b80ee42e3af22c9b126775ec13f9467110b39;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e749b26308d55438bf8e989689a2a135c9a2d4306984dc903de5eeb7d82cb922ca3519534dc536ba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h415c84423891d4f38d15f5d44c978629837e8636a1dcfe4e28d6d259033d4c7fb95df97077e1466d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6ed8cab60213cc1f55b16a59fd327901a3e902bcc594c1dfef19808f2103e54f6c66761b24f7fbd0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd28233d2a818348218c6f1b46e29c0ae42c54de6b1267fba9a8600a42e96a50235bbe6048a5da4765;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f953f29c8223faedb655b103fd42c82685bc4efdd26d447cbf8e6067e4ef7c0213d2d3c7ad053702;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0f964aa9b5e9a208b2db7678853e1270358e46b992052ee54f18fcec784881f92564bbb029d0e078;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb84e35966a87b869f42dc24c1612b9f9a4cdd777e5bd27271a5a018bb4a0f8dea4827d605c5ab392;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he397a8505a88dc7654c1de3d7da37fa61775b11a5721f2e415509050326684755f55dd973b8f140bf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83503a9d6102f41ccb09776792daf80887a6456077e416f2a6205ab42f91b7d9bad39690733b8bf76;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbce02889f837a7379d9ecc1203b67d26b7a4ae873b26b09281228d3d11f41ca2cc1f0455d8b5ab52b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2021717ef5a3812eb8eb28e7ca2e428895fb3969f659d9a8139eabb8490e947b64c2904198075fbf0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e0cf54a425febbd4adadd46d549631bc8da352f076543480e069573e8d5df1725c9a27cb3584e536;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff9212f2801ef292888e57c60c1a796640bca24b7feb95b43626facc81731cb4f14d5b7aa992a89ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9363ce1b9af914ecd08f35b5c67c34fa0230958f86598b4b36395f7974dde308cf1fa81becbf9ff28;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41dcc8784e9c1302eda7025e1cf0a14166f37c113088ce6e35279d977032392974e11cc30e90eda83;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd88ce9113419d28443688f093a855be82503e4fce720f1be5b5a47977b83eeeb4879cd827fc2e935e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ae749505527a1d53a6f0d8c507e5d8c1d3e3dbeb7cc14b9c3e4c8ada5ecde9ef621a93279736b284;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80f851d0be40458262dda684a804527985a80cecbfa2d42467e4184f3f3b0551d6fb75852a9a9d010;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30954e0723bca6b7a1e7c3417b386cf529d2f07e987c4c03a321fb2f2f5b0de5e456c9bcfe900b918;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd192dcb85e0a045ac9944c5e0f4035eac723099afeb443e3065a75367ce52ad49f8c14e3abc1b160;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bc86f3829dc1ee10a69d9ee37acffeb9e12c5ae195f16f928e3d8e9b088f543cfbc0ccc90fce313a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4b65b08cc71e74a88128110ed473d6fb4bc6600e589db813261c4fbd4f9c69309d6f6822568345f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ccb3194233dfd99aff94939efa3a0903777a6d25de78cc8a92adb848f14e89b0bd354fc5fc3cb124;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf44d832229c7f7389982cf3072f6d9b803ce0d13e5d5975052092f0527d3c70f8d1c1376657f05348;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb650cf242448883ff66d72345ff0385cfee5cfe0f0cd213da88c55501b9f948c22465ddc7b2e52834;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a368b6e1c840bd33970ae943d9938ff64dc5698a58699d29ae25ed4bc51cd99a8c0c1545f1bf5b85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2408738b8026508dbe1df17e95db93f6fa39468c9ed22dd238b3adf094c16f7030e6f697cfe58d44c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8eaa3a21e35071ac7c1a5270f533c4cafcec9016db8bb5faa116d502fb9fd7bb1b13115afc8e982eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf6791e311cabd56a74f70724262de7aa918f010b0db2f11d39f2a9fbaa34e42f9b17197b67d444d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5b25cf486c9d8556795fe1e1d7b6a9e324cb94030adc347835317b9f30f04e42e805e058a6017096;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd79dd494907ed7ba7ef2d654bf652616c5715882957276c05d3da83b4bf4820bb5d5e7ff50734a69;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbde246ae9f1375df19884ec9e829e36a67d9e2ef7258716c27b1fdcbdb1dde225b1f84e0d9215215;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb69ba0df32fe4ea8e8cb5a471346255131d80a0e3dbcc90032caabfb9f2b5e5dcbc0104ba4d9149e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5836822b2a61025891a5acbf5b9cf67f1f7304d62a387c17f7139214f84ebae3c24369168749aa415;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34ca3c19e3b83a63a92b2c415b4b623402155a8ac3cdcadeb0f3f1bc462d65745dfebb35c0f728c01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16f30cede7a861e14290c3e73342af82e580adf0e927b19ca6313b6d0e8f569145cde330586bdc00f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac847a0d28ef0d98af7e0d34478c5e48ab926904ff3f31f87293779118a5eaf1c7aea1e19dd8ac3cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h242e59ab9011bb8637a068f14810c0a8e115b1fe382c18c1f9a464940b169c1305686456e5f2c25ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he622d1a14dfb7eb3d2904eb9a734b87b1c70d0000dec0f1354919958ba99804a696056e3d6b1fe26d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88640c31371bd0c383465d0bc66bd59f3efb545187b733a4eb72b6b5d6a5748e91bcc3ecc0c81831e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h160349b90d2f925715a1f5459fb52491b6b55bc34e8064ad1ab6568a587fe3d0ad9661812f4aa8e7a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he8b4f957982ab08709b1f32ea6cfecf531f2c6fc48c6df1c63eaa4bcf8742367ce96005783c88d220;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7fb8dac67fd5adf8120c897de4d87e66377a32ddc6292594bca1e424cf15d89707ee0299c0bcda1e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4edea90d0fd189e329ba0f591c2e46147c64ace81dc18d20bfac30434af95c3291627ee81ca0c51a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h547d6512802dec3124cf30bc4dac7a9c882f0cee086fe015a60f4d249e028cdaf82c7f9f1a6811a2c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6195e56d87b0ea696b9933b2549ebad8f524adfaff9be57afcd54b7147c71bf212df8448cf3f8270f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h276e0653b795e49359429d30d9717ff3bb4bb1722d0fb0d151489dccc9b2dac6b7f46eb1fb16fd1fe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ee418b0e987ab24d48d3bcd17af03804db5f152a14bf49a861d9a2569d62ac6f8a014878b42bc61f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda6b59b9f44a03c101f6d4f3738068976a810dff22fe8841a64ebc79c239572ac42f06049150d326;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d7cdd76970f0a1a79bfa2f7c57ea26dac71a1db4480bdc5ff16ca4e4c4301014ac8884e7997f3244;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e92310ce5736c9ab157e0541237c4db021fa0097c0dde3d483b0d500a2fd6065a69658ef104f6272;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd2df5d78eb53539c275191099ba3b8c3ae1e85bbf7c6ea5dae080afd84c86cd76e0a996800739998;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h73615172a3881029e03e9561c342a9181bb375f7d8c593168dba5967de689bcff3bab2c4e3aced61d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf3fa9a06561b624bebdb8a3ecef2b28cdfcca7f6c91240733232819800124b9e03e297e71e10c8fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8593821d60d0003843fce39727ad86c7ca23c9984bfd44be271d38ae3f0211fd2b1311bd355bedbf3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58f4f8c0be87122386666c081fb24cf615d1336e9c6d5021d2981484011eca9809801225e4804fd87;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h947c690b2684124bfc4ba97cf8105f19d1c49f6f53accd8c283896670e09df3f7b88062f88a30136e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77156d7b334aafab2d7c09c2d0341d9234c103e03887bdc4f90b0b460a11a3b1fe93db59372d5ca5f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61f8e74ee60596f71dec08b3298c84e6236ead2cdf8aeb699587f52c46ab4a8de47a815051d048327;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84640776539976a732df08f864467609b16900e7512e656d22d748747f0aa5e83526709ba33df96cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he94b13d337c28658b653c5fd0f8fc2efa3622127350ce8f03ec9229209901336328fc27d2fa974daf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e867f8ecc7e4cc7c125d51413cbc915d5546ec986060d4f5e94af5af4c679a5216b0d9814b0702eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he751e3ddc0bb70eed2eea938dc9834b2fe9b191992c5462d93a1b712ba3a49cf03f9d8d10d7dad84d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba6837a565307143ca5ed249eb878610523397f6e838ce77ecc75735758b5736e37c3d6165f180e8c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7868d88a5353216049f99ed4c1d85f68bb60a8e22d8fcca35edcb5d5a736f3bf691bf2fb0b62eef78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8301b4647a1cf05f67f4a8c89adc2972740509e07f75426b63e7d281bc6d5711eb530bf633d354b49;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10a68b2f7013778cb8882fe34c03acd93364edf1bb9f7a707fc9898fd19844562d3b2f15d9a50c787;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb66f82ce829c9aeddd36945fec10432360f5e3b323fdb0f275305996575e4550c6225663c8aebe5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac2bb1b703aff682797fdd5ddc4b03faafe3df878bd2f4a837ad312ed3066b9e9426508a064b4e9b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79f5de11dfd08f78497a1083cfc0db4117c0c0fd8baef97bc396f346205c8333e38c5007a1ffbd6cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2874f6ccc41403dd942fa20efe5680765d7d7e9a0b087494be22c8f1548f9e9cbd8a4404bb62900a6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30aa19cdbef2960161e45f8b102536ccee9bd3cf18765e035dfce5b55f09f2641d28ba4beccede759;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8774e64de02fe9853d148d4926bf358b77f2887e0596cc73e01dd958d0d18065496bc3277f69b716;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64d1010482c8561689b3b23e0b3d8e257be270c19ca6de30923af4c5c31075c284749496049c39cb1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f31bbaf4fb057e92b533dffeceda78b55556ee7ce2059c0686f65aa1b4be5fed0cb054fbf71e80ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67e20309a7895eb8c62d504a35971f2d9c68a18fec4c3a9842086dff2b4d8b0416a020325fac6c64;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6116fcb51220b9ad05b907f5fa7075dff7c17a9d4423cf4d6be42fb5b7553b59a8106d8b688e6e772;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59612da8b065429ff93729928918600932c7ebd1f64732e5f0d44f5bef70291a7598ac953fc0131a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67d623efce84192baee634a152d28a0299c950b88e7c5478cb5d3f3ae8f920ea7946771b5c48ae608;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a02dd007804c5e94b1b11fc1b5bd288fbe9ece144900c119131f4a2030726a4dbaeefda29c09ef8e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dd5571c3840dd46ef2f17aac25a5db75614cc8a90789dfd52daba1c00f6796b30c34d9516eb966ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5eaa815088a2bf25cad7a11c8fd2417a3577df9c396ce8a48f21f4198b1be32349c15cf8e49de7cdd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4df66c5084f6aced1c007758d1c9bfc05450995d6a6de489b33908ccc47e147d5f85a206bf1d55493;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1235c7a19d6db6b7d4ea95ddd5dbe2a16213ca1f9b7bc0f8fe3d4fd45554f479002db792f7a346618;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46ec7ea2f337395fb37f52bb60e904b1ed318277f4d6ab42e3ebcebd3d5d7d1b7e7c7399558bd33a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6eda0d37c8db79d7056f93d738cad5a8c63962c13cb078d36369d3cceee575e2aee4cd00153c2c2d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h631fd007b9f4efb1a58cc6fdfe245a41b7f70a3ab9c790539c5e3cd60f2b34530f97bab79cd39ed47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfacf6c817dad6730ebce12738bca963231d7f9e446494c717460ab3a25f76a59dfc88aaa86c14b3fe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd73b51b72b1c71c1e686831a9c6383ea49f1df40c2ccfb6eccbca529d8f6981ab9733d41a55480af8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d3e5315c95e89372683d85eb7bf2ebc421fc5e1e42691fc700ba03c9a5a0b5decf39bb465c4fd5cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a7c98b84cb2d988f3e2348d18e906f7bc8b67f9ba788f4252bb3cb06c18566fbd0aea7da7f95a7f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3e771bcab7114a7088c334060eea0216b26579d878a89dedc36b9652fda87fe9b38baa41d2ad52f1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc663548c48fb3bf439f92166dbf56f33a34e8d7ed6b5f05f671c71301b0fb5f1cd6649dd5a67e4617;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3699cf5b1cb8d06af56513c4c4868b185c50d389d52a741d7a0970b1de23d1a0b0bff11bd4390f35;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a4332160bb636a19e2bab010d1dfff4147151b60b0b44acfb87d685e4d5e042050cabf112270188a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9376337b079cd7e721c2671d07e4b1e7ea9bd38078913d07282cfd748a48cd31e6bd0bc06ad483cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93e83aa5c8cc6d6729504ecb5262a6c027b4cbdb39052e942776fd80e6cbc021a8475549f819080d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h784e4fe94b24568d95ac3aa1895608fb409fbbc1d14cad9b97236b99d72f0a7b615192f9ee251b1f1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d36823e2970cb4de588584c286ab183fc5e055ab9b900d2f435c31700bef19042a5b15b3a374bfbd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21a119a90b12514eaa5a906c037b91cb96e48e6462c26f15cf9b08cc838589977d00e21d936568a19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dd8be2f7f2848952d7613a7f1579ca1e726b59be5edfb0c2c2ad6d113c839f8c0e404efe12eefa7f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd9ccbe6f3789e1d02dd7f100d17e2b72f1d1d5ce9753b16c9f03a36a9e56c0d3e6e5658195506945;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha71baade33f378f2b26b4342d3f58743fa87fc63b29fdd8f56343dd9ae48ef36e799cfa8c95606ffb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b037abf555da78e9414424f739b860b13ed25acde68b79ab2ec9eb0ec2157580c19710bd086d9b1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2c76c0c23aefdbb34ecec4700da6d75349e328b58fe0c7e0710bffea4818beb2bf244ed1eceb4364;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0eaddca61e768100024f8b8f891d42b5b58d4eccd661701deebd8444420ee3b6a9829fca3555aebb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd905fac645b42abc3960ae3d733af9a98bc3b9fad1c7d0cb61ee3c5810aba052f8114064bb7349dcb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1a69ed39226191933a3217faad1ca22096e1317bb52eb2ee19c083cfe7b7f8bd862e7114d0afaa7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf15843c038a59466d82439073b30e017caf4157f789e1f11efca934472426c16b793ca08bdb97e4bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3994de78f5bc85d282cf8c77feb246d330e692cf69eba45636486c6285ec0a2551b3a5d2cb7568b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa99e2e5e61801582a051ac410502f65e27de13287b9d70fb245a54fdb156d10c46a2b881fa85062f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddf3892f73c03034dea16f6558254d0e78a293ba0ca7fc98bf1f13e20f1e5f83c998becf55a9d9bed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a0a2f98b2c9d8e3de793650256827c2bd844eb6345131b122b7a9f821e38aa3298a25a57c4019f45;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d3a3b3d0483efba7d2ca0f0cbc4a57b42d6229d6b5dbf3d4183de1ade3d8bbb1eda595f991883b9c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc51cff468086322f3fc68376af05e8376cb34bf7050632eaabe2017ebacb6dbf798c283ae3b8c7f50;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ca9c027acaafacbf3138e9e43eb063338ede3f5583fc601e5734d6f0c4812064917fd4b06cc14a7d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb63332b201b27ff982d9acf713edd15ff6e6a3c195de7792501bc53ac85f873000a3d4546d1436698;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d78e2baeb849c39a031c11353b6ae7f838840cd7447bbcf6b4503cd9e79197b2333171999b1479c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4f3d77957092de6ec1d6549c31affa84811a3944124c23f91d1dd54270d4e69b165bdf1c27c1c75a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5efcd79eb4c3186de76179941e6f528ab46487897951cb773a99f6d8fc47bfac07cf3d0adb5716049;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h724901aba482a75a5c6fda9373523c37b801115dd1d4e6677271b0475c53f70049f3b6098c5f26405;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb0315e52dc483fa5ee9dfdde0e769866603f67985aa306d73ddf4e4a9a518fdfac53d581d6b35252;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6841c1dcbe1174470fef52175cb32840b71aed32c37a0832971484e33f252ec29a65c524290762407;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h299464829b40c3d6126f7bae86af0314dfb4e8dc0cdbda6cae87f14db097f44a110eb79ae5cd44185;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd096d2abf106976ec6490858cdbbbdb0c6fd7f5120a07385c8a7bdae3ac1b76acf4986cf95690f5d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2483ba732983d6592f903c5cab6e0f2ef37075877aa4ed99cb1fef2a7cff82fa5c7bec64fa3163fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb3658940bfecbfb3e9c4d08604ed7c9d4d1cdec2901b640dda8ebcc16143691be0ca758f32108158;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff31c8b0c9c54c82eb8ca29052d356d221fa90eebc4d98c965619a2ab6fa475c7ee005ec83134af7f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43078794a764825f32691c7f665b5991bbd17fb57b89a3bf3c5fcbeb9233f31e198d0d1b91dfb323d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf7adf849266a6871b207750fffadb1da8c096240624601f4a2e441094ad5cb8272a02c8459cdeb9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f7bdc0c254c58111cf7979b177fede6ee097f5544880ffb0fef28843dda8e82daebb705d3bf3dc15;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5db72de62e7bbdecb12add761e2d85d82a4da8e7adac0987af6795010e36cda8dd366e6b760bef5be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba07cc11d357a710ef4702706fb88882fb5006e88dec4c8d3cbc00286044c08523f936c66e2a9609b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5dbd8513e3fce302d436011e4c407f503bd0bbab709b409976cd103ee654ec9c2945884195c8cfe25;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7eea14668590069a67fdf368940eec4cec7ae93375fa8f196b2b03607f111869d4c38b5cbe320e799;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2303888cbf602cca557fe1644b613e4cf07d7f20110004bea66b73fc4783a5f391afcd669db33b1f1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he045d484983b1fc4853b475dc327af0c94bc6b666b3f3e25d7c9df00e51a2ad6a088840a49065898d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8fae4cb37200f3bd6acb4b75f4abed230f99b2bbfd6f15a8cf913cca6fc7e1a7017544a9ac18984b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h994e079cab3bbf5d83891aa5aeef3ef8f26bf0639251d1be4c7473f6a4f699963776fdf4bbf0e9ec3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf1a07a8b49077efd8f41852082d1ff7ef80050c92be3766bc872214c6b96b3970f7f329c3737ebe4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6ca0e7a693dead7f1cf9dd1e3194ce6d4908f1aacb638fce193df29a64df94978ff93341f8815a30;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fe12f48734b27ba19a82f425bd84d7d94f0404ec921ff6b6034c66b44f86a63f7eeecb284ff54c33;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49ddbf1e4a28bc1e0ff311b6d01055b26ed883ff79ab104b402d0d5d971901120e3efcc6b8d026de1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he157cfaa005df043a6408d0d079442cefb0bcfaa60ecf97b6203377b05dc4442448144a982dbbdca4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ba962459943764c05c079fd61961363a3cc257639db1ab0a3d227a1bc46e3a6351e2f10940b8764;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6a3a310b0bbd6387a4fe7ec02f6c893b4857cb1ef4cf7f4bc9af419aab9e18b27c19babe7b027df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c41d38c78f0be792eff2c9d2948bf75a1a516e17a54469dceadf704f74554ad2007f23c3761fede2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7cc371ea118e370c557d3709d8c2191b24c42daea14ba543947e010b0abc5fb8ba779ce82f50b439;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd03aa096d0d664974c01fc9569b0ecbfa69d4022e703c626459eddbab189b90b7a346627d7a6cb13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafe852cfec2b42e9101cf633b376144333bde5e39e88138b32472ba75c2365939463668c140bde008;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93702f5382ea31f7aa0c4f4461f6aeb6ae82df2b25115c503b46ab6a1389bfbbff342f92188e2f0a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc2f1aa1fcc7dd57aace62a377649d3c7760f340760c1083182072ad9f0d11b55d474793257aaeba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h615be05654f20eeffae457dc69e95f875b8f35fae16f128befb9df24bd7391c9133a08cd1c867c8e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a2b341673ee3170a2c895edf2aec6362c3ff9075f778012b6cf278bc2083f2265e159bbd994c5879;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f2dc1cdb6a160df4f37b128acc8251fb1dba9eb92aefb434e5bb9e6340ed3c3c77424cc8dccb7c08;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b79af3e61b7cbcd1ec255c05b77c515ab17355216f146a5b0a5aeeec3f7c16cb28ea3f12ee28ef10;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d53c2862263d198b7b3f114f036b2c3cefb83186e02d825cf69b175d30b1922b8c74e08f8e1c2be0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b6bc49818f9912f984b782d7832aa585a719f04d914dfe8e29aeca8dacf8231d9eab658b389fa52d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3700efa66a9012853ac39275299d887eb47d0e80a6169a17b4c6db9a1496eb228bdd2dc915644ac46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf65b0dfd590a7575ea51816f62c271bea91e1e7f3e08bcf298d37aa9b7b1cf19eca8469b77f2c131e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1def0d8adb19dcd67eba9468c390f72c7533192fbea39ed6302d6f953cec602c4f5c30d4ae68fd2bd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he636932c3c6e5eb107eeea167d76472a28c016f6017ea488f230a80d3c28f3c840d11bfb817ce17de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd091c28542d5a19b629c4b67de63b495b89bc6a044065be720426fc19520540cb488a711358b53a44;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81012bc34822e1e0326ebf5ef94c9320e49ca8a96be30f06c42c0ccdc8aa1d5d3534636993d1bdca3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h380b4e328e7d47f04d2b324e51a4d187a7d5e4a8aa8dcc77d99286cdc1e2c0290a2dab7a164c2ba01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1be4e6718334fd96313d5aea1c389e016083274c2ec357c4a8cfd23f107f54bca3a06f9df28d4e05;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4172c196779f2d1629154c729299fb238f0a0190f5c4433ca8ac8fe8210d204e4ffa57c0d598e2712;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7e6f092e8f0797a8913f9cc7a321c13c4854306ae8b6e51ca1108997f36c011e786ce1a2568858bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha187d6c9b2024660540ea186f3c47b0886d136cf3f2212048c8f01199ca6fd81e5fa769ae97fa5ac4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h966ac534749cd729f00d35d220dc546e1eb2c6659b1bc015b49da40488f183f19ac84845ad8c550d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf529e2e756e725800c8af89ce3c6b623a2eb986c617f08d2a2e7b1cf31f511fde8226082f667717f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80d93e82ebd942c7a94039abeed4ed22a107b728ca8d98be82008c4f1bf2f6fbba81ee453e8596a25;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9196bdb774036cdcebb360dde1017e63507e274e81bdc5b079df6224dbf223383c03c13a2de2aee5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc99f9f9077d1423f0144486b67e97a02f004d16ca22556604bca29baf135f24ab347a911e585df9b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fcd68e435b25d2b47afe6db0282a6faf3e0865c8317385f175027b1f7a932e6a1f6cdd4cebb3ca92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hceb51f7fdeaee0d900f1965bc7d26a89b63869f2a3c2269f5d0bb76cac994372135985a4438347870;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfabbb5527872a8251e4b45fb07053e3fb721a4552dfd3a6afe4d142c53e1907d16a3f0cc52f5e7c5b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd3d8698fff21e3dabc472025dacae2ef43d8049e180d2d7071a2ef138fc14fc3f4d1b6d956cfbd88;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bc6cfd5ef5ee8ba32c7b6230de9ead46ea37ce1f289af33cc88d271420e93637841b6aba188fd2e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24e69f5ba31ec50601dbab20c6d8e242f30f3d7e6dcce8ef3deb3e114aa38267cbeaa24889c38a77e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he46292b813c5575f54ffb490f070b509e9dcee3d7c280a7620104c67b62cfa61078eb5d627c330421;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c3db60fd43758a0a3995ff35be4b19214e6ff948734f48863d8d0abe1c87dc94ebf2d83ac20900d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc35e4cbb2595540e01a757c5c2777520eb3c2f70ca1f22ccc2ac0df325435cf83663f1fbb63b3d652;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec0a12741b6494b0fac148130c46b51df4a091184191c9843387e0f929b2abcedcfc8e9497ee9afac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h885fcc1709adade676c0a44b8bb3029c3f7601303896f05440b2c4e8603aa04eb73b4dcbc274d003e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3825634055bcd1dfecd9c903eab8a8d3307d8f3041f784884f37591c43d2423a2450fb39c05895cd9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcadf0744a868227258d823d3a31b251e78720da622c06f9bc30e8b7a39a074ee90ebd37adbb4ba1e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h83ed76608a17f8a8637517282dfcd4470db1b733b13fabdceadfa453f1a29a06be84bc94f5f53fe09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc797f3b5c128cbe4a6354783c3b41ce751464f96f579688698e4581538ddb8e1a4d1c396953f538ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77da77bccb2459c6e0cc451b684ade674b9fcc16eed3654c35492e140c949128a1ab9497a3d117029;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18d9335127abdb8a40aee8a50f81a8ecc483695bc2bef98f31c06ed4bf7a408aebd9f097f764d7c93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8798c1ae3ede4fcb8befe34feed4cff877d3ce84dc540569515bc20a8d6d7c34caa5eed9eec250505;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae459ec046995c0a27946b894de9a83e173fd8826377f59b63d7902aa01cdec7e4bf585cf7a1a10e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he847419a951af2e4279043742fba715f4cf4df1312600856c3442ca08c267c7687084b5c0aa0092a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha22f2796520f643dfaff5678a96da9dad53a0962cfc714336f4d9d6860eff052c5d0bf28e301f29b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30a795a6f719664cac5597660e228f46cb36f3b6af6548974bf399cf232fd7dc7475457ab80219991;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b39481e7ee3c3ad87d1f3c79e3a642ebdd35bc8f33d39e20a80ea076a78569e0b70eaaf88b3396c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37219d830de3c9c2c1a6ccef62e33480e44cb6dd89c0f32b286dcd73109f5a25a8935fbe59e4736e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe60fe49547996bf98251fe0c0560c0887dba95472da8fd6f9b9a377d7f58b0882308c588d89b86f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hccde98cd0906283fe9cb3232c5685d8ec96a646de5443119b1287b758e95d40433d1214637c80df36;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0edcfe3461c4dfbc963b959c493789a08dba7fa2577ebd876a93c97b9cfabef9225f8a6ec9bdface;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h847cbeb02a3366e7e24107b127043d21c16ced57d7c7052ebcc4f0fa71be044ed583d31e7df9740c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74fee3a4f963660c08d355af804d58b6b4bb2761888cf9fa0c78856a476b4ba2e19b9c91fe76dd25d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5826621acb57a8220aa670b0843cd4cd710bb9d1c1a054f56497227bd4ab27df13f59404b84665a81;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda1d4b761f487f18dbe36e4382424cb25c897b06401040f338b0ab8545a6983a25bb9558f39d24c09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a1664d814d5eb2c51b97bf541917941b2d0a40765ea74946939a5e9f5a2808a6c10aeb6cee64fbde;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf82147dbfd0ca983cb03e3d94c083368341ffaf86df7cabd02bee73c6e9175cdd07d43298c7628d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3577cb15b2bccd7228acd5653d689b12720daf4cde56bab5895694d0fa7d11fb490a66265e7ef93da;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h711bb9518adcbd12d69b0ca819be4b0100faf713c79a65bbe0203ac1d223bf332259a579ece8dd459;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e15f1d85ad5b167537f1a8923eaf2dee7edd4d8a31579c75d69f7135b613273b667d18bcc9fc50a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he040cb7d00d80965d499e18aea482bb488622745b2e64a92defa749d96c36980d0e5b68161b826f8f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bcd2ec64ae03856c7ce3fc7c11e6eeb41554635e13ecd4a3f118948006f3db8fee046c41bb06034b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b2ddacf76b24e1fc6c269079b60d1b3ec60bf5938a719771c9edce4e608d001ad3baece81e7426bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36fa9924d58805898c4bee8a64417b12b4ca433e680ba474aaad876b9b074021e0b42f8f589e80ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a708fe6229f45791a8bbf473286419897677c504507eea70c101cbe0e4d3461ed7360f52475e94db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5619ffa34684ed67413cd0d8d2fddc69af94672d79a5878f805832bc97800bdfa6f1fbf073c4889b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h645d8427f5c36050ac29d9be3c5556d2a84e48a16e961d5675f2d4fbcfd74985aa593f780070b0822;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32bf431aec27b8c1c3cef0722d4209b112953b93d60e203973b4cf7086ded84926f4246758a97aec8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9a5bc4791149c464a92ce616914b643254746ef0e3fbadfe70098df9fdc99616f3fde1739ae029f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3ea809bb3cd0aa308380417cc99f73771973285aabb771c2b807a42de5fb799790abfabab96385e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h734169b3689211d80011084d187a13978dd3f86747a5ee0c91dfe734561a5d72f363a2fc9f9645d07;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65c895ddbe021b6a13d9ff05847097b799a110fce54b5f2e5d0d59ee595fb808fc6dfe74f67ab4096;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77c15800eec257cdcf88e4515f8d9be68c8085b742d6699fbb2dc97ebde38accfc4aae28a0b0235a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4406343b75aeed536bd36a5abb0ba8517ce5f80bfeecfd3bf2ea698cd16b920b2f77566774cdc67d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1bf58a09dcfa472179abf1c64e71e8429df5590e910f9ff512f9698d050158bea6bb4bd6e35917a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb7c38c25be766831f80780846f83b0a9e77d9965aa9875292171c5525c6748c8f165772e663efeb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc07cd1efedac18c07eb3e56a46d9c40a0def8abaf55c541d9fc7428665769cc5f032921182a32dbe9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd661082270dfb60665ccc68ceba117d2ceb33b058c65a4056a6a4b23fbae623e52aa73fab322aa60f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6253f8e3b3832d0f861192045a4dc3cad84651dd84c708afb16d64b084692decb97933b895a2d5f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36c31cae747838bad644335e43e1bcd9fca0e5948d0829b1b438870bf2a62ec9a0a5f79c1325573d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25752f443f2bab48cd8c72b6aa8eb497ecb566bc3c7bfa5c184a8d7b1744894f5605f82ebf94dc1ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd43d2a3707fb5b890592ee5584c303b99e7037424988ec566424102052a877d513a4cccb5290625e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0c894b44e1bca80b4640430b57cef51af2fb71fb8bd27e60a3101501b7821360c7a5c177df3d7cf0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3bf7a3beb7f5eef2561927ba7e6cdf1696431bc24b5c90c420522e40bdc918e06b702a9b6a71d3934;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb379f3066d7aaf4b1be64e92080fe6ade9be48492b12cc5b7523c363cdb95be0e72d2d3fde4153347;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8890d8435b4ef2a6f21c8f248f31a15ddc103481cd7f42f8c130788f813ff31b417ad88568d051417;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h570e83c67e38d543b19bad2c9a492472e1c78ab94376ac7ad35dff0de76f7fecda07aa84b1af0f2d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb44607a9e3adc70333e9f57961905d41c38215769fb22c4eba1af01180da99045d637864d9cfa495f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h785423cb206d6d0c8324d6080e5ab547d928f740741ab584aeac496b7f675376e751dff7f0be22a0a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb92b278235840723783dc36269ef91a2ca60403ecf50eb89b2a6feae560427a6dcdf24cb0dcad415b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef74afbdb245890f389cfbc2b634f76ece210b5fcb89dd377a93c4d6b637ea4ba32bdf0945dd8523e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5be9b5e6196b7ddbaaacf23c6c972a72bce101a03bc6b49bcbb219f8eeca46f95f94239ba4661e943;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c62a7fbdbbe167484c8cd51f9744087000d8dcfb97159413e4a162ca92d05037b4463aca7bcfa644;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87134cd7e3b3858e960cf10afdbcba638826a86760846a44f57f33c0b35e5b475912703ad5420f92b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e214a5284613332508dde51a91468e43ea1f8ae9894e9e5e02190931263edfe9461723b937dbff52;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c1dc7e68dfeeb82d03d2da66a22af43598c06a24212cbb5b8ac9a3f8d1a99db8c19aa5c34cc08ef9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e7af5e653ece26c37bdcae9bc225c67ee2b9dd55b17f35d6d881f95c3d9dcae0c647cdbd4c39d0b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc335cdc028b237f3f36da973cd475d61adb3d7cc1c62821e9b73c4e24bb2414f3bcd6c6a7338551c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb11c921cce5204501d9ed4e360a51b9cbb31551ba60d7e66e4514dc34d2d008cc9a6381006137e34c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3410ea96659f8861a8ad6af9f067ccaf671bea378caea08ce782091275d85697156aa8b97172c9e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7ecb9b008e655d5d9381550b1a0e862f5866a3ee2a621bfa97df04d6d2209248385b31b620849eff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d186c1ba5751444a7ba53a916c44d94481d70a5e506bcddb5b9977ae21bfca87af1faa4025206fb5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfee2201e461eaa3f3934411b4a5d3a1857af11cc935b8823fefaefb9bf7a0bd2ea697fdfc56b512b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15b774dd06c77f0328ac5dbde8573e2a05058ff55db5337c891842f4630e127ede2370ba5587dff59;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2100f9702da55cb539cb406a08021fc76fd8da7778233cd7525c706feaa068337cf89d4ca50e3a828;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15ea6b929748df0dd9f1b74ccc2c27c163ea5584f56ec9726a4b5f7af5c883cfac808aba949961fe8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd531f07170a9d52ca9f2319e9d18233234fc23d83e6cd141f89dd4ba370dcfa02f42a51aeff154eb9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4b809e5e596991821a09410704bf119860bf6bc9fecbc3ce5295b2910b332e3bc9282e309835a6cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2a5a9f3a61562ba991eedf82cb4a7889491de7cce090554e3b619823dc6e871ea0518d8588c35f1a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h225fbd507e78dc039a36cb84a4cad415c7d56f5e91d1f81fb809a264ffbe1075844bf08c2f68419ab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha74b949650ac74b9d8756d0d1df36d904bae586c8a358a06230e8c3a999f8400d36e199ebbd34bf25;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd89e06b11ebceb6f9c09941132714172b1cbe1b6c6a59321afacb5ad8d98446e9cd58449a427c7904;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h517a62abee00d160fe505ae994f0fa879637b0ada1382e356407faaa6dad0d3a917fb0f72f3fad732;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf284b2d1b7bf1d259323ce33336ea06484a474775596573a3fb187bb429f62f249cff78b09eb70b46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77da8463af3aa2cd3258d578355b4d1b6fab4a07a18fdf3efad504e9b1b0d89b1f5d5d647eb2d768d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha1c4d5d97e1f96863df9a1dce5dd57e8cfae0e8ef5c07a7d4b5562d000529305338e7fa6c4322fd5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44a15d31bf5fbb69cd85fa5b6c9dada84b00eb122a8ae2a87336ed067adac54432dbe23effeba386c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc38f62c14c963c3dd9ca28e86d5b5513ee50a24740f81fc90077d559bf56cb00ee7c1a111abcfac73;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h357c8f9258df48607e1ca4301b89a21313e45943c338ceebc4266119d172986f3304e8b289482b9a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd47711dafe7d09dd7214a879ee6e6d1bb2681454a35859d5a276765ab30a7b5134c082f8251ed46db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4cbdb3362405edf0081cdbbde7eb5bc8d613b90125072ea15662a2c082fee3b292cbf2cb019e4e42;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb992c8fa5b510828c5be8bf08c708c422f037434c0e4befb64c93c43583bfa1d3092fbcec12c7fb54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3eb7baa18f85ed8df2ec90a72715ba890b435a1d07caa39423a273dccba05cd18f2bee7875409a2b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d531f110540b22f389e37eb01b9427dba24e78051dd1fed15d6f8112bf4cd40ac4b92ad6822483f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he084e5287764a7dcd2193e140fa37bcc509beffbeef6f8a4e59505310b02016e0e9108875729c5011;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heddb4ccbe1f0954a8dfa216e15cc0dc6d67e60001d0f71eff99abf8b04ec5f2150c4994ea94ef9bec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha80a2414bf014b9c1a8eacd20e58e31f874782478cf2c05550b79bb7e712ce4fd967f3aba9526d571;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5002b90eae5e69b9d0f92d5bda8d4ba76f790d06cacf102cc0fc81651e7316e1a5b3266eab503e31e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39efee9aa8e0701bb7ec034be0d68288b3acfc5f6e7b2af9fe82cc7b4a85a9c74ac79c91968e662b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ca745d359f51636f9aa791a14d198d034619642c0cdc21c2260aabf29f184b154a3bc7ee161327db;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6d25021ada440983dd8f7b67f714b51eafa4f55bad88fb02ad9345e3df63b856ddaafb694130f690;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1d8c8750abbc5e9bafed2fe5bbd2d1f2af1c8cd009e4ae30dd4c7a9601a484e0801302bcdc1adc62;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82805e798a8073cfac342a03956921d4de91daee2ff2456b274e6ac07f92a593bb7a19d5440c3d89d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcec3a6712a70f3dc3987011a8fe1f042895abf09441cc8e56a67c86aaa5cfb644424861f601509636;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h947a2c92e8845555b89c05c77f9e792358c0105e4dc5fbaafdb33c233d56d781c5ca5378103c3097;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h106bbe93efa3c1b7c87337cea68f8f2aaac8793600436e7d6c991536d125a32fdfb382df688332163;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b3104bc8077e2d90d26138d3d7bffd7817b8fc8346ebe07ade06000d561b6bf1e7e10903fc6516ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c3e9a3bdf7ca6e45adf311b7ccac2a196b04f3721a56617fdcc72112a3822db6948d2abb8f652fe6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habe5b8ba6fc24e6c81484834cd18ee4988c5e7a3e3bfae95e5056bae89d34954d88b5fe99605ad06d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80d2311205e173d758799a40d34e62447bbe7095450ca75d13d40807046bd2ecaf72dbd2f7483eba0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he191803a64c65fdb1a610ef4d0d5b1a730cabe99344b95c3ba50df4d8ff4806ffad2a9fab4be3a585;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h349b758d4a570044b80e326f0e6ff4c434c3c3c66ed70b2ceaf827440cc44fce53413a438bb893ea6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f69c004d8a2567ad3a6a3ed050684a3c7b7a30dab1b29e57ae7391ed390bb424e851c943a0cd038e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc2ff06bfafff7ad3eab1dc9ab529623711ea08608abf5e97e940593db7a38bf7ef16c8ebffbd5dd5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h971a2cdbf464819e0d9e711f3dcfae5ea962b82243e8c1146d813fe9d7331825ca47a0f50e602d731;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7de776b2b7962e6a67d7526bafd0836619cd8f2faf72ea38141a22f941600caeae0c26fcf32167c6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71b2f4049fa5176e073aca179410e2580de1efeea2cda0a6ccae7de225f6ea5f2bf41a14e9e240812;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a4f4afb849a68d30db999b57d5e0e0c0d6be249efb2483776bdd4915ca3f64cba1e2faf36f6e0a0a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f90123dfa5fdabf7fe04613c1c9d046cb78fc6fa5fcf5d85866597fc6add8fa4408bd16f977b9894;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86de5f8a24b8efdccf07d8078d98aca51f002c98bb1e03673d7519493d68d66c6d65272797c38589d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h271c944f0d6f8614e8c50fd3166a08486adf657f1c786de267064a4e7ded26eadb9bdd3c244fb02e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c7e7c86bb0143b7d8e489367f227ed15bed434edee9b767c3cd9cba62323c73872e9ab40739b93f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65c61a65c5d19d582da243ad20ffc6181016abbf4303b79cba2ee4bd61f0037d2f984bad9704247e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94ff9231933432f3d6abab01aadde47f392863c72ff4f12851a90bccb5b7a301968b822ee786b9190;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66debde71ea4277c7d0a31607418c3859d12d6f01e60b4a243e1cb389f74d116520d0a8864158d7c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h497450cdc7096e8549b736d441f9117b614752e0f59a83ca318d531033682f225e0795e1536afb4f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4545dd7f792c567960205689fc1a5204c903d59c6495b3c30d4469c359473c463f0866fc8be1e998;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h872851fcc0fa38362e0c9311f3a50c5b718781e837e67d46932b4adb1c8c24af6c60a9009f597411b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1efbe2df6825c5a4f7c6395007f27f00ab03171101c56e136abb92bd9e26e5e9d4250988961f91e0d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99f1dea7f6e2e7663babe6eed24b2108b6a73cb3598070c5014d7a959aa90ffbec9c4da0202cc4846;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29b8b1605698281f425b38f386ef1075d33f01160dd81524f9278ee23a7f9d493a9859ddc39a2a778;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f22366095aa8045a1c7aff5e59421b992fd6fc4547f6c99a2cd947e7ff81cabbbe23cb8ece3fd0c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5595a218809d103653491f7c2d27b7e8f266b8d9354dc4c5592ba7ed7a04badc6da043ca7ce67f866;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e3b384ddae2e4bff58ffa6cef20b81cb12d882b475d9dcadd8202ba26ca947188625cf24dd40fc6d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd66098004306002bd7b7655cfa69f5d44e2b71f556a9fcd49b269c9282576464b67581ab066a1bf3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35c22b686450527cb6b7bd00571abe43bdc324d0785e6a310932c6f824cf23b24a7164930b739ff0a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3895250ad6905cee4953fcf17710c3bf5b832d93e5d464db7ef870e37333e4d15e7a61401acc57846;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9fa5dbebfe8e1b32153d2ae0775e58cd1303f64a6eb9f9aa405e585f2873c01e2fbc5569bf0100ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93f4e22d2863bcb1dd67cecd73c0582a8e00bfeeb80b1a42d0452ee6984a94c3071415c6479722fdd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h749413b5b6d23808a31e2fe86a983dba1da09d11d0dae75d58bec602f7b4071d399b3e97ba755b118;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fde560e853f53db40e8acddee730022a2ca19580502f7b4a3e1b10fd0e37cf71576a5965225ce703;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d4acdb926ff8e15d82022853160969dc636738f99f33ef8ac0d3784c0e02142de5d91d97cda65bf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf93073ad2854812ba8a3f6f9479cc75afd9e348d66273b7d7889e5ae80e6ac5856fcb04e3ffdf3d8d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62c8d9b6a2f5dacc7236ca31384fd50ebe62f5e21a2c222f95c791c1b29b25bcfa385b04f7c0c041f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcbdf995fe7a7c8b4d2814f876760b9a5fb34205a11050c77fc49627a3aa9be56b4c1359527a82b246;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf620b4b6ce21cc1df466b6f18203023176cba433a45043132626cbd6cd4222dc1e3112f6898e9fe13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cf35aa1e651fda723563c1e7d68c5aa055379e802f83899b2533b8886b8edafeb0113af1da83b317;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h132ac85e0322e23484c95412d17694a911fd4180dd60946bfc1bc9f488beee03a938ed9ba680ff6b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h334749f27daa0ea9155bd4e4a9ea842b84f4548cd6156628edf8831954dccb9e01f01f9c275ac9664;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8e2f28f122bbc6dc6c8ab929b2328247a64a34f16e3b798d0db0033abc44baa495df684f09cc80d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53d1aa90b4080a1d9b5b439c21c6f1c72d3206309e1bc54af913cca7e80ff7f373925d1f701afe0c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc26d13d5613bd6a9091b05806e2abb0d7ca3eaf875146b715d64d97863022bb02f118bc505290fbe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4a89033b1342931fc16e13659ab04664db1a3de01e467c3bfb6c80741900bb3e9be656c6b41fd633;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7b77c9d14d000cb03d65e40271fb449e5113e83a97bd1091d242c36b403332a55892334471137346;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b2a2fee22321c2e88f7dd916018f27297dfb0eb43c06edeaf6afa515886d8a77202b12673db41910;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88757d52ec59b590cc5a1ff6415f42328ae5327f445f2a857cbf7e02c39d40cb3c3ded448ae8914a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h622fc378efbb9da992ce5166e6a8469a536b37b07f476f90a0dfb31676ffdc29fd6d4ae132fe21be2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h124d62d33f767e44a3cedff3af9da469c39981c6a8f2c02f9fa73f8ca51eaa87a0d744c9bc1b93f3d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5bca5d4e923d8e2a002fb59e1e2914e0775df8778eb0c3c20ad94cd93b1873715c336c8b59431360a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd51ffe5fd043e79919a737e1ce59b6e8ad2a27923b16cff16f5affec5743f9253b2bee7567ef308a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc12fff5ac04d6247db6600667c44ee8f0d4e610b547ba558d242671902a0cf312e44c2edb9fb69bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd57cc57c400fd309fdf238aaa9bacf0c33a4448b626d3fa88544a7a03c330821e6ed6d184ae33f57d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4877fe3157a64e6b5495db3fbaca0cdb9165b632d268686f701ed2e7c9a2c64482c263a49af0ea75;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haac40899bf25e56b9c40679c42df81073d6c62f88b2eda374949e84675a9e7321a448bda785b9ff10;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3c5efc5f67c3f01e2c5bbc4e286c5015a4537fab0c5e342da51914370fa9cd3a164b476b7cab244a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2971ffb510af397d0e61540c18b8b147208079895f76fb1791eaa0d5583d852a26ed6f59105c6cc6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e3288079a3b5ac3aa2e03eefa619edea379c2fcac1a1eaf88c29585cfd2556ec0d78f19d220aa598;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22deaf37e2974a66ffdb20837279c03af7424158069ab2ea38db682fb9562b9a4efa0bdfecd521924;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9b999d8d23a61e3502f6c72ef147b85093140848ddc65372d128ea4388a7a706fd00ccc63ddf56c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e9159649df4a552e2cb309540a0ffb6260ab8a58a0a2c24d738860bcba3bff3b0dc34f6e516f9772;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebdbfc45900375202e19bbe886ea038db8c99aedc4014e90d181f412cc8fc3fb33a4962bbaa74ff47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b8b145cc49ca01d034b20625a655a2455afe4ee62db577ecf7c3107e2464ba28ba176ced03faf59b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heeed67a88dfc32fa642e28dc68c41b19eb3d72009ba51c93d504fe0d33070fa7b1f5ee1328423f4f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93f04157bbc4b8b753e255c6bebca7fcbe5f21b1b2c3ef5befbe83da8e9898c853424625990f5f056;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5d7d2ab4e8680b12ba5e649f7f9be9070776710dd279e1085e102ee9e2776bec74cec283701410eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h585d51116705da3dc60ca778242e595474b15116cdd627a86388d43031f2279645243915acd07ba55;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa632115fd90fa57714032619a9025b521824d3fac92bff3e5cd46dfef738cfdefee15a246c0a1730;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd23df7ed37dfcde20c2592179e9ceaccba44701a554f4c61c6090647c47ac24da5eb3347b46e3fdb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45002aaf89d02986ad20f2d7edafd2f76ea1af7a69ae5c05a5ba99c0f4c9399ed553c312ba6c5b6d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b8780c160fc903558e95f80c74eb4084628451a290217f8b276bee682b1b75b8508ce94ea8706233;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30d718b4368a76651a3175b51d0f95a3e770c1a60c5f229d707caa037e1f26faa8709eb6825850fe7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f1ad2d94d10dd7864e1fec11042d271eb50b75c3025f888d988253355f3ad867eed62e94730a59d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20699101ded9fb0a16b54b83c0099e2b5658d8162c2154f213c5e7885f556c49417fea1e09bb2ecd0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haca9f3e5ca98d3a4f94d6805eefade2df87539c599f125ef6e6a8657598579334a8c9f45c58e8351a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d09bb41ae7ae5f3dccc2945e9d71268429bd856176cc990732a4623e6a2e9ca64d5f996f755878c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h601dacc8caa87decc61294ed3a8520403b180c4588d6d967c8f700fd2e5eafe77f7182264b6f28ee4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd88647b7a4ff1fef36674c168dd3408c6d5df03f840c6fe07d63fad3e57904485d78cdac2956ba92f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50c27381d7b6cae18d4ac0645263ebd8f76cecc09b33deb11699001606eb010590947e17601aa6070;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa4fcf69945a9eb3e43b33764867bd5936c353e00338498d064295190ef39efb3af5773ddfcfd44fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf48897926f0281326d3ce1a89cbd2f5944dab3aecf685a8e6ee07b6b48a52659e6bf9ecaffbc62baa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb10a65e8a6be3180cfc8b66e8a289402f083f47df3174b4fe0e2d212bb0299cd868e4acbd70682e27;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97429077ccd5c4928a0f1baa24e157e771c566c9768c4e30749794239688fc54393af7b0ed29bfcb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50ac8c88349d5e7ae5688627a40dd04c70cfa33376c2c02722df4009f3cfd61518c62626f8018f534;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c2fe4ba61b70e2e78ba8be387cd2560d95dd30d6fa97b7f46cc3c3bb535d66f11189b7c01162b1d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ceac3703af0cf710b38f23c90e3af934cb511ffc63cdbd0487ee91da51401adaebe5f5e8747fadab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc381023083e9b7dc7ed6feecef021821684a222dcb6022235510b70fa5b1e0a5011117b2fb28fb4fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha588177cf6d0edf234ba45600acce8583561790f3038aa85e2d03340deba47f6c4aa2f2d1b783b83;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h486081ddb34ddd8b513f51df3489e8fdabac7dd9e01935ebac77fe622cd334ab71a166f5ebeaea9a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6aeb154013a428d2390eaa113c515d10b951415114e35ff6fde37141d882218b11ac4eab2fda57547;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbaab3648f8a7d41cd593379517bd8c02d6d79db7fe1c97c4f11cd0192b7bc60ec2be3e8138f2ef73b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6cf146009a1e4369f2814bf851e7f63281ab39a73ffb47af349eb7c4cfc473de5628529f218be8403;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd7d84d15102c56ef10c8120c096fdff6dfc91bfe1e202340b91359672aae33e06db5ae362fb6a187;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcba10cdc7f2c3b7c005f81bcc3105124c3f760c1bcd5fb8046c7df0c4455afb85633ff95584928a65;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc09474be0553cddd91575156de96b46f55437d6001701eb33aa796204a779a27f09ea5c2892fa7d08;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h846b1e6173fd4ecf8d5e73a28b11da0c81de69711adac6f60030d61e2876f23575cabbab0748e9e18;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec928721045c851b5d09b99b17bd11764a33ca6a9adb21e4319df6a65ab1f3ba665c2ee2cf19fb0f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7993c0404382d96a7695570e06c9023e24113432816c0a76361d5cc77a91d1cc13abd3da9636abf5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd561c258cafbe1eca007a0b3e9c7ba899b63f356eb1627ff62f47b409e2a9ed7e23ca6fe3031f020f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2e9f96be4993391992b1b27080a67cd173310374c2bf7724a41a3b46391cb4b63bca4eed15722044;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf41c66a85b13afaa0ad5df1df9869ea7e29973b6edf153fc236f655785fff84cd9d8718bad6e0f6c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec94e86eba4f9057139b6d2a6f60b781b9622ff38c368b4fcd62eff52264b5bb8800b3f2924a8f7a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h283f8320ffa17689f899527f60a1ab04c9440f2d56f99e7e3474102e1d66b9c97759855b12b448517;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb5b30978ef014beaa7f99559317d2d8110bac6b8f4513cfe59ea33a185c442faa69b12086cd7ebfc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1f334eeaae4bdac62c61a04590c22d9e303339829b8d700795e031a70f34817c8d7786f75ba05e8d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2798d94afc1ded58affc0984333c87ec6fec44c92fbc1f4e66c851e7486eb28c9e3566de258cadbe9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4e1db087285c5c336eebda761cd6cf68ef7464c1328687251bb83d7f69a693a97c886dda6df04bca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8437994f60c3ce363764000dd58be55948a661be6b47c7552d2c902cb8c7844219ea76dbb930c79fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f8c75da9141aad7f82205c2daea373fa54f48c7645b2a240d24e989478e7c9fd312eb66c4dd8fac0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8044a383e671a406b8c669f9d7df254655c2d6bad2e277d6105f39f0b3029097c219d7d2aba91dd43;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3d6ef3c6eaff78ef94d8fda428f270db4c0a2c04ec4c384b38783859df0531dc25c9b8710508385e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h294bd524e38b4f90ec693e2046a8d2e3379e9393fecb3775d31f4bbd2e6224c7c719f1da3c6c43f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habeb98396889664ab9b71172a4e20b2639b48027367b69be3ff00b2cbc72cd5bcd298ec05f7f77339;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d381a5e74bd07fdb5b75134e42d350cc717115a024d4561c995bb4e52501eece01024f5d7727f452;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5173a3216e381b54acf308ff1ad2233d7c4ac41b484ecdd9a1638ea37ea66faa0b181ec49c6d7c83;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb72871bed483dad9ac5b92bdf699ae9dcbde401d72be98084a37e292ed1c1b8c01eccf1a8164c7d4f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1bcfd2465f29e0d9179a2dbabbe878dbcbd2101e7ca4a870c7b66309cf2839e2f047d50e5ff09d349;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3b8cce5876c3550ebee90d22a56fd27f63a1a17c0c5408766b4455ee0f376b625f5fb7c479af39e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he040a4e1f29e92f3f46bd6143fcb86c979de75beae785008137244cb19ac3fe652a2f8dd4b7d799f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57ba57441d78f9ca22c26fe0fdcf6377263840e18afa4a95f38b0cc1daf4e9c4b2901e20210131b04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f2246c0cc3391929242ec1fd507f43ddf80641e30ad07a6267de37c7a2464ce73c994d89963cc2e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5debbe580707d41290532970bf72b5b328b7589b71db7439e73d16909d91bbc0cf6a12edc36d36790;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed468bad021f3e39f801d091f1ea266e3bc01ed451da3497a7a620ae49cd2330f74778f5dbaa0e106;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a3239af21b29d552318e4003c1f427bf8a0c4a2c244ce9f908da065fb69bba2222146128bb7f654f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d2a0e4e3329a7e4f8653f4580346cc288db334b4731ba9838b6f55a13b95133fb6f7b1807d74c8ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h105b473bf15806c15287adb823dc985559c992064e4c3d91c2b14b3f5584a4462c43476d092bc4731;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11985763de7a1925edf691b7f8611444627c12e0ef88eebad148fb7560df6171a1058fe3678d6a7c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0774ad77199398ef1be2e3d2e9ef05b193d548308e61c3be9e6c842a7d35468ab4496e57f23bfadc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f3e8ea2356ef4bd9184e391b845fe3b55ad7d20395e16124127671ad74e5ddc47845d21a21803fb8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28b52588fccb2b66d669e205794e1025972fd6a34f265e29191a397e0565463338324457e6275aa09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e2e7f7a878ff2e7d4fc95155031c5b317261a4895048e4371775a57f48a17929cd6d9a9fc55c1177;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea8e64f3f9ddb3b9dd4ba48c8977b0dfed3af2353c75bfec274c3fc360fb20d65d961270e1f488a37;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36589ccb832f3894c000c65cdde9bc9545fce273925d0b6742ac87a571aaa056d95da8311ceee21a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc8fc67492ed6ede6c620da625999bf34e589ac72f13d889488df60f6f53eb9eda060a33301cb53e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6549b35fdb5806f151a3dccfadf2e19864c71b4f5161a5b7fecd8a360ca0c9f7134ce20a5a7da30bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69be2ef23c50e2c2e47be1920aed9b94d184e185988533eac48e1aac6e5f9dc126ea4b362b07b46ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97705b34bc3f34f7a9753a12921e3c16c6d20b62fc90e88ed4a22f4470f57790ac27fec060dee2bbe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1dcc5887ebafaf7324977db481eb779d4a1dcbafd138cb8fa3af3d7b1769e38837b54b8c889e80d58;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87da94558a0ed8e5088f0e00be987d96480335d99f32cb514a6352433a381837cbbb2c9fa50e2f573;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb63edab0112d970fc779ca6f8900306bad6ee31348fabbb716e6ff3a9b9a14c29c0286f2641f35a19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he97d0f9d3fbdc723d86593e80813ee9bf7b13427d9c03f0af415b66ee35d042f24a092d54b645b0cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88aec6b3c2f6f5843b59ac5c7bbd8fec6d71f8e0cf1fa342a84ba9b45775820008d031f62c4aa689d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he679d2ff4afc7276da160c04eb7d870061dc01e7ce8efacce64f3779a41195113b9b71562cea46e20;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d86341a40c61b1564e95c57ed69dd73870431b6c967defaccd6902c5bd0511a7b0d0f7602a4b6d2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ce6690fcee73b57ce069f4cc64e89bc10decbe4bffc9c94afcf79fcea143663c1fbe5c76e3589315;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4ee183124b7e39dcef40502ca9ee542444db91b07276d6e22dcb314677c2ca664ea14c7757325cb41;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habdacdbabfb8509047429ba7f4faac5c6bcda37c055845d1717b73f03c5b08290e6226c1c82a3035f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d22a7cdf8036c6d54d76439c979c0813cc280b8dff5af03cdddfd24188f98237e4cc95112c0a038e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42ffd9232e5783eed03a70f9c17998500a4d456982c58f80065f99010d63a5e2bd5e42c44184be8e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bab32981d982655beef7841415d9b1025c5f0f73e42a476045857b70c82013cb6a85bab1b322a212;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba14f25bf684736e36b78385a3c3adcaedd5ec8ffdf91d9687ad4b33b8782e469d7d872dbac8b0c4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2409f7ced97112647d8568c60b7d1ee03326c0c3a0bd645f76eee4ed8a49f58b0e48991606190d1b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddd31f06852368038054b86d90924a2db9a230d0912997aa495b32971886fa5037453770201f66e94;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc09216c6e618decabaf40fdf4c9e3a243b0cf4cb6850f6aa1ed428a0aaa0721d08ff6df475b6ac22c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffb4bc147fc860d2a509b258035d663cd63bebd7b3048bcb37fb37b71d195ab3ff1cd3654bd719c19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fcf6578c40b247dc5c43b284f3562a4438ff22a311c0389796610c7794be7a7aeb9fd87a388072ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a5007baca608bb52f82c8597f180b61db0976d6c0950218533f6c5eea0ee3fec355ab54d5c59976e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h387d65a2f993256bdfed67bf614f91718b6b401218c359b5f1c1e2963f27a73d614c7168f4549c9e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1b7e24311277a7171e86c69a31c251e2768b9429dc2150db1cafe65330fe89ceed354d6f380f7a5c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1658d8cf614e349ac2f8938a0cc5b6eefecadf3c07b3d589621f600609114a263011e223319cb5cbb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4fb09b673410c29a3fd5b9a230c24ecd2455eadc20aaf43e55e0aae5380e19db51f18bd94c8cf013;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2471706a390b6864206c1aa60dd66443760e37c94f9e331009bfc92b460c423a35fd44d5c3842c99;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce607c1e5661824c42616ea71f16ff9aefc3caaccdac978852150b2c999dc102a29b8e8734d5b1217;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h32f83a22d66a2602f9ab72a05980dde83fd869e06dd85f2ef6749e10807e6299d7ba33419e238e46e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45324db05b74a7ad2cd9b8baa11901a2a67883e0c26f4b4c600a62c725d52175a1d732f18e61c6105;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h445efac35d296e6da3ff89870ca6b498d762c699be4de87d6859e9e0df3f3eafe88ccabb4c5e1e8f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb607b07cbb2feab3893578636993819f03fe63dae0324e10b092dd5a12b61f002b910a0d2deee75c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf83ee55d7e3987c7953af34038e279129c3e0e41dec686ab5fd94c71ed0c36f19ce9c850f51e68af1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h509bc6b476dd532822f55df8c14cf73e00757edc97ce881f94f7a6e30db520623075873b768ecc0a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf642efeeca66ed0290115ddd5c3fc8fb9962f474a6f14fee3fe8744d3d137bec4e17a66b2b1507890;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c04036e3f989f7cdcaa272266f2fdffe4ccd20d4b43ffbb8dcaa1c034f08ba6af8b5c56a72219cd4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ce497063f96112229d618d5356e9bbe6db280e8774f6207020b91d8026c71045479e47d34b45e883;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbadceaf824b9101b0dbad91c6069a50f4da1a1b70c2b380de2b6c84c35fa03d81f75c08d08b2ec31b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7ae5e6a5e936c1470ed2710155b00334271dc45ed3a757699bc0f631e33f20c9ea2d13ea4a018db6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2e4653e838227e6d84d17336dfff51078e2e2a2df041ca981fb81c5c61d4b0a891a51655bed66db8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h625f021bb48abc49c1cc7601c154a532b92c1b23d61fc7dc17c4d2722b3f510fd711295671262976f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8703358fd1d27393089f80bd7c0157bde986f92c8c612c9805707c7f40506f25056dedbadee8f147;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he57abb317a8243ae772536f40ee39a31c0eae5cbdd42036a5243c8708a44b04cca00b9e587db1aa4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5809acc1e1648b0d2be87c4e3c23f31feb8e3432ee6b4eeb738d52f4b6cb6721d95a03515d69cab98;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5d7f7d59285ff73eeaae30ad52e5c86b803ad0c1da5e8143c8bfa26f2b8f43a04b9f160e9427b742;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fe6d44a54c59d77904ec99c4be5aa29930fb726a63daf7933ec86f2c448e07ac4abd3bdd23379b82;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7cf35cd449534f3ab7d7c436beb9f14c416f68952e8530a1a7a38fcbb790f0b47f2a99b9631e1113;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca80c7942cb6ad679b01a6c73e11c9a2931e0fa1a12cad38b8e1bd78eb20b47e8a0ee6cee404fa1d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87a00781ffe63729176717ef9eea55f33d8d46e429a059cbda6ce9c2805e941649d295788d93b3265;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h372bf457abdf8ad428c0aaabd03f3bff779238aeb9fe2a84cc1d46994ac7aee3883734694ccd3987b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9f9369379b161bdbceb055e57273bb44e1e6fe99cf39b5203983d79b6bf9180eb84979eeeaef41a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a8dc3ae659421ec95c6abade19ec8f4aa4584df81d34c90e020af67409095ef71a0f30365707f68;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d92c66f5155e70ac0c0960483af16788194078a912de3ebc8ed9e430c8924d0e019410a5c90be78a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5cd793f367d51fe1bd9b5918b308ab5e33f2d447b2322e65c060f93437548367db1a77ad95599f2c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8868eff257b01b5b6312dcc84898939d85450e675b86f4b8b16aa168c48dc5ba6458fad887bef6dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he3b633f8d574f80a836616387e5eb475d80ac633646f2d82771c1cc06e64f8b376b80e826cf998b29;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2e76ccb4dbc4e4677bf81040d397dd00d5e5c35ba672f08d180d1ee474479419025bc71f26b5a399;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4318b95d1e02afbe32fcd257bf61a0f3c84efda33f652fbd99f544215d03318de5b41a659e10dad7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h746a7738f038aff51b1b5228eb24e4973e509fbcff325da253a85a03f1e574c8cad45a9de23bf7195;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf5f42a7c55d9f9755c1513ef6e00dff9e1f91f38436d492f5eec0cc1d69102152c3dc22c1b088db0c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he88d19b51abd6ee79e085b8b136c8eb29c8273cf7c69a52c8fce94beab4dd1a497ac6e60b9c3bb855;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb27cfb8ee3964ff57d4b8acef0466b612da147717496558dce8e82331641494e6b8a6a3edbb67f543;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31c735087cf5787e5d0478c61c80cd19ee024600b5b84c17a620a9cb2132bf6f7a9b3aa382ce7e159;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c51bfb17c27dd652edd2b4c944be045070ca430688ff327a83a165315e16c4b296fc307f5cd19ce5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7e2ee105843e41ed1bf53c3c3efb9af45b7454125a8199a19dbfc9247cfd9386e147296f6b6bbfb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7572074692e4b75f749a8c3b78c61552557aa031e5150ebcc72273a302d0f4f48535e669901dd5d5e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h836e006b34ebc6a75acde2f0fd2940e219de8069e37af6dba91adde25d4daf89b66918c49c5ccdc16;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h513fb3ff83245318e0f3b9f4bdbdf823297dd59b28b6efed89ac45e48a6d82d7e0f4d02a82cb2a1a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6b43a093f49a119a899763fab206193991b8db068de0e4861579fa2a882186bcc2f1f4829ec05010;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba1e6b96ae5f86794670fe1352be830832cbc44283533a5523feb1b24795db36bef541bca96561c09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f3955a886fb2e220b9338697ace9273e0da8ea5445eb5980b168808980ed89404ac180cf1fe5bb11;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4197c4833292cf70b594e39295670e6c2b0f43d868617266a21ac77743d1c845d796b6408c30b8c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h623ec1b1863d5b960e60c236b6236aed6c332a27bc1bd03cb512571afc422995f96743b2083d7e1e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he66926d083b1760a1221149938978de8cb45c99a92763eb44705a5f01074fa1a4eee2656503fe1525;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h653f84c261c208c0211178d80d6cfb969257f6c5b07e638dd38f4f1e8f0aa00e487648de68bd11dbc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h415dad0cb743d9c5a4d465a77972894431e424d9d012c233416feeeb4f158a6bc5eb83cc6103ba5e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a07531a9703af9e3d51bd970be5a0b10dce7d277f0c3f9ddca8c60b55b4e9aafe6e628d18fdc4522;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h694911bd63d7dcc304035b6865480382859e5e21004504a17a7e1fe13d708f1f3758222bb6aa3675;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9039af53751c463ff7ebdaea02f0a67c5864f14f0e9f803b6a523c05fcc239963a0256473b1b00103;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ee2cc0cad53c5597a92e1f5c4131cceaa179affc4946c45350c9d83966736baffff7a8e1df665054;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc75064e2791e2720a7e535726e91d9c01e07349144840c32fb80694a6e481631ee62cb36e23333f16;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h552df1f5b7549bbd110aacd2cb327f2d04742ea8b0cc3c41db2cd085ac6ed97c1c3eb2b3a9f79a893;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e5d5439836f363303fa2db8cc38c877f2b2b2f99c1af07e0f39b3bbdf623d8f1251a26b6639a61c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h473756e30041b522113b2d5c7983144b613fb008ef2564c35c0c81fe0e500ebefb19146438643a162;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2c785d4517111b1e35fceb7550bcb591bee620e5166670ef6a905f652d6e71c0f98acb02bc252721;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bbf17ed923f4cb8a8aee2f8fffba1357254dd10d63fd66b8c23c49613536b70bfddf77db4045b390;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77ed101da12925901b5d181cc7d586060e410b226ff7ebc47eee17019fefa78ccfff22fbb93083e5f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h51ff799abf51848705e220d78c9238831a441f7790c92ceba485aa4a6a2e7e1cb075f6d02cd24cdb7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1af2cb4eaa5666972d04db41ee7278b653ce0f259f8489a0dce7e29c118ae2498b1165086b5736dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dc3a8eab15f56907fa42d4327e6025c556ae567983b8a66691015bafa9b6bc3b10ec639f084acb2f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9aed3e6110d2d60d994799752c3f2878f2cf20278560d85c9a22587060cfe9961367aa3c3ca6e6bd5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha303d45473e1e00f603d08c43b46aaaa0b59f07646ebbfed3094560c8700f3a678b38a6e30398ea54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5ca38c25e02d827f732017410c6747ea7eca3c6f94883016a79a505555b211ee1d9fcc90ded48ebd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ac428c7ddd97f98f0fb06191827ebed7791bfd24962870c49d7aac8e240855f2fc6013e866377a32;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b7346c7620584a7165bd37d60ec91fc5d78d044b37d1a826ae2722b77f3cf5589f9d2574455df977;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80b17a94cdfccb873f94ba7d27f691602df764a5d92b4e29fcdb60b892dd7c5e5a7359a91d8526fad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71c24caa0457f4309e1f8c1fa2a73df4a89252cab1e9c196841369059a3b84b3bea1907366b87c366;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd17370bc59afed22a26c2d934df5b1534b9cdf9df068edd14a0862cfe09f66e8c234e33dd2259991d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2d303a6c80762a3ab8c1c58a6b04321c830b8670a0fcacadcd280742b8ca71c0270769cbbb896d25;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3686aa6be334e3db4f350804491a4e515b1da1840abe2ad58cb100b415cbb514eb783acb56090b9a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71857251eec80c6b440de0513c7f9c813e56be9bb82dad59fbb4011e0e464ceb68f6adc92718e61c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53811e8e08d1edc2431762818f59dd2a8ad5e93fb341bff557d940d8fdc249272fc5a8b5eefbc4324;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ea294a88414539275c53326738146cb840f03ccd9859c9cba4e52995670b744aa3793b419cb990fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a3f7620f56590e003e8c37bde3909469e51d00ce06d98e8271385b53aac52e739e688f3a2630361c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha345c687e958aec8bf8d30375fa0f26ec45c02ba74f13f7a6a66d8913fdf1b94854c4a88c51f4bc8e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a166d2271f804879363c3bdd6d84bfaf7432efd79ec850fa124fb872ad9359b89982361295cc1420;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74b925073db72f0067824485f6be0b3f4b0ad4cb8fdcf34c6d75ce93a12a929f7bd59a00a6afc3347;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23ccf47bd8b81f95cd53722f12684714c45d0f9b60e08bfd40a678d384ef2dcc31f4f6edc0ca372f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c4cc8a417c146f07c299666e4eac6c89e0f260a0513427439f5edd4ee481d9dafeaebaa0e8ecb9a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef683f88976bb930ba4e12bcc903f9865eff3a7bb272704c1dfe5a28bb3e17cbe9ff61f19c7638654;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc98c551cb386714ed9ffe6b495899715dd1c9045775f01d0f8be173df4b609955205b23497a3e8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7d4677db54d9aee0bafe4a3fc9fc519ea844b8936dd071a358e30c8da28bdef4c9bce7248e626202;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6546619c777652bcbb5c6e4137ed6785d9627056df02e48568304bc4675badc3fb2c62390c19690e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2010842c4cf62ba3b448facecde1e251a1efe5ddf47715661ed30553c625d0c587d5e2214884513ab;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b6285b6e633a971e99e28643e3f7ff7e612dcf76d5d7e7740bafbaded1fd81e49625b665fc040a5b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde54878b14d717dfce48adef62339768dff9180d810a2b2a2cbb4a77a9abd5e96e969489847f900dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97db7a13ccbf1ed2570f14338e30911c0c3eebdc210c7c8cdb298f7a3767a66ccce03e43714da9000;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0a67d8ede5c4bf8a0de9ed2ffb739a5c79af59087867600b07131313c7663df01e6accf48fdd3dc4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b457ff329b77ed0edc27a5ad616607726f10ff00c722c4956446507eeddea8407fe6367fd94061ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b552e3674932ae3e6a7346a333ac55dfe3da3655a5c317943f8b8a67cbf39af1710e8022741dca6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2855dba10a31f2407fa62ec6596d18fc86f45aa87aeafdd5e695809284940ae1d027adf8c75088411;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h447776bbcfd2550cbb258689559a8f54c43de28edf8ae7c67204f208755cea2f5c98a8a70f8f23222;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97593edace11206fd7c173fc7e0dc49545557bb90dd1360253fef6998ce3969d8ec90d91207475e5c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4757b098fbbecd4b1c2d364224a26409700ae6d622a8589702d9c3cdc4440f7354d31a573db6f0a23;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaa8051b220542a5b71ad6e4e64eee8db05f46b2d9f6d5c6dee3ffdeb6da9f4ed6f59ee173fcb00c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ed51ac8b214add7d9c16fe193e90029b1f6cc9beb3df6a1cc3177e8773c0e76dc47bec1bedec4bd4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86e60d22bf2ba42003af4e043ff1c8bd19b18f819e2f285debce0901806acffff09deec9d1f1bc56d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94d4a9d45f9d7113114ff689e80cbdb108e3dd16e3d3ded94da6fa559f45d965a36dd8943a48c6f45;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf74b11c28e9d6c0d5b474958fb05a288879b9d3fbffae9f9ab7622c19a4c3a3f3fe7ef7c2a1e5fd0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7da935442841cdf453b171d724af4cc3f4e798b4d83b702c3694bb35fd7ba9f328c9fcf48325b137a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e7058a524b0a2b6227a341d6cffe9450728bead4828b7776f69b1bf0a6a0de05221874df5fbed990;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91153510c007eaf3f2b72505070f36eb1d13e357cfaa97d4c84975f83a989fd65e392e01dc5b17018;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bb1b49857f821a70e668ee7f01b6e88f9619de7e3476b718e638e4da4edd0f65d480e9db7e445789;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5130fa6ee9f98dec7efa007a55511e655acb0402f225dc76c2b87876acaf339722f9bb102127f3186;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ba6971b8b9cf42247f7c046160782f5094db301c75982a827b3983c0e36fdaa279e2235e44950213;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45ae5e930a61319b18090e04c4597481c37474ed1639c075bff2c7f20560746d1cd403960b42100c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36ab46a508e2d8d4a761ee017ced6604a0e385ca4fccdfe53eaca892fe7ef0e6f246b166c7f8affc6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcde8df2b93fc38af60cf58e2a95a134455eda75d03b31bce768681b4d1a29ceb27aac22ddaec6f6c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41af90ecf0151882f5696720b33a7691295e15a9ff08207cfbd601d98a52fe5dc39bbbe6dbbd47b9c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha836d55234bd8f8340af918050314231879250cc509d87c17ddde62667477fd7cac257e334b33e45d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a4bf61c2fe3dd5a411ef6d25d1e0e8ca4f8bd8ca3b41c5735c2ffa2a2a719e8fe3cf56cfefa70e4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa9b2daef3945c583e6aadb9073f5dd3a58607af33afaca30df39cbc1d44d5040624d5772e5487db5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6ce685ae7765a66d82b85b1f95fc7f810bc1cbc187b7e10a01ff6532f01889dfb4c8a9a3510fdb26;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2bb5ef689017a666491319d6966bffbaa040a9f5a3eb67aa5671fe488875810bf02cbbc8207b683c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h226f62883c1063cc7b65bde72bcd93950cf142e92b1a3bad5d78b9d5f253c3d7c0f4f4996b8a822cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6e2a039e00dc6fb82e67687fe3bcf289b5e92242e3053934beb21a35300d22971772932b99de0c25;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ea0547b2bdd38715a78956dbe9d2ba4014d19ea197cb309f6d75084faa8f781426eea90497beeab8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4af991c6c9e75aba952f33745b83ac52261e0133b4917a85a3946fce4f88d266bb00abbf0fa2d3976;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h295a2e6b6d730a3f88e2324a4b5e20d439575dd16456813d5efda4b7bc686a61a6e696a45c46fb17d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5bb68f19ab70c4aa98af16ac742518687975face3f2538d7111b704b1d03c6d9d06a8d58e6312fd9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48157da606b94ef3d4d6d6a1db52111f9fca571326d7c192cea5b844409e0ad19b3c2e2842a092a1a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcba1097f8c71572f181e2e1b1dec9a29922e4ac385231cd641843d78ae9731268d06bb369ea5b821;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27ad4090ab06a6606dccf051186e2e078298e561893a473fa336f414994681705c2b7f3ed23e1633b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4b5e36bb25273565d8fe5dedfcefd9a04631aabb91963c65043d7b4193b740b444db29a15906845;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b2549b1c74786da2abfe7f69583e39fd02ed56d96de9279716c2274ba5fe0ac6cd339df608aebdf3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59d0d045bb69d72629ca1d2cc6480a2be396278fc5601ba3a0d3fae8fa506355f99f9f94df649a27f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed78e636cbd622ef50446051bea9643a709baa7ecf8517d75c8eafe47ca8227e80a3c16a95003ecdc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96e1efb301434583d519afcff0f5bb3cf31ced9cac64fa7efe287ef39e2959e8d06f219e90867d6a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dc6a25dea0bdfccb71957e81437ebc36417adee5f9eed416d6404b8dc1e7ae75667a44b15558976;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h779d9f2ffc769cdf9d423da0c1e60950a828782235e42b4fc5e4fe926ee3ae0b3a20252a48f70701b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6a5636da3c79a8b459a76509560bc2a29dc9a361eb7a2efe476641f1c4a97c8452824e2105d25e34;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h270772d7e915dffb6431eca1331761192e91d1126ae2399d5b89fdd9f6f917d8b133aced96b3d9593;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d24f6e38b01334b244a7f73466a3dbd4095e6b1d0db3a482e50f7977b16fa3262243ff908b8f877f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h175ec59fc6af794bc247a36cb77c5276725e6b8cb21fd1429565551b5d3bcc1b03cadaeaafdd34cfb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3586dfdd22d7543faa1a368b828eaddee849aae4651cba1c34b96a3fc4503e53a55df8b40e84c859a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e442cbc7a3894dcffc7373e29ef37cedc3c641843c49ef062eecdfb06f9170b812d92fdb5490fbf0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2457d622cbe256242348ac6fcc01c09e4787e557850e19628f58929a925a12566d08a3a5bb8fb2c95;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h701e8d35b0320eb5e84493734a941b728490f4bb025c0cc382b6c4433b2d20f7a1736f45e4156737f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8027c19f06cac812ae6db10474d79b41a015de39c5438917ee08e6fa7b1ea643b94aceef4dcdb6ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96ee48211d7405e23b66608c62bd85de4d8bfd93c65126ba606d0f2c073b74f7838ccce767af97eaf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1415b0f289a4faea6e67c5f5f1583b8a98f078ab06a7060ae774fdecaec09a537a297bd4efd649dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee46d4b85e96270a2b648d0a8ad2ac882f7e2c42f9a1d1548e9ec16e0449e0ed3e495f81eb32feec1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e355dfbf85a42a1d6e1da2e6b973c5bd7dceeb5341017dc5d723e4bbda140f64622bc630599dd1d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cf6f0b7695b91e618e574fa147686324266fd4f6bfa8c4de4906842aa9521e3027dae3484a2dc33f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e80a30bc3b355507c9bf001f75e684068ed7318350044f76f164ab1c08cb4dbcc95fa2bcbd11f3a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h914cabd3fbc0a1f0e85414c0b2df44152180fc979069efb10a3d0987dcc9ff77dfabcf8596a6a4b60;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34eeda8deae465005cbb749a8f06fab7d4ab527959ca5ca239740fe5ba5d05cbdbf39264694986262;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb226de210ad6daf89a0831cfd94c9cd04ee3a3ca4e5c38528c9de3b13bfc8aa659adbb50e4bc1cfd8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h908cffb8ed6f6ccdf4941001b9a68e6b81763d5b4960d8698bfdb2cea5b4abf1fb964fba5329c6aef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcffa078d4a8e99afacb675f17c05bb2a7e08e88c722f50b9be88a096d8a71621171ecc1212f4d3189;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd32f1a21266626c6b3be1cc3cd7d693a0ceeb92300b248f52983186a1e1b0ffd520bf85e36e5422c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffc405ac9b4456cc14626766132291ba7c501634ebeca397420155fc98a2c2e50ad20d4a80452ee40;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcde4320df67beb4a110911a7a74214454373628ed92e706f45508d8a4e726fd54bb0c075607bc7c87;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf09d474cd4299abab69b28c51b12d5a134cede0ff81203be2540c63a8bc5b36bc73304cb07886cde0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haca537e1b84f31c1719ab7c7cd1eae425b1a8ffab2047d6f3b8a72a2838c66fc4941021e2c5ea6406;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f6ce4b64bcc8dce433b84e401f62a4137ddcbfe7d169a845b5c5dd30c152dd4c815e2d0e6634e962;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93ec3cc28f532fb937acc93885e532d99dc503eda46b1489522190f4eefb91797255d84d4e3c2a41b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef9a704f92431e2785d1a3e35bca72fb721e800fe6ac56bf453a5777f1fb42f344c03cc5a4fe99110;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd936298667dc8a08d89b529469d666173b0d205aecf79d9512ae9b974e24124e30598ebee1451a317;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h459e7e144f38b457754db48e639d2abaa2ad16b27620e43ce16936e5c00330da27f50406bafd51d4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb10b6c7fab9d8cd799a457f975679c04a056bbc04fc3623f1b44c5df41f0dd5d69c73a97c9f681ab1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h646abf2e04387e766ffc7f08ba326dbe373b8459e3d2c9918bc1dc39026f2a737dcddae2278b41557;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e5b972a78d55b8a0f257bcabc90f6ae24d5bf2d33ce0907fa50b7db6f92b0a94ce1122fd985e9ff1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10dbb84269097175158c65cc9ad677f506311ee8bb659f3f2bf8507f8fbcf69daf2b8e311fdf4806c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2255ea681a3851ec40536ad7ed052a17a77ec3f3e91dadae3beaacb72451ef5d31b1935fc379d08f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22a0e165c5c209f0a45ade3549a7c583eb5349ee37037ccb7413a428fb7911f5797bf0c4511a28836;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h511f5abf9b34d5c42ddc50249d318adc501e188457a531cd6cafd48929984b1fa386157b1f3c4d878;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87a699aaf4249fee7ecc61469facace0e0c30cea6c09457f4d9fe7c15ed431e8e2a754e432fb23d46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h841dd571d1eaa04348f7987c691d7d09f5e71e7ec0d4e4819e2d06d8c2653674b5e0f72622312da8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42f0fdb7d02159fca898d8538da96afd4d8978c27f02e953fa116c089cca77e1a02b6a5e4498211e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fe430a786040a2c4c23b63dcb1a157cde0d2ec07742850f062c4131d4de6d8556e1164594e76a40b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b4c0fa704966c745c57f5c115724126ce5e0eeec2861d5de9bf270d541236e69a57ac1dca43300d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e514cedb6b7fa5303c877411577f566ea45a5e0aa50c77156ba67d4fb29747a88adcaf614d671cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f2afdc5aff46b3a750703ed6457a41928e8cfdcef29e8701966e454aa913f85038b2fa75dc6daac2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3a01d7ff209426a1b664266115069cd7df800023195f529f8371ac7e554ffadeb77085a79604e01f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6ad014ff4960fb3caa56405e30a3e9798fb42d3baee18ffbd4e2ea8306f440fce2675c8cbe11b64d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e7345ab34fe9af5f8d3210ed7b22a560f2743c8ae94d61aff5f968d62340c4c255e10db55e09e0ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfca97dc954b4bc3c6bd94b26ce4f51b020caab0d412cc8570bf984a077c2d5e15c9e54dc8e37a8c1c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf43635fe583f7fd4177e80d806c17877b8375480328bc201cc168f501af3409be87240b540204e2f5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3499f4e65cae71488a3a0d1fcc5b50b226a0eda9f041968dc8884fc78d9a69ee0729f43d15c83adb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb7bf5add2ce259555fc876617d733c1ec714529bd10b68cac9c9498fcc8c18f5a325fda1ea6c3fa7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8dd261e74960de7f3c55b97ab3f6f57ab0e2cc2e481da4f9ff59ff244d1452bd1ce4f1d8d20b138a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d2a8a3433488bced0eb3e6d9698e6111d7ee9808992e93bf21c3f7a96d381644d252be9769c28f63;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h587d9ded2b637be5c62be71c4595de726a762776cbb70f2e12df04c6da81399dbae14a8ba8156720;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h442e8cf5c6c2e5a0d929017b9262179c56ef25425dbc095c93ae8622434c55070ac626746ba2da4e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba355e18f31614f0dc4e288d67c8bfcb3cb1c322bc97fabc3079e21d6d4cd055256f99939028dcca0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6af0a958ab54eb634819a76ef6bc1b7108e7ab2b5ba76393778998dbf92e5a2205ff9302bfb961c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3b89b913c1d8cb8d61a4dedb632d49d0a38145c494943fb16dd7a8348984117a7ed0d34b2739c726;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h342c17bed5103bc6020d85c2449c641f4a11247946f5256d264b1118070b5f10a21d60460b720ecd1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44b0dd4380afb9aff8f5b62b39aaf2a8560ead79ca129cac1ecf20e1d9186946a7678c22c940ebaeb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb14e18f21fc62ed531c10b16fd343ae63bf50afc40aa637df15a51e23562cf0b7415ca6624671371e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2dd023f27c143e86bf70c84e2eb38eaacc237b0e76f87acedf907e61946dea65329bc712e017f34e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafddbc42fb1e9e8d396be5b4168ee315254c2a3e9dff4ca5b6b926484df6d744eb4b0bd718da22a1c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77d2b4794ba92bb8d0136b622a1412efd29aec8d8641d6a9f80a6638f9405a33a7b2d3afee5d53707;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce5c1e4d40b49b80cd7aa20d4afabebfadb64bfc08ca82365b7e874c4d0e3dbd14c4a3158e6b1f28b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6aaab3a71f76c1c673f55b07b24cefb23f546bbe5d8fb0da4643fa94693ebe337ef14ce3f6811959;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfe4a0fdfae56d332d0bf058756dc7810b593ffe6aada97fb78c48e4c5f56025b19c255f61d613179;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13807ffa06efaffd8b8ebb9ed9308624b1d149fd346780207f4ce0664f15ddf309f9ae010d2f740b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c88cba842ae417b4cdf09fb200f416d7eeb6ef4c4f540a94290db633efb9b2956967bbbf18a4270d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b312b77b2bfd9cd666623dde0c54c73ea3bce90457f4d92819e919a90eee8377772dd6c48dccffd2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h625775b29b34e33abdb0dd46b0a7d2619da6010aef8c49ec94af4855841177cf80b20739433367ea9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bd1481b6450739bf47910fec1beb6eaefcf529ccf17dff26f0bead4f6b0452c1d2166db834bbd320;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff393c0f0c7bb99857cc4596a74df0855b91c8cf9a1dea9b8def5d098c8eb5898b47f31bd30d261c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68f371aa630b785890ff0069a043c070e109b464080a6fe0f5ebe8a5bd5de070ddf7d11b84c322dd8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9f25496db34d29ebeba1fd0ffcf91e8189d33c1e5e5969e3c000049c0819959596d97d56bbc19d12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21f74f0b9817bb217465ee089ec80f451cca96d3e4486c74c1ef2e10682aaf7e32e830be471a03595;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb751f9b85db86d5ef19741e359741b76a5cffb226aa9445f00b0c65c0a57b49feb3a698ca8b7923f9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha93c7e07384417879d753685171cf147158a724b22f348ea8622126d82d8611c7dcd3cc2e96a40bec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1b9d8422526c130f4a6ed000828c72528a6fb26db587408951153a0540682c9827da8b7da2662815c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a9fc570ce150319ddbdd38aaab0b0f93d1f3986d5e0770082ea16d8529825bf43beb5352046f66dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h117dde544032b6045360b0a8ca34abfb6fce36905b0692f6d46ae09a334449aa3b5c0cd9e0b76f0d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fd8ca85e88548f567f254e1251874418d0f1aabfa356730506a2e9f85bad90e0abffd0f0c15bf23c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5ae2d41e574072cd2f4cb95a5baff4ffe87db41e25e82cdfc4b5ad914a578967466097602e7a2eda;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40a200a48ee3a956da9ea481da01981660fe983bb537185a5609550adb1af8bee21960ed1bc5199f5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1768edcd88a33188bdb5fc101d338f19f62dd63b4aef927df870e1de4153c993bfefc623d4c2b0a7c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfbc4855d39d58ad1058f3994eb81bdab72004774b8e2554fe7a884e900c89b9999b3fa813d4d05c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha69554b28f5e34469ef11ee6b9bd6b808449a50abd04e205c501e154d380495ea504b55a8f3fc0b43;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha138277f0d5857f2277ff05681f0495ffb64867af28e3fed19369ebd8270fd92bc1095b80daf6e46d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h812cbe9b16ece41e6b1758a4d273f77d44a6c5f2d179b7d923be838d6623ff07d8b7d5d8d3a2640c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9067ceb4f597cf30f50efdea8856ec4c83f0c0b6646be6911799f455dbacf15813ba56daa7ff21b57;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68d9e43305611e00bd1aedf5e0f3c672f988a77823e112354335111b7c7236e608900f5900116844b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc5f19e95b921053b119bdb52bceb800663af61b74545864308f6b28d4a5cdaac6be8215e16dc0e45;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d1eb966046bd8ce6f47b3f63347dcf75da8aaeaefa75a627c4f0d580bf32f7971860bbc713f4b5ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b865fad514555f824016bb7dfce8656c828a74d80a478ce23f03d96a4b1966f4556733f99eba93b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h946bca27ff0fbd0f11e35cb4d396cea848104d7219a1f06576eda7642a3a1c32cf597b99175a3a751;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b74604e144d07513917380ef612f7d3b109ef7087503a263ddcf3f3bdf4b14d6598cbf10e404dcc3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1c6ef02884f434fcde839d86737a9f9b2aff584d0e68549e6d39dfee0a3ee9666547687443062b85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h201da4f7d715d21b1fc8f12eee14b0b51a1555cd0581ae7d9c72b7c618f210c6c16fa4eb3248e04d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90dcb26bb420cc27f702653e6e938c8795063b40d3b8b416c632196ce8fa7b50ceeab36d243a3e3bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7e5a61aff4729f90354af7b05a69362222e27c4a35a86c411587faaf240043b716df55b093109a330;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59e021d880cb9cc1cbb198d50e53ec52bbc99db50f7577c8c7ae37c5c372c8d34dc823f9e7b5ac965;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb73bd6cd4b17b8b8a0d7bc6df1fd2d10a514294983d8849bb5140629257c67df12e6dc4e91bb3cd78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6fc2b6b1237f60a6aef40ebc3a03f2536dbaf0166529afa5e7788cb42c3120d42f15ad9dae6ca582;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d48004dfbd8d951d8d1487796e107395484a4977cac687cd0ce226ccdcab4278a006c06736b21b46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf765f78da05412b47188f9b715ad45c2a2f0baff2309abfceb7d4858573f67f9760bfaa02674035;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4a75e4ff89a9248c628a49f83f828b60e56531dd9e00bfd420dfe8ea0beeb38cc0e9539d80b18b44;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34ee00b77d10fa514e17a19c6402f1516de4cb4f69efb41b611fc7a209ce16e8b7c062b8bfe807104;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20d883f155b464fa317dfabc80509c57918759f7cb0522ca1ec3b4d061c9d4f07421d97f468cc3483;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab5f26fa7f8d02e07ef16bd003ce9601952a850812dfe1ed469703edab20ad3a54ed89b95de629077;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4ddb901f665bcbc94463e8e0403145b4c7aee07051ce31b5cb338cdebf8e497b3834ea33ad253ea7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18d1586a2b5f9e52ae0ef030aa9715e0985c029516698b7bb7c4fef530da2c1db036852151ad8ba8e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23488f972f9c5605732cba3ebc23503df958d333a94c34ade7bd35e5d56eb79a3b3b6cef1fc8a06b1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc104ae5bdf1ebaf8651ad783bd306bfbf31a05d1c712431b9bcb34748f97829efbea5c46194d32a8f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fe84eae6eac5266a1f9a3a655ee1e7986f1a84f494caa1b0d4f6574d398a875dc51dffe261a232fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28b78a1972d0697f0e449377dc47d07e5b1c592c00d0c536b47bbccf98be85270f9f604f01a42101f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2424c2be08d238c84bc520402f2c8f9fa805eba9a4b9551be60126b7ead2b043f755bf2f208b2a48;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7d4f3c18e708753121f3570cd2d1f4ae5a69d3764e12c504d5f1a843f52667a03e7cb46341652204;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5879f7b62edf7df35101d707675a074bcda7fd90239bd89f1c498b3a6cce8a13d6dea6c6bac4bc0c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8516833ed1cfa3344800b21f5132e4d57be8f34c28c099314452f717549ee3a039e91b72031103890;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefaa79de7232d8e9fe54ad19f5cc662ca0816bad91d817066f87f122bb98a1dbbabc12262732805b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16451bff0e7f5119e7cee7c0b9592993ac29310408bf887affd09021bcf14e05899bd5b422729fa39;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb163faab8ea969f850a5fbf8971720b79542fdf2201c851f6f053b4cf746f118f07c3a03273b4514b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a7314d66488a0c49e498cce1bd277f5a831b8fea2faa3f1d56660bef12092db26b61bcee7ebcdcd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heecc859cd13ea5e9a173ded16588b0b3ed505d3aef28639d6ddee0e0b2528e6d2ec0ead300255dafb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2917145bc89574aa5a34f55a008a65eadf8e61b09d2ebedc40f827e06971ffefa18ae64d0adebb85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3583504f0c303fe87f94e6acace9c1a4dd1d13b57d9cfa4664b3aeaf3a1ce2ec85f7a2bddcfdfab9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a8bc0d9505043c451778eecbfab0226befadbd9bdfba50351586145a60f1e757b8c23a294e7d39c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha624f7b9b478115c0103da173454d230f61d4fbc1665ffd70138b4adc414f4c214f6d5f16464982;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h28561ae64bded85f8495ee715dbc8cc4fe1a5438183a85bfca759f1d97209989e447f8c1eab200bc1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf340b87eda8a47b744d41672bd3705d241a9c32b5f0c5ff2b3bc6585b15d5f58d16fa55ab17a06ca3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82d9eefa6a83fea53658b64187adea36c2112e40e3cad4be130602c578c800a448cc99de1546c8506;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3e86f53297fa520c103ba65c05a6cdd4ca0ec88678989e87eaf3910d4495a2833b22b31782dfa24a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha758f520fdcc5226f225ca514a0f6dc906575adfeb4b12a4f883561be4ea8e7c33a9a433066afa8ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5729d0da50cccb2f9a34044cbeb23a66b97e0221ef8ec273531fd0491273871d3d8ed6c831ba033a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b0fbdf125c002cbcd00532669ad1eb6b6bb599d6ef4be90c9cabf470173cb8b2062185c7ad3d50e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0651da0cd146195bac0b71a616e8da248567e35e2f3dcc790107ca1f0569c220e6084ccbf3d56356;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4ecc5f4d507e97ac44f5f64d92754b2fb85afd7f503f26f196764077c32040d0e013e714a5baa60;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h231764bfb0a284ca009a742be0b6fc2b4c2f9153af09344ceeb85f92b829e9a1e9a904b500165fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39f14f91e923c87843518fb335f7902e53d9d0e66e469e45aa7c20ca7f26fd83a976b319e37651af6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha26b11e405473c0f3347f0db35e643391bef34064d7d1bbae635cbfb7d661c53d2326acbd4d20ff02;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h538213cf512952b2fc7dc7e82dc62bc6a809177acc9a56b10c76e56a6354e3a04450b061012795a0c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd1804a3eb3d456de192f0dcea1478278dc60e22c7149dcb9a852871f24902c6d79ddc60ae3e255d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he79b50862952eaac15ad7152df3fec0bde65116fe542d8d3a63cd2b4ec97f7bb3c4d866f23f86ea1c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0b1d4472ced38a5d5003080f54640ac472d4dca0569d2da2a2b73cfad267f701d531a86245835c1c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c1dcef43558c6e5aa563726cf0b763881a4c0d1a70b90258853e7a989a0a31fbd2801c0ffae94d81;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a8d7cb497323d7fcb2dd2cee277c3df513f67c6095717a71cdbc9c1f552a34a50fec81ece102ae6a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h953e2a7f394ebcf47d35500a355c2752dae473faba2548b7b9a20df665cc50e0d207fbc72bf7077e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd62346c8ada2c54d1a0aef5b8ac153a20a8363b906946335dd41e1b21479424343318c06dbe5873e3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5046a8d78cb12794810dfb3b2060c7fe0ce4ea431396ff725df664b21aa805b2464f756ee61ee1b8a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h332d1176d72d6dc31e1b9c3c56dc5cde4ff03a80b8cc020f550497198bc64b865ab672c6fa3485c8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72880920e810f4512ec55bc3c9928f1b20c10db8b0daa5558a8a0cd8ca8d33fa089f609ceb86d518a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h729adab78a79596611b16078b30dce681bab6276353ec77c3fa981113228c7083cf02fb19197a1183;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16aee3ca73ce943a539c6207b43a0aeac5fce3305a5829e3d9f17f3014a354bdb2191f97a92ba41ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8daaee66acd78d75819c112a281c494d9569507ac79ac0147d6f81eca81bbf4962becc1efe9846fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbf1da7064f4db70bd6707436e67bddeb1acc33d3f1c36bbf7c84222bba1b2a1afc4f006ff9ebb2ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf39f273c57de2eb5bd341e03944f1bc5519cd022d4237a10cc9709c662d3254655aac9dba2c9b6a64;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d22f375f4c9faaf4f1bfeb48448145819bc377cf4a9a884da113bb1b63be7f11d48e8e497c38f2c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55024adaea8e41c002c026bc7cc6b471fb603e4a4e94b2fdf2416c72ec153fc503426a54fbe28567a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf6668861a90768d89a746109ea786711788b3e2fa15476980f9f3366b00e4f52545c719400ead061;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha08520e67e5d50ebe1a7fd7af62a13fa9545caa2b3e3f467857322dd0d273dd99181312783441deda;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac3c29ba915821c19dbc1733b22c2052a541f9c83d5e615b1f6e216e84e50de5da28e123a300abff6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6728f1ce297cd600e4b381b3eca16ec80672759bcb8abd0e4165f42415c7cb5c19b9afcaf3988ea2f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ab2b6fa603be01bdfb860f19cb4f9019f4866d0ea73164f8092c42e687ece5dba9918898c4972a10;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h403dcb7c2f26dedf64f55ef336e59d7b2bfc8f4bf46dcc4f8f30fb074d6798179c56023d3cdfb6be7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9962177ad90258f3df22b59b47319c11c464eabd9b88a7728a7eab7ab51b061821e2795d7b116504;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31810b1871292cf4e572864582474c5eb235f724e6d8001fa6c68b142040460431c9ce312efc6d7be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb09ca1ae27109aa4c2e6df2a20059ceeaee99c250a1b3da87aa876881a0199c6f58e1a2e64e4db570;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b2ec48da3818c803a3974862eb5dc0f31f48ab9ffd9080af49acd06e71a5e4c62448c1e7dbb7dc43;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h898100ac01dccaac7c70124c6e615d9ff070daa94645fda3d1e580aa05bb1ea9a8cd4ff2ad2e0badb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6e28b37adedd484f6aa6a4c7ce4a49e8f0e54637dc5c1547dc6d66a9fa4607e9ee28a38e471b9732;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2e68278fe239b219da60c5d929478cf115e4f6a5858f23d85486ae22ee5bb435ead7dd25a3354eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h119740b671c1dbcada427a7d2648498da00da9e2ec19b60217684d43005c6b239a543f6d198c5e011;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc961ae30bbaf5b93ae39969623383e4f0c9a9a10ed71d3a49ed413827ca3078ccb34cd402ad2d1770;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8b81ffb4313514e6e27527e262e9823b1e2b8accc340c14def79cccd9e2bdfc78cb351d2e339f2cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb57ee1699a3722039c4ff60958c962d3a133fa3583a9f90471976b1b97194d172d77838ef996c59b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91277c3faf530a968a3fb8e1f161246d645def65863d564e7079844eb4b1594170e80c2b9f3ad8843;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8dce1258750c5d96a9325c22ede38a6a2b37302f7ef339abf459e922324ac0f9f1e4a363cd199e2a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ef15b22eac5692eeeb29945719779896856f3874f18e69baa18f7b4229449cdb818fbe642589616f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d2f64f50b1300476477ae9e1ad70e1d9dbb34d6ceca0cddee0c594a254eb7552a6094b85004d263;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd93287c588bb65b33fc848eef9d954d8c383508747b0da31ab1f6792b33825ee3eddcf4f719ffd13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9f3ca134be58eb62e330f26debc354d60e22ba5b0c501efd12b29418057f766dd28015eeaceee5ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcecc80203e6c61232bc9e109c2de28ea2fb0e45f7bf62fd102ed3348ceaf22058ff49511017bf4ede;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbde47476c84590e20f3243a5b903080052b5372b0b9a8e2bdb6d5e3fd82542e2dda8e944b7f002c43;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h670b51b7d66f319bfec4a7b45fa425502c7c743849ceece499c787dd3b359cb5d83f2a8fa591f7452;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2071b2881f62fbf2d94553a915d9aa2530685d7966c027b9d2e6c3f08b908b8e54c0edec595d281de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb6797ed07896c5f545d542689ccd753c996d4f38a877a465d8a62368de2b62e6dd335bdc9a6f130b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcd739820c96955c31c88729b255d75a0e83aee98b4f7d7d50436ef8ab9ec94c3849b241bd14de1ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5bc576fb36a9da2499a5ad488cc43f89a621b17f7903c830ed966f0c644a5fea3c929cfc88e4201d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd14669ba0a85a576031f7383e0d166018471380a6ec1d4cf6011454bd85fb0284dd8f3659d1e97256;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2622dc8a3deabcf92d90eb84ccb13a6abf244b3d1321bfb85a6cbc120b022dd24d0ab403d3f301198;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdce0f1af0c40b744fcd58bc578e3bc3d27de8486f64f29797a3715a1748964afc7800581775cf388;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2f9c6f9b53023b25d7b4a53294e41d61ce8f780e90d75d6776b905684737efaa55322c9ea1f96236;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8da0d802a0c357217800e4a0b6078c18207e057f9126e8ea1493352145177df53a61035eff639cf7f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec305e6ed8b8a781af4b200e3862b6c427ce276fdb6b84d777556a9cf3a268ff6d6d8354437e7edde;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h768d8983dd89ad43460ea9ff9b08988305bb1b10798c98d1eafd25f8591cdc17881f1ecdd423cbe93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ac583fd1b0a2c2fd09185a92755167790e1f5820091ea7dca535525338a14b10280abc7ff282b26c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd842ce3a25529df3bb7d817225eb6807b6da278d09dbf809e75786c88edaa57005510055d3d149901;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ce3b76869ccaea3e787bac3a2a8f01097a5bc4ce6a1975b5413c2fc3b48e4d5ed544083e000e2d6c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5152e24342c8782c36d4667087e7ddf023a47a999c90867625e1c85b050b764870fc3694e248eac9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab63b9730dc2cf70ce5ce997d8a541739581bb938a3caccd146dbbad44cb2000e928a23ef3456fc67;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc7423a240aa330c9f88751e491630f3bf96227877b818e9e54396fcf2b70a2a6a6722318f32b991a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h974d28ca8c007c663aa47b3383aabda1d6cb4cf29a013d87147db787c8594387160ff9409afd75ba4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb61f346a6eea7aeb6858ba84cc7b18ac1cb9986cc8b26277b1fc026b47ac37639f617c4f22e458d0f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e5e8a9101d8c1b6b1938a82df1cc1c6b87792cf5da22c7817c92fc316640e2a53e1a8b1b3a187a8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f8564098e22d77a675525361b026f4d7f490d4b43fef9b6732aef22cf442ee7b6e13bc5ab356128e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd21bb21aec65c99b5722227349b4324381f47b1325ddef64ffe27bee4bae3b1d88d6ad23f2a463c14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ebabcf599072e879366e3665c4b996ee7295a34d1732a65383f35713cb9c3e4e2f0aec6158b16c44;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea865e171678482e94df0dd310d131262533dcee2f0c110cfb7bea4fc00a6de61243d360d2ae748af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h864a20dcf83a47b59d63b8cac389260f4463a40d1ba0a29758d5bdf0ee61113476e3a26448d49ed78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f231d1bb51caaf02f5b6951eef08d2c5fb3046225a29e74e13a77d709c153ebf3d0ad596687f05ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86e49030177b7b79139d737cd36d42dbbad179345b2cbf63d0fdaeddf50023dffec060365ba06004c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6ee3a6b97bb0a84df170cfdb036a66b07de640e7a0ede2058670e8ee07a1926562467faad41370c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc07b813e7ec6da764a9ba8b0674a975a97cd9a7358b7e5ba6f23d5147b7d9f5731d8f21cfa2af48fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7b525afae3cd016ca1e73746b7caf65631e6e7c3de5444733a69ec9f980ef7c9be2335b7b92fb3cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5fb90e683686d729215628fb44125b89148c02dfc23719cba6e139d4f12a6064d6a598cf01c261ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19b438826c56d8abc4646e877b461fdca640b2501303ac3482dbe52e336d07dbd1fd356f7aeabc1b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he497086057ff006ae4e81ad45c5ce0b8222e4000bd40c1ae8d7504f543531a62bfb418c95c26b747f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe99be6418ac3e7fba12617cda8ef32e03cf496ced5ab1a80a27bc9f730abebfe26de30cdb6c2a953;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5327768afe82f192d7ba159fc9dc4ae10ea77852bbc7bc14b2cde94ffb8628bf6f4433dc44840c201;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h45eb24e1e5ac5ad27e0942bde1097956ac6db8fc12a4896da386a3bc5d6877e9678ec7d2925cbb716;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda2441cf0755b12c22921e0f47e262c004b7256d7a817f05b0e6218f61931ef03664d848a8bc44c04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h825409428ac8567ef2387dbe74aa2fda5e5c651155db6acb270161e05e04cb94e9b0ebc8125f83b8d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbcdff25a7d6e8666047af0dfc14a7fb69cc6784578aced734ecb402ade4efc3fe2f249f1c07e0fd8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb0e39192553fa35d85a828a609836a741c3f0cdb33a42d664dec35d4d24d950971e66f6aea066dd34;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb751e7b094524b016438c14909436b21c856bea61750c0e1d7f5f141204b635cfc4a862a59de1ad51;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h421ea46246e5631b4ee805ba6ab0d715583c4d08e07a1cba931a4b5a226fc982a3bb9af74d4c4c866;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60d9b54b4d00f8cf937e3cc4e6a255b798d0ceed65dc2c2349cec688c2c2855094b0037088835cce4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he313debbd49cc52603466b5a4aea34e17658727274abf1f966546df2a21d11ce97cad18889d1dbedb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f8263853b94070322324bd25c47860e3b9b3e562aa445058962bf0f6144cc64b3d52df9c08eec4da;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae99c697b11a2f97d3aaec201a71f9723939b4310df64790bcf0145cfa55eafdd5d8f0fa231e2602e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd2a7b0df61c958b5d373729b38f1a894434bada244e7a0df632272ec3ca3bd4c4a958d508840e41b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8785ada5b9b9617a96908e0170cb0ef891043885ff8738f602fa09bebef34887ef4dc4fd172571ca5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb55e195176e1432583b49956a314ee4aaa45aaf1f281ae88c489f8fd121e7c1b9226c9be2236ace3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96bafab64996c202c58d7d17a09917712fe060476e3da289518ffc53828dd3eb2ad584cb02bf7e9fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30bf92dc8ea5e512d8e4c8264b9cd1c1bddc096a0551ada3ee5fcab2432bff42371e3edf28308a549;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63f89d653e56b9e2631593a890138e28fe1aaef47bf6e9a68021335eedbc481ed6a49e0c69b1285b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9a36dc5069af90c40ca3cc31bd85145f1da255a13459dcd69dd95dcbc529b307e2dedd910fc4975;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5881cb7e0f8a7978a9aecaec597a37c353522e030fa1253a5c1fa689e315df56210a0cb07f7765c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4009531a34efc990d8d6545fe562b1788902262ec0889dfd919c35ef6220bfdbe8ed581d557da05ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d9b009ffeddb70a0d569caaaad72f62836ebfc19ba875a572d0ce11fc71e5ba332cc0e557e2568a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8887c97f68bf19d9fab30c584c83b049314102874d71c90fb327ad34f0156bf89f808a464fa97ea0b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61838e91a485ac94ed5910faabae73ddf1622aa15c640d8cfa6cd356c86ff24a3f530d611dd7e9100;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7552bb6aafd88d1fe0ca305731c8c76d3ccee88711aed3435b84ac61f1e98516379fd601c8d1bc47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h735074360717cc4a7bc7f7adf68ab1954580dea7924621373068e1a9a1340a6d003d7268b28aa5d23;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h221137b47dd815a75ec303f8f2c83dfe5ce46c04090ad6648706e2c9ef0f17e6000ad413fdec2f45e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf154c228e13ab7db294789551a61041d81f211f06911e21912a1a4121ec1383ce1a0d5e04a9fe2a4f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e3f82368169ec9e8af7147afe321171b872982f9864db003fae551f5106367a8ca7e245a0259cd93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e325123d8577c41279a1f5ae96cd20714a49e1baad477d91340004c36990184b1bd6cbbd1e03c819;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9037348846c74a810b0d443a3638282122c6cac29c801ac330df176f487d852d11d2c313b65635b26;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8faf145955668d889cae14a06c06e2a0dfcb2c7d9cf6efff06d6c7431bb680c5778b4bc1287339d12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67242541f6773797089180acc62bbc8c4710e63461bed55966d34eddf03a857d4b9f31b6e38a26fc0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76f0a23bf96bbbb3a7faaaef8b79d4f1a3df123d621cd6212cab89cbd12234468ee878c61d063d3ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f5743236f0e3d01bb1f59db2fe7f39f82e48c49389b1a46e90f13fdccf4d0cae27295be27db94ed4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h741e1a3d864db3c17d45d471efdd6b7e781ecd7b0f6238d889d05b600f4f1fe2706c06d094bb67972;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd41698c4a9f8bbad1135693988dcedabed70afcd78fe50cf8bdb1b10062902de7b41bc9b8b5c209f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe22fc61be39260c7d70a7f5b35ad2c1ee3b17ced88ad1a2e1743dd4b0e0a094dc00b3abb1ea5f329;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefd4d15ae6446dbc1f30b86a0e36d0be160e67de8d86d4fb2fbf397991196a0e35504d83b46fffe84;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4ebd8932ae497c6f3d880689cc1f77fc3c0e35cd97da7e6d6b0ece2bbac3736dcae4e39dbe109814;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c2c268d8d0e03261e39a5eb1aa1d20aeb20eea85fd640e9d0da2d13db612dc3da5c896afc83c5db2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb63e5da91fd9dc53c60430ab7de3cd882c783d1464cd9a62cf62bcaff49c8d6ebb0191cd3a5a0baf4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfd84895337e0eda9f213a89d226953268d39338adfa8648e5472210453039c8ac99331d14004bf13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c76b3791560da4cc9fdea75a7dd432deb99c6264143632499f3d2afeed1b5f3425a2fe33147a9659;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85919db4040bd6cab1a7e884c5e2882710d620f1b481a591b85dd9a1eb7580a9d8d26fa8442e04307;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8130ea4909549d9d29eab0fb8c566db3e0bb4bd91f7c870660d3146617392b0b496bda821cdd9cb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h735d08aaeee10b5a7a397912d2786bf5ff613c52c3e6b8b83bcc9ed04292518bd0602ce0850c530a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9c6159f477ee041e290a288e3b3f95d2227a41697649ae7859699fc8dc71c40ae8060f539c584f1e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h265706a5b9ac40a1d9dd998a6218f156f041fd176cdef341fc2b8de08be63b3933339eeab3044560f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0826e18b58fcd8d129e8d70b9de5ee22249e6f0e2227e43871f5cbab3e14274fbac11765e54c5fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1e887693998c1d2587477cd444f9ca1a4393de91cba903a0b54e1a9b025c74372748f49a131f3e76;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6616e4eb50ab9001c781a0f7d262b86e4db8598816320ab411c6d3d8af197d32257f5602a09231f42;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4af61916c70eb412f3362acee377c2ffed30433126b0deff1c366ebe10292deea2c10436abfd6e0dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30d518767e2d5429046ef2443b2753ba4c950e02c73002e2654f051571b96bfe3340604ab3be7cd1d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79d01ece56cce91592f60b7e0abcd36c86bcd9efda84a53f16e11d3a3a3ae75f15514d4060980d646;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9cad338d32129eccc95c3536d4e8c910cd056da0c169713b813bc77ae5a058f45c89a68643fff9c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d9b0f940d40b35e14c5d6505c28df751698fa813e265441f2e6fd561a752c6e5eb6f00de1343269f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c6b8bf23243e041295b6b25132c4733ac50e1ce9a292235dcf660f1b70d4406aef9c2e810ea4bf03;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h142c99a6d44a2d4f71467ec58e8596f17f4c5ceef27f099a1b373cd7bea539efde09080a2b83c8365;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3142ebb38a76c5e03dd933d308fa2a8229d3580bcaf77ea6d3213ca1be9bf6d930076e3563d5fa721;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba66fc0940b1d5909b6e89ea25b443b91e86002505d0b2a439b2cf6d0fd698b81ee17fe83f5483cef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf66b06ed5f43e15a2d415d9505a5c48b113c6b5c0237a11eeac8869fc0a71cbd5bc4f43a8941866e3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55b73a579c12fff41f9b328b56305d85024d1b38568a75394fa35619a86d2ade8e678c709667de002;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9355abffed3306dc931a0e7e8c0e9061b0c410300b6f077709898fa0005b9f7f5e57d727383a3a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13087618d98dece781ade013e5c6ab0b8da967506717524b9e7c305aefdf1367a294d4934f5620f17;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec4d7adc119289b5cb745f6fe59e7f3f2e9476d8b66f2aaf984fd2a347d83dfde817b6967eb46c606;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3857c205402752f21646461229890e28e229018494ccd9d88becc67cee8911eacb482fe272407cda0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc284243e15bbcbb08ec8eb7c38398185612c84d3dfbdf0cf4dac04f2a38dd49d3455e015d66d806e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7acd28aed8b970f61cb63e0eea2b5ad4ea4b14f9b68eaaffd25719536010319018415170ecb5e4a23;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdccc2c59641fdd2f180e73589da29df916ee7fbd1c938ebf6c59f58aa179ab48e9e3ff1c82364c6f1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3b2f0224ec37bdb342511fd7692db90d1dfc30f33c58d3ce12da50246ae6b976a5376a1ddc2b4b54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfadb27ba583ffe022883d1f654dc914044a67024c301bd51e01aa39ebe84cc768b1deb906f96987d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h443b822368a7f63014f6d2afeb9b3044eb11cb8ba1804bf65e04c7490355879a94080319a259fa71b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha085786b70308ff89e252ecd0eb046ce1398891cffafe4aa80daa6943c2933dd33ed405bacb4880e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58c64fd668fb03b91c1d178eabd42addb75aa09bf7ea690e2281f11e6b4a486c0f9ad2ce7fa8fd288;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h195460e8f6134d910679c88c737ea3d5f3f9cd8660200b63bd613413903033460a22639bff6a47786;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca42e9ba4f6d1e341370f5aa36d73ff30218bdea452a13a8dbd147d01ec77b3da326116a1fe5f9537;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40e2d7aa973cea6e18116769fa3472fb14aea9670eef208bbb4a077cc601ba4b5b25f1d0920100bda;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h822c9e9699fbfd44451f64afdb5bacbe368b589c73c2bd318fe56245ff15b08f654c4cceb3e6141cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h546db600416b3f558174af66e4ab4545bf4c7e6c0b962d53364f3cfc9d86e4248547cb3fbdbf5ac81;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98d2f035de548d897b1795200e5b0f83a59907b4c72c7802aef82e37399d3a7d36ff89afe96f480d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec52fba4574f8675f2bd0305350ca8c3892fe1eef0c5edf5c681583c780c240362c007eb2c9209806;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa92a245fb118d7aa0e6ce6a0c4392a7701594157afed2589d4b4496b86b03eeb4a8a09e77a3b2b32;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5911e689d3f0dbf51697dd0da4bdbc82650ace686bf35994b5544732afe276721988a54fda624fcbb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he47737c78b6322622c82e46b502ed85f4b2943ab29a2b119e9e7f30b1407960ad0fd7a8809acd123c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h27b08d21f9a1070cd59053c16a184273793bcacfdf17cb0bef5b69e9294d3ba630d4dc6f75eafec9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c08f6b06df381837fc22a267b47e555740962031efba9243e1fa3b41e023b55582632549c6f5c8be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2731d41332f27c966bf659d6b41cb6179b1806371cb5c16bbe4880bc8efe57da14ad13e0e274035bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7796b41506ce1c2f88e26ae7835b2a594b7a6ad7da671da10b233f39e283eabb61259c38403cbab85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he477c7edfa0ef951e1751bc670eeca7f665e77ba66a38a2d9368928b684657ed36c0202b2d21df13d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce654c87e89ed9822b17ab20bfc7d5f2f7bf79861a7d970c9a33af7c05b09b95e3037d8909a345fce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8028f371c4d976f481ac502fcc9612fdc8697c433f9a0fe16d1a408e16e737aade9c875c47bf8e59e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e214816ebd8056d28ee631d544d211508ea4c28e49ab03711d6f749500f13ad1295556facd9077e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha412021099cb5f8dd2762857f4e2a95c0f37d88126f5438ba81d54656c013197373d92dc4684d7249;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb136c5db700839d4b68ccd03f46ba88f89d18f1584f16ea66b65fadeabf62e760f667d4659b85daf3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7c4c8a204a7d6f0e7251d4bca892f54948fe53cba74617c95746ec7a765425758386fe3447b3bc28b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f30184a80c285e58799d5cf99a4bb5c2dcb43bd66eb9bf0ccb7fbebfbbf5ad4691d2c07f441d0834;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heed5f5e0a7c9a3116c20d3341ca2eed0f0bbfce5f34728b7fb06c3ae5690ab0229fcb2d8cdc89b466;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h905485de2ec45501afa9b294916f7ade1405d84bd41c323465462d77cf590e08c09a6475b3c571950;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a0014c460fa541593bedaebc5b4b01da96d3f5bb89e368f7ff6812f7f0bda0156a493c1b792fffe8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h253473a76800bec7f3da7c6152afb2568eecad2ce59ff9df76af1fb600f4d3dc8e837d480abe885b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd19d6fc65ed5ffd0b08ce1340e2bf1118fccea16b28002aee7ec47f52f1c784490e8c27bf25e25bd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h829f0c1db860d9a20873c2c89389459316deea22e96e9c87306324fdcc594e038fe6b11859367db5e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16edcf7fd1b90cbcedd6172d8b24619a463a34126b7f8009262499cee62b11c9a3e82d2dccfe42682;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c4bbcaa5a5528dbb689013a0a2045da566ea0ebc089dc8d2d84d3d3b4251501f0acd532cb6c80447;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7bdb5d957e088e79560cab0843ec1103f2e28e4e01549d250c8fab763a5d5572628f10a0369e44832;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c3c61693826a73c4cb9f59691f0d7dc7e856a2efde32781cf5f5b3d17a707e93661fa5434919762e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc01cd4c9df56723a87893de7e0d796317a82a9b4251e32aac51211c1fbd2256848856340359e57d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaca9cda7bc74e3ae231ae194bf04d6cfcd9a853aa6e1e8044961473ba34bd3a9c22fa51bc052c483;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fba9b223c0c8bf5f07990815c3bce28a449bbafbe68dab1f7179952063bb0d9e82bc4f864cb8ebf5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c252d743e386a89c0c04ef5d84db36c0ecb05a1bc9bcf124c319e9ae0f413fe8a68039704e493e80;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4aa31ab48a7b8d8ea14c2ad9e22e10c493fce904ebdbbdd5ed57c1861d9c92030af734fa55a3189a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2647fc50e83072fd05c798354f9657a7744388dc01a19909574dbe5324252c9fe8485c794c247d25b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha02528279a105411898a91a4353d6c5847c422dd902b235bf93d118894698ee7fbb3abc9a2be354a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h316a806e4a5d41b7541598bddb50f679578e99e32087559b63a372e7724f77d2a92a1a87729378fcc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4544f1d2e60d3eb7390219ba184fd0c1dd7d31036ecd9652e4d09fde865460b37ce51e7fcb00d26f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12b2bf3611958b21fa36268d9ea04f068be9055c083833bee86d08fb428d5746c3c9c8e1770dbaf06;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9ba7cec0636edef57d855ca251bf20a908e16cce21d796bc93f25140913f4ce9591ed2029d397f3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16f810f5451b8e65ee451bee94ab73e97c7f8d19034ed53d68de7e266f085970769745c3b5ad33a89;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b47f8e2572aabcfbde2ca63742792dea2024cc22942bcd0520f069cea971cf757db147ac5b550272;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd8673ab536550727f81063bbe46743204227f82341766cc82bc417298d40fa3d7e926b6f32d22083;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h25ebdda9f4bf6767f53fbf955181f5a0155c2881d7fb725d7af0d4dea12ed095b241cf67c47361713;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc8502dc1e92d26262989b41825a8f1db0234c49e5cc936c7ca7285fec8b51556e76ec0fc820fe712;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h409e2436b55a76b63062273e0258a10ceb47327b597356afd712dc1189c26698b651f6137d1f7eaf0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21308bd87f5e5f84623429f578bbbb236ea744d782d9f71672a1cff32bd2c532891ea77855b600f71;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9be843b2f572cc450b1ebc8f7ad4d3d42d3f0f3f4c240655077b0f19c4529ddddb6b4f821d336395;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81db8d1ce1166f800c9cbb8c5891bb47adeb3944770934b0071e18aac6aa2f1e254b4eebd5052a39c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc23574062abe733493d9c5fd0af425917d52ade9889f3891f99dc117dbd6056a7f30829dde26dbdb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h193bd3d0c2bbdbdaac4b073854891cbf9dd36a7c3c39b2281d70e8742459ddd77c757dd19ad27f967;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he816b21384c28cce5abe052d320489a82ee04aab01ff33136cdcb78797a75bf21c8fe29e066f36a19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd18da7edf91c433ec669e998dbb2910408816bb1cd12a0366e26e24cc82b5e3b7f8fa360748db511e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h391af29245e2a70559f91f4d5542e1cb88a51c0f73c7903d4539c8f030206a1a82b83a874451f3d3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f7f7f2d5ea57abc091b124a8385acfa9aae6391c7a04393a904352a9bada01a0284a18d26c49cb5d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h329b65278bd1df686decdd35b344b3905839ff0b38d316e89ce1544ff5fd9df9fc02aeb8a7137da74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6d04f78bd04a93044feef63cdb36114b09702852937118bdf6eee69a61e82e46535789f98be59459;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ca6bc3d4227f16614488489e0b99e0fb2e2f33e803b130d6b9d05c3e54c918f2788d1d7e1fc26a54;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe79b28a870be70cefddcaefdc442d6b05bb47150a192443ded66789922b1f13feb16e894e1200180;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2c914a8243c280a2ba034a77338ba6b214738e2281abf59c88dc1327ad2142fe63cdb15cc9797a146;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h276bc30649f1c4959a00607ecfc04c355712d8a4739c1c5e8c3abe7094a9f7bbf9de5259219f55ecf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80c62f022d9b6dfd1312f11f5fe87ad2db8ff33c60011a9e440634bb20e7e885a1390a98b14f967d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5be4035bc4ae66c6924eda5f6118c249c97906b70c14cc017ef9147de151ef31b171566ea1687970;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ce1117d059a05d725c62a1d03b981ed2c19b4be2770ce1e164a394727b41a5612443c5ee0ce60502;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57e36c456d28045c3661025c4d34c087eb75d0f142d4b8bd540ed48b851d7ae508b5779acec61abd2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1416b0e3968bbc0f309a198ffe465d8157df5c6d8c439fcea0441f2f045a9f91ae4bed94885762e9b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47df74cde7e6079070a6e08473d817ce106aa4992deed6faafe10212de27a244e6f1afbdef299852f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3ae0b23d2cf36ebd8b00e2c77660a6ab081981d8c14502f6feacd6ca4655af47b6943367e1a5987cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb560d016bd297691a49149c43d8810d9d8050b61ab81ce4875cbe9e3547359348b2adae1e1e47a08c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h642657b685426e1b6eda77386d0edda1cd408750713471d37efab7187f9c4c2e4698b78b6b79a4a60;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha923a45f125437235b34a0253a0b8c22d0fb393feffeb4b6051b14d900b1648a5dee3fea01e242efd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1883e36fbafd4ede7ecb2da1b3d0e3b45fcf15c61445e08ee5c66cd6496488de6c3a6ebaaa4d7f35a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3cee74d4ba96438035d55856566df21b09caf38e3d3580f5af17a2fe358f355c1037b3251d7ec6768;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8597863cd22d50a288846fcb24b22b16f407ac30fc31e30ae66d462f630f9067cf6e2e247cb87006d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f1e62d682262399742a524985ff1ab5f65490f2ea3241a4549f0be8a23cab459a7bc28c739e6e9f1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe2fd33ee23d9a7186a8f713d02aed01dbf2f31e5aae9f62b21f9c7095fdb148ba82e4b9e74e40bf3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h820e1d5562acd401df94a805b9c326627ddc1937a2a9b6904f337be98b1076a26db90f698a3c9eca1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57f30cd88877501a065e5b137560a4c2844cd27bb188c29aee346ae394da72798faae4609aadd7cc6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb201ed83d649c0a21768fccd25d6637fd486c56d257367866679c958401304411911c6e62b6eff8ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h999642fd77c3a220b6d53a11ba5a4acbac51e13ab3ac8d0d132f88533be73242a5ff4229262d603e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa98ec1bfe2d4b5edd3cbf13da14cf1df9bb5c41c3e1a65374a9c1ec54c22a0cb68a4e1dd9cefaf2f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26596ddc4b98e447a576a14ebf3b2924386b4041f91a173227df9c04082dc7aa0fb04b4d0609a5a14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc43716dfd565ccea05c46def2eeb68f11ba66d4e7883d185bba2726672fbfcd2287c2e6634886b8e3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12d56024b55f08d83f7cf1eb8d79e8553345a9978ceb47cb1cc4a4767206874608c5c6553cff4498b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb0f51777dfc88b50a11cf976c8ff2168b25cadce07c0f2290bb1931c8a2a36fb6b0244ebef97897e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he632d55de04811a01dc01625b8c8fdef5f3d87b42f04ded882ced3e98abade829c235599f046e111d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf821fc98bb711be0d321f7e536edceb9d72633f0e98a81ea7f72e2f19e4ffb463407d42e3645e4d5f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b383211c329c896b7b94b001ce9794f46a4063196f4cdf5637c19ec4cf742c523d34797236169a85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ea4e20c8293d4f68d5ed51c9556bbb316de474515f34432d798e63fe5593d1e755eeffb75014391b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf455f3857f223fe19fb482f63b6fbafdad983e7c00a27c761969c89b1ca2bd0af32eb0a7d51fd4e07;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd80f488d1d74d7005e070a851ca6d5966310555b35f958620ce14ff76ac635c8038b52ae64cd77f1e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3638dbdbbbf1090eb03b77a8c99902e940db68d5c4332b553ec69da04062cf4769bb59ab5c2ac4d66;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf8efa6de7ad1b8aeef49df104c9d76078a256817f7393d98cd8c62a18efbc872c77198a2f9e210001;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6aad5ace0d37069c36385f9edcc964a4f881656c80fd6d17bc8d9196dfbcf8341da58104d444581b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e223d192b5a01bd3b9900369e667478df2ebc97a91aa9d403715de88352945494c9fe5b1744fad0e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9205aa9334d46327c439c27dc8892063e141a336831df03e6942aa9b7d6af7d7321e9ac023fa0d0cb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8232105dcedc52326e36322e5b19d812348c2c4a0b866d5ee80dc991b05705f44953337939a0e4b58;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbf5c4bca455e03414997df65e5099759da07dc7ddffbe550a0f87b461bd9ca5796a89609a1283ecf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7eea721536951e649dc59061135465091d2a6459531c70a200bc3492a4b0333379a23f08d3c74299;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7597b2045ebb910f7b5bb385f7445a393ede0e4ea857bce6c69bc74bcbe7ae4c1ef17df5e5ed5c0b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h883dcb04cf023c579e97c5f870c865b1808dbbd5221644ff8dee32631d425b17997309b3f01a02cc7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbea34ffe012645db38060bb31292ce08c8c587ca1832924627f27f16d58b00b08bdf6689211d27ae3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9059ecede1e7bbf7ee5807182a3320b2006ae525bd9d1a3dbeaf464b59d054b737db27287893ed909;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11c70dad42a6431ba72597ff3d06351cce48f4051c8f3fcc5a929ddd43c914affadc21108bc4fe716;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h940f0e85cf3550d5a6e5e54447e466862950a49a974a96198d35dfa0f4c3ed8f23c55c969fc8d2c31;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h914f4cf4a6d78663bfd03186f78eaf5cbc48082257805684af3ac75670e4f83d4e909724ff322769b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c67549636587d4769fc4bee7ee49d74a6aa42efedeb24a446a51a0336e6272187c1e2107b44ef3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1b1406f6fbf765bb98c8173077ec5b190816f7b41176dd72843aee779d59528f24024434af68b14;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58799c07d33d1e01a176b7e745326f9d695f80663c13396b61412d33f23ea11aadb4e1ab745fc43e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd89c07640b491a597f940b33036da50fac05d395f51e1ca535146e6e5ed2053e7d259187dddf7b639;
        #1
        $finish();
    end
endmodule
