module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [36:0] srcsum;
    wire [36:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0878c06758339c81bc26d5b3594332814b33016a2f53703a6423e82411b9b2d0522d0f86a79a7145cf0ca8dd41cb435e4b635fe28798b77ef027b36990e1a98b42971e5db22be508906dab42ba03831e9b4109df914ef73aa9765f508b2a9ef2c24ae4e01170281cca136c05b0c161ec23e39f1a53fb1ac4f259e76a3006ae7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd0d8e91a5517e05875714a6a825144de4ecb8e666156d7a59b94c7a4f0e078f169f8c77b19d40b068afa0c22fddfa2eed586983267d6d28a6ba1c52d439bc0c680adef562573deaa0074310af93ad287f45f12be00ed18bebdb96b6f1df8b287c05480366bb5ee95f79e2ebb03c7b1ed47e4b2e9caa490d935df72080046a1d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23c7205d8cb9d33b4c0c6d33393a97b1b6380ea614dd5612269c4bfb700099cf5810a6c0f5446b8915f0631c0f736e579fa2d4c43e9c902e601014929ca7da180e250655e3b81f753a36823581c746eadadd759795a103555b2e2945a99165a7d105e9a5c44bfa292a41d469256be1fa750641b5639eb3b201249c2c132595f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h765738f444ab739b55c0ded16df1e3209529600577c415048206972288165db4e02b265e0d232cafad5831006d31de28febc9842ad608eb98043b818aa587324d003299bc5d39d391e78eae8484b1202c0178f0660948edbf024e9e65a61cfbe3a2385e0be93e668dce4cac24b18366634404e45f56ba83aefa9bac51d897084;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h934202948a4e1a166ff8612f18ad9ed82f8b83fbff1ab3341b984422d557954ed7e6979ae8dc5e492d350950678651c4a98b620a79d052ffb2529e40f40d7ffd8ae4be0763c4e8a0973713d708eaad3706482e4a8b6915e510f9a8fad77bfb4a7ebf9cf4818d8bd35abbfaf87fa3ac329cf7ebb6680f678e11a28163cf5e372;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha32681e1df258896251a8d0d41389a49b75d124152ff2f616615c9ab3727a6e3b382e72b7314dc9c67d64cc22057d0c6164b682c83f6f1b61f154f3b75facd9f91b9747477bf2f29c1b6ca4bee0f4e5ee4d93dc34e8f5c70ffcaf033b70f059b08daf4e4a4ea1e58032e08a10710014626a2bcf27fb85f3893c762ea98f6750b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ec16dcac5290bd9d4d153d6a0d1bb59cd17102f5b300ea492df9814dccb0446809d2ff64064f78604812dfa83a5f37cde30544f00a3213b31186a309178e0360dd1d19aeace33c1e35bffa95b378f52d4372cf2dc3279cc433086d7cf787409e1d26ab3a04b9b4a163d8f23723dcf2ce4c9733c729e0ad81de1b2114531dd22;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff13c62013e0f43f5a3506a69d18309b03b4f65b88c80fb41a4bab6a158815fbe90b4283d369048d57cd57e85dfff882986761b14f637558fb106ed65d47cda0eb0df3a8e95d626aadd1ea01df842c91f7fbf30376e04aeac6fd7afd9c7f3514f87af11b36335a17f9093b4dc58228044d65e8bd83cebfbb418331c1852b6b92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7f01ac8fd5c52564a08e26807641acddce47a4904cce3379e205cc3cc6bf718b9ce78b7d52dbd0bd3851f39b832ef1817e78412196ef3de976cf783918c464cbb169a74a0670e2780a91338142f07a4727b961ba48808185a488d7608e532fc14e4e47e7f8d1eebe5356d44fa01fb8a46aae2024184e4bb81ada7b80e9e215b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88c01735bbb49065cf2637980b4bba72c97d8b7761ffb87f8e3a69f846a5d5b2119a95a4af095aa46cfcc4e13ace7231ebc0370a9ea26a1bf9468b9ea0ff3a4ccf3f14bd7772f1a7fe386c7c75883645d11b2b0ae4729bfea68578c14b50be1ccd6f203103c57227ddc13a0d53cd4f105c215a1b4c09d40914719ba18d6a5235;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4985782ea9ea88d1b809b700ad8945efc4b58b6377c28b68cb0b230473510ef016c9841e5d5f78eacce2bf92321ef5b037f3f676e05339fc4df59e8bab087913cfc4a39f8a762d37803eab8a1a542224418c31ca3d4466dcab8cab7617ed5bd7c518499b4c48bc3b9ca7658b51165323bed14688a4ad7aaf49ca1683f403a7f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88871059e935418064a2f65c4fdecf5454019ccbfd2e6a9d96b5b48639510f9f46a4caaf4cd66eea83e40a1dce88040f5ae250e1969fedc57360fbbaa23a8e9a6000be7ff37177ced7dd857f55d8e6eac2a209753456f5e9a2793cdbae0de635eb0780046d7c851169d1749cccbe8c7dbc3333b0c6fae98ff104ba78dfd9b2e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80ba46765189768c45e01364a0d0fdb5171e4624b755d80a14663a6691cfa10370aebc8483b26e5127010d1a8666e33621d15db81c8b15e8afa5a8fd60886f42bff40060eedf0a2d9011fac1c5faec6ba911d5869044253fb626dba7e7cd901003f6cf443b4273843a69a2da8e350eba60df1d60f34e35247662b8faf7f06d51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15872015c0b0fcd59fd3d75360262c45a4a941cd77ea44a934712fa61b9a41672b55a558560f0de19ed88f89c193a9d07dd1f6a253089ea23b6701e14639b05f2b4d9f65830d702f8810c157a3fc1e8103f2c71b128a1140cb9c174aa3f610cb3a18571d6a99de9586a6c597ccf7fb5e891eba734e9b6f34a7e006743bd664eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3acbc8413c3bcfe53034a0f80beb571c793ff76a52a8d0f6a9f4b7356e5ccb62a3cabdfcadb56f3fe2975ea396aa8f9e68155fe78d552c85a9792d8e37d02052d3df7d8e44f3519b61f34f9310ccb58adf0b68e8d71418281c33e0758364352a286b43a4e13928831e90b595dbab7d12da4a04e0ee6e73bbc270fbe83b5a5830;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2b749d0c8ecbf4b5a385cb3fc6511b165e500e6605ac983bc3d564b16929362ace8440f2d6d9c4dd740e5e68ada5bd80f10439708f01856b19ad12033ac7c7079e2d462f3a6c9aef8bd43520101cdd725cf4cff4c7d9f2802b3e72db57c0b54b1ff1a4b6b859d18b7cf5a72445c6db74493f464a0603fe5fa361c4d22664654;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h116cc2b93b68e991f25b4ccedd3c267a90e9175fd79975671fba46be705dbd6e854959dd39f8a4c1c2f072194142a21f04ebe68cbc607faaa847ee7ed8b903f6e0b24ed9c60d8844512da9a8a03828cb4f46b85258ce6086ebac655d8e5bd4ce7e06298ad5fdd68cafd51a86ebbaadd042acdb39b15dc2d78624cbb43064c5d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f976ae176fba65e33ec1a42ef620ff29fe1b9aaad000353859044a74348c44feb69ac35339a90342440ef3cabbecb5c914308cb456460cc3ecd5c6ba59515b149ae560c450fd3e88bd25ee31e91e27cc7b2736f73f2a67fe3429c0ce5312809207c03c70530258092a5af1080d7dc8e02973cfeb92c7aa1ffa976c594502b8d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf12e285a44372fe5c7e86d9900a8ee4c6144d9823326cba068a4e876ea2c09558a13e5046b397f9fea73e80e625e7a3283a4b7fe9a854885d6a80579819e97b22f46269d8f8a2c4460f665a8b2d197d13942acabfbdcde97d861ed5dc851e87c795b6bf981c2167467928d8a1766e0ebf267ce957a7567a8c6bdf237fe3413a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd5b01b2ab3ead2375aea829cb08769dec9560ccb9a6b0b9e14e679737084272bf81ad8d0c94667d1770da40032f96f032124349a8a93b0543df5e727690abc3ba1d2448feea1587907f303daef6ca88d3454b1cebe2c071f157f7ff3718a6dc71bbc1dc913c9742e32be30e844956c38256ea16f6cd896e1e3b39bdba51ec5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38b8f02cef9e28c6ed66b3892de5383e04f5ffea1cc83f5b2b3f89ca9cd75b95198de289dac8bbea7cc23796991ac5132e2f8706a9b1b7d7bab4296dc512f57d4ae7735e4edd8ce945d0eac98b85d3ab8ba93095376684a4e5c2986e40677d56790498c04af2f4221fe2429f98f56b138f6f29609cfec37788a0f69ccca76d97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h965b0e8bd11dc1cb5dc33dfa21530eb644b34cd246ba17d61025da63d3f3c89bb3b55ae3a0e51f7b16ca6570b70713c6fb317b3c1c7f85efcea2f0cbd5ce6188250c4a464de3544ee621b8fc4fe33aae3f6bb4f48ee09722532e6230b98660430cf85627d2486ca1d4705bb226266ad379f5d41111de3f0861c5b64781807906;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f50102946540c7d83011b3f68a34697681e36327abe33062cca7bd053b257e306008249f71d19e3ce312edf519e20e6610ed7d29730396a1221826d7cd8933e0a5cfe725ee489f6170bb78e2296b6a6150770ad36e2cad3f027635108e4420efc0f9ec22e5aee22c76852fe5674fa53c010ab2cc86d75d9b0a8d3ae957cc24e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb53f28c80a7cc27cfeb7fb73d76db3f487b12ea50ea6549d692e6d00eff927b521151f57ec49d897453337975347c176cd4006679b59772bbc7199f70a3a009d99201583be21e675caa522a9ef69ffcfe404f9b6b159c6b74511b1ef63c2beb9ae230ed8a4c19bbeff05d4fe01248d6dccb7d72d663e2ffca160ca2ed9b24ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64917f7f17a87e29b18f155ce383598ffefaca73816e2688571e02da058ff535bec25fb4ce6921ae73506d57ecd21ae1a43d4cb51be0f642829903884a4a1cf018def63ab27db789ee858958e64971c9aae4d398accee58902d90d2fb01bf759e53b85fd9c9971cf3d4ce156124e0e426ae80e59ff70d24a581c2cb110847e40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha40ca97dfb3f0c1c597af243ecbbb6110638caef2e6adb6f548890f7bdbc1ab796411bc48ebe89e1f23b2182d5941c398aeb644f1efa9e73d54ea479ae2abe2f92164e3765d5e72d5ccfa1c1afbb18897984bb497037cbb17f160e57fbd1897ef40bcc313eb5d8f5a16400aec8b177a6c26060cc5d45563e2770ce4f701c7a58;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25290baa16386bbf50d2f3c2eb2b7e26d09f0111e02c555a244ce0b9384595723e88f83e676004b88e7a315d5b9cefaf066a85ad7506438c69b7a8616f95137d234155ccf22888eff76366d17a2539eb49d5202ab8b359f6a1b254a2b44dc0b5722648e400d99adcc21b08b06af276203f980a828764324285ab1e9b0dc91e21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe8e341fe18f9903ec1f51a9cf1e9db6b75c25334360a3ef6938d29e1aabe8d3a5f854fda95e4e89ab1e70dfa17627dc65a5eee4ab013668daea5ed86602c15fb9b548371d5239e103eff17a2704328ee395cce01f61eb0c299cd293c86fc5f5e4654121d2bcccfefe3a2426d680b7a6549302b92fb3855b694101c67b58ed2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7534b9bb3d61a2baac7db493763334e3947ec60f334a05cb363aae8d6440b497bd15ef68945cb66ea80cdf4719e8864ff07491e325165eb8ec1742bc8b0cd9a2046333e2d95f8f203a9a7dc2e97ba9cf2dffde65cbd329a45366c1beb3eccc9ca5d2cc42a326b57d2c8aed62465533b2652dd2faa50c85a03603bce23072c79c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h519822a37a54ef720cde29989ba6f07803d53148185b2fd1248d76c06669b5aedb96e69544d49399c61cb153d4a140cf6e3ba179a31e2b500d618f1cc58d9d2c3371a270654e0732e7e4ecce2a3f6e110cec57bb4c1444fbc0c2f1e903fe3a62278660488282c7ac6762458903fb325647f46888045f6f0139f85c2c290079bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48ffd88f835eeca92f5323ff05af50770a2b56505e5698b93b94d346dfe7b96ebef671d7bbfb639ee7ceae4acaae26ce568ede3fc5853a4dfe21b1f3512ef05340df11e9feb3c91e7baa702dbaef238ac72755adfbdc5f46225719714e2539319d9feab8d69f11690291830f03fbf2abb036f7515d02df60fd9133f40827f98e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8181f5e3622059be22a60812a7463a72879027315fc1cf0d89cc0f3b574a8044ab08015a07cd9ed8e269ac959752a10868d7156a6bd650fa2e081133abfc082c91a9f8187f2f51bf64f7527f804fbe7ba396674ea4a3ecf54a6476287f6e9387f99d28e154c92bbac865a72fb0dd6bb6d5afde5388f8d0121a078f1c7edabae1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5530592e9a3930952f2769687f23e255c479d28dcf36edd5488eb9ee8e5762e5cd4a6da62b7be18f95d8b4e1c87c3f199895b6f25050a8c0bd41f0b6ae571f78936d5bb741a1c23df651091f1db324f6952dc2eb539c7397b1f2bca8e8b54c937983c90ef8410aee32d48e5dea99270c6958158a54a75aa1459107e66e2c0ba6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had43f34648869f60c69986fec041e1f760826339092e65356b29d95caac3b81279be337b4b52e04658e0fdeedf4a0d8b988ff3f22bae6f146c6b7c9e88199b9a4b8de67a2ee65645c1151ac08b7178cb666c19f31b989d0e535635d198eff44c958b2c00e6d633c572d5801ccfa201314fa5d6bc85a87895cabfe0640123b895;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h512e646f7a25488fe1765802ddaa62d6ffc0134c0b5e9c7c50cbea449a1ab0636d7310f490fbce7d3514f6e051a49e6566cc3946af39c7706d567687f865749f84560b4415ea1ffa95eed62ceb16a2ce5debcfbb84afe16430a95568296245a5c551d8ff75bc6c3c6d33dae23e43fb5940a7775b03317c5a7b7bf9e2c5b06c45;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1edbcab0dd58903ee5a35116abc153e6370dc8be8599fadc7cf11abb848fc2b63192eccce1c9050ab2a87bdeea1e7e00ef95030d297ee0521a659a285c5ea743903e3997d8c3e9fcd8fc29795c9848fa1f4239026bb051187dd9fed73061daa59b98883d01d27fe6fd296291b1a00f52a264fcdfa2dfb716682f01c0d887660d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2487b9487d0b87f89a745d74489c5561eadd6166f4ef6a7cf60aa132ec54fcc4b12c930bd2823bec17ef2900b6fb5de57da74286b558dd6a843afcd338c918882f3f1dc361e153b637100301ca7dc4f53b715646bcc1b951ab5a881b3731197c2fc6607bd9df0cb6f7514425c2af48306f988c44cc9a8fb4cf3db388f583286;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7a9570257380ae0994064d7214992d15a65d797f306e1d2cb2098db97efe8ba4b6df5330c824ed6600bdac33acfd948b0ff437aaadfc98e1ea4f06fc3b11df429dbce252e51247277edb3e48702bc9dd754f6566d6b2d62db9537175443b2d89c905af9c0938300f7e13bc6b4db57a8af9056c7787420e76ab5d60b8f4a3e2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10ef4ba884107488428cf8573a1ffc7576ac43d3cb5b4efc1ac2b830dcac4a95931a4df4b16c59853aac0aaaefa67512255dd3e650109cd7ebb2965b01cb9406d242e8448feb7ef6d31ea5cd1ebf9704a6998c9e5a395bec91291ef6b906eb01ad9f8bf353ce517ca01eda7be7be90520ca322823b816a0c7427768ddde79b0f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1730ea481d999f50cd03a525d67695a94edbb1e6fdf172063a4eed4b730edc3b3893116bcf7a5b88949c281c3cd96cce3e4470e7e88d11453e0230df9fdf4081ae8ecd58e4994834bc2135a664199960846f9e6615eb6e3bf2cc4fde572fafaa3a7a89cff3dd1cd39a78238c9ce2b00cd1e5278e2cbaf38634b537d4d5f628d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h791b00d048e88ef980c816092506c94116bdd4b89708f915564f1471db83a27843639e01dd11e268bff6d922adb30a72a733fed111a6c7a19f54a2747e4fbd2f255531735228e7586d0b7c0e287dcc47dcacdfdcd7c1e8ac5c4dfbbf09ee62366f408e3053fdf6da854b31018e454c70861fe93a86f328804f29c70476f8f2ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1daf3d59eb34f09ee6ac9d79e73a87c4273ffab4d7898716f9428c9609cfa28d78a03e356fab2e3154e71ba2a2c7f737591864737ec0ea5d879b7be776e1b33e1e07eb0d32f620c6e90a6938c40311799e6d96caaf6a04f29dde4d88baec5a9513604a6718667705184ed76614bbf62df04f0553bb6024ee5d290e0259b0e64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bcbfbba425782a0368f80c1b347fd51757a5fa799547e734280e6e99aebab58d8bcbb22fe2ba3b6d5e75a07875ea6e6cc64aeb7edcc057dd23bbe52341f75f9317032e46ad6610777e97088183039adcff626a6a8c170e18a0e8cccf2cc46b7633d917517ab699aed9ceb359eaeb66eab885b4f109cf5855072755e8df251b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1b60ed71a1e123cb3ae9773694b7925a2e630a395e2f3afb96f72a105de66c331b1e614063ddb6c067a5a3c8e30fcef3276fa25bce97dac588149d86772e66cdec3181b8b991ab48fa4537190020bba9a5a654e5b0d760ad198343786a1ff41914a9a44a65891826f8430f91f0a43580ae4c086fa222f9c9cc8f50ae5cd5703;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1603d8fef3a9fa6a76ae0fdc968f63237240fbf6810ee4eb7c47cda0cd7eef9b40f650bfaf22c6c7d21123a856e114a4178c70a4f5c94313b2e7bc8e58e2f532c681546155f7e1b4c464619e11222d8b89904ff6d0ee7951b0df2de9d975f77094d670c64c5eb4e0994ccc18fe6bbf0f76f76dd847442ea4dd9b6aad26a2388;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5bcb6eacab816c14bb154c24692106a7075f1e10eff1233e4eabb4f6c71e1b7981782ce70df8698235e32f699e48784e98f7b3723dc49745d2c1d06e011af17817b34ce400901d5ada7d0a3f14845f7092bbabef7a9fdd0d2c02477a7e939f3b86715f41e5f45ac93654ddf06b8d9074681a30dfde59089e044bb78a7164a8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c44c034e6437bd2bbccb52ec6171a4b8a5f282bb83d6eaee67bd8e19197fb7c0f27eb8e9dc903496ef4efc43443daf402544c3b83bf173fc115f8958703c9deeef13131c9b0487eb7ff480f969e5ef9153c8d5cccfade19f02228b2b639450ae81fc6d63974bff1ef5bf4b3e5d38a62e711401f72bfe9992c9e491b252e650b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha51bded6a3b58d0ac7dfd137f94af49d850ceca6269abb1ae4763f9e7566b7d90752e01c8ba530a44d7b2c594e5332ecef19021fc9ab293cea154ada2dd3a9ed1c10a433e52ce05bb213ef2720a308dce4452a24b2deed3890af9edee970f865547a26cb1769495a2cd0a556e827db34cb6a53aa763bf8dd94bcd75c4ecfb672;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc3e764b135d486d369bc8588513730b1e3ad2a8f531f5c4602097f63e122b3b572386cfaf7904e9ebfed2062eb33c284eef024e4307c647129e8079c1ebd8a66853f798cafb46394a5349d3ce505a9a626939fe2253c999446937aa6fc0137ffa9476ccbc4a54d5970b60aa6ca25db38b8ddf34644f1d1da2fa38e95a8d7b69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h458c0b5a74bd240d4826bfb750b1e94769dfdfcfbdf8984f6dffa89b137cc89087a9b858c79a2a234e0ce03f37bbb4eccda11c579f71e60899cbed73c6c0f239e9e46886581fca584ba8c78d155095829d72e5254ac5385cb1b9f0229e7665d6694e56ef260f8becbce916cde85889fb2c8f8e2912bfd606c3470201bca5ba06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heeedeeda5d96560eb966e5c134ba4dca19a25cbf384d4cb7cb6a16fdfd6b2b19b3771f9fe2ef2ccc27094ea7888e1813782b02c82eba91c235d71c55cf432cb20c9afefb49c101841b08075b83168f4fee095fdc87c34e2263857828272b8b23e5c2ab26625fecde467a30336d70718b92ab3c7389e72844e7b5ef8d7b04c580;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f263478b139abf6d7735c9e85de8f0739017a152d282fab8007ad999b2f1e3de873a028d96907cc7febc0926aa2bb994ee16eb6b1b125b509761dd9a5168d745155a0f19a2b716a1eba2ba036ecde13c58bcf8aee95f58192644c851a21474578a2f0cfc1615de50ddcdb50d9ef1dd50ae75a65380f2c0c07a65dcadc3c3b45;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he68dd6b070322d744859df7df19b9060fa57b8d57c895afc9045efe5a15ae7e4c0738f8c5c1c1c4ec6e8e7a60f335be8e72f461e7ddf31b4339089e5323a4e66661aabd1fdbf3944a78274717c390babd59e0a95c5157144556865de1557aefdac712a0343c4d3fb77a07bb75bce7caf2311f69281aa43d81b46745ecc97caa3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bc526de29e4b23419642c0af9cf7be1f2e64dc0599a9faa0290c2497cbf514701e92abaf54c3e6d8468b103ba28b64c957ab25611e71e49e185859cd4e2b81cd6a7e665bbf613085f48628665d1e7a389a25d996a78553d02417949b0496efd734f9fd8a0cc7c9138e91fcb8a87c1d26d26c8fe2fa13ffc65fdb62f511e93e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cad9a3f037470e022a6f78a8ecacc0245ab17771b890c88d809325e10571ad1b181c283f671816ffe69f307a8c18aa9110f891c16c1d29869eb17bc39f23e99ab919188217e0b96f2395e404548becade53ef0b60c0a3f6731e6e237fe8d73c9328e91b0f4ce1d6b8f6b60e8303720d196ad7f6197778ab43a2d2ea332c34b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35bda35134fed8d124f6f49b32bb0c76222507ea345fee47a59a588a172e4fdc01060903740691f010df04d0e64a8aa87b0341170cd98c7d4ebd8abbc80a01c1663fbe1ffd450c2923fac71286f7a14a620628235d32ac6cf2e9de4c34e363f68f63bdf99f9c23d9071e9a4f0a16d60af4acecad71c2401ba945b9cd297468b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cd80695c38e1b2fe9994c0567e31cd4be9e8ffca7ee0c177b15fe9029201d275b4c9bfcb26450f6cc580318362cd82904682c338455de98c4f937fde17e86ddb7f98e6fb7322d3c1ef8469ba052be8b6cb52f1e0ae3202a1390969a2b53209100ca5002b8248208b145067c6b694589b05209e3e192f8a87647e88b59222096;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71d07eaeae55b92e5f3256073453066306e0dffea3f5a461bc062d7b95e02e6a7bfac4ba8ad8449f29ead4a09a69042a67daf46e0ebb3857a697ff99af3fadb37417cff39e6f27984424fd1b0653564514fd97c384f64bf85fb3be7fc99bde374912546c0bdc542cba58e79955dd56c0d43990122e2eebadf8b2fbc394d2f34b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h16b89a4c63bd7785f798738550630086f7d6b931cdb3d4b5977345b95e101fb88f0271aa2708444a0ed7fb273a535f63761e4a4da33804e2a201d0a56d57ac18e13fafb4893a27f44a800dfb1a0f9f80e09aa96538e55d066f3567b36aa2917876007e8a9ef8e9dbee49fd13c3c27798d50faa3c8f121b45cefcd8fabf22eb36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2405431c3ed435ee447da52cdee536b85f75a395adff5a1aff62fba412f86d7b47c09931f94903e08d6787f72815966f07034f7a968010b84ffd1ef56461f0c95f8860e227744b1f7c3342435515d16dbb897478d29eec81971b8132c7b5e39e194683b206813650896e7ad03813d727cab7216b6a25d53203ed59f3eab9bd9c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h763e44ed28c18f0488b7afcf5f0d75e56db831e62ad4c0437a45488af9ee2e99fde0d05cfe6423ded97140e451781935ed6ee8a9679595bdaffc18b9345b7cec1cd9e5aabc1bc6e4c0d5a8eb60ee1820a58a7d180fc440d9fc0cd4257bd4ba82568b6734fcb03876a27e5a97392f80b803ba62b997bf9b6cddae094b61bf41ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f10ff68e1d0102accba489d9cb6bcfdb82cc445ada1624db02443db027b65cf77b7ad09665346ac1f97d19e51d9687dd6eaceb7904160db6884f59e1fb0a39925c2339deb8f8662906f12f78cb244eec432064d31b3464b39664b2842cf38024d858069732d3504b18df0985c2e394b16b00683cfb8c0a6fe256d2494a26b20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0b744997e0264ee620dfb563b75023aa68ff1d972a20957bdfb853c002a5fac05ccdf940f0fee2aa4e6eb90c7789819e894a855e1c188b39b9869c0d9218e2eff3d97023b59271fbe966c0bccf72f618084448894182605f589e0f7f779a50980dd7600270b61a66d1856364a8b68d43715d535c27705669053720f38516062;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7110757b463fef62d3fcf893e94a6733c4304e01b2dfe3fbd5da63e89e6629c0b7ff07deccf2da360364bdb86453a41dac379d76d06126bb7521a9759caa463114608d14729c69bc690a5e6867a62ebdd9613fc0fe78f1b66d775c481dcd8e47b23a6a71d5b429726ce32219c965d91a64f777afbc591a33b8a83fcbf187981;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8735ea53d0974600d25cc8023a8c295e7d16d56ef754fc5dfe6ef94556b4754177a431088362e80870f707952012c6f60ed88213bb78477d83afed147de5624942d1fca55f981c1f6c9bdfe99a799b5913be5fd17883895e883d051008d3813dffb308ef86d137954e91e1c0247ac5f4b7eeba22c7bdc2f9f07c9db195578b88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17e188e6ccf6f9c8f90a37992e06f64d9ec654aa135687a853b6308e454553deabc19fe0f0feab614e0a907a33d12a2a83ec2db22adb70ad08b5a15fef68339436b29cfae2b267e071016501cc4f24cf7f63657acc3b0d1c3a2939416d91cc9f2919492a0f426bfd80c2714619f1042f602a2a1287c3470d62fcfcb0becc74b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ccbe57524e4f3ecbeca49b292bc7c625a28c40f1252fc5e4d580315b0021827a32776368bdbe29285a665608aadf24bc25d1903dc4a6ba42c382bc946dff066fd99d879505715b714005adf8802710b18b3f9e1e59f883a951470caf5dc060be9aefaf009ae5174339b5f0610e358e9ab8094210222cc0a5ab6e1cbd8c29f43;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49250d27f57ce2673b40032549f7a4e4fdf716cc00c0a555068451ee22e167fe9bbf2e008c18bfea3181cccde362f65b0a50f091db19f941542f62448a9e3e074b62932612cfcfefa1fa39fc7765043042e1ef648f3e37fab1efade33d26daf62181ee7e66a130ce2ce0142854e91102cb965317e5fbc6095b3dc542baac90bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a3e29d576cce93162ee998d31cc11114314edd1152244378bb1fac1aef03710f5db2f15f063851f54f7b2df43a3260815fe8889000aedc86a883aa52738a9dd452c24a04717477f67773560d3d3c73adc633d107a3280ee47c01a1de1dc3728e9630f6550cd7c2bdc1b526ad35611374dbe24575e6994dd0e9247d8887a7051;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d259c6af416e1939a5293c68ff87f8d9a56cd2b9d1bfae3b35e94cf35910abc1cf63a3baccada31b5ef5ace57b0e728897f2f39d3c82e61eac870b46db6c5cd9135c60e3ff03b17eaf3b73ab67443d60babdd1309c27b4724c2c30eb7d32d77b1ae97e29fd3d7928f43a342670f78b68436807d83dc47bcd1deb6365cbc9dc8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h600b30feedefff0fb6962a026894cc33f8e6cc83e63f0b15846b0e8a0d6aca3480ce7a8b1ddec07cdc83ce44a90b7e34c7522ded56f783cd62aa2bbc9fc65ad5f1f83d9b8b405cf8e0b5ec921b0ba896f3bc6daf1d294fd111acb808ea4927119e22ad1bad3b10b5dda0e8e16e08da143e7b9c696a363ce3f595fed9f7111652;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ae91af497b22bdf6c237bd503fa8e9a74d3987418128b87adbdee4b744dfa60009abf145d9cbe7914907e0b74eb6f90badabc24239493a6d75f5096ed0b481966fbacd9829e5d40c36e0841348626616b0955dae759206175baec8d3c2e7c1a00a2c7085d750dbf6bcff91143043892d93eaa51e94ba0b577f93ad90b35bece;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he75f70d135369a698ab237953d6c683d76ba5f8123e5ef8dbd2bacbb3e2449d7674a8a7e83d303186d012176685ffaec48376801712823a78e56d279f3fb335a9ac1219f00c28c938b80d64aa0f6014b9ea97e01b3c5fe0d31f4d6f3df7da9df80cdc7831b2904f67fad37cbc71870fc6c3da4849d718d4a4790a4ac57a4e40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8372f7b92738a92bd1fe5027b1e75a9624ef4f47661c68789cee3165acf4169554dbfe8923133b0d72626686acad63c11700561e870636049afb70c99e45b2b16564b84f6f16a020936b01c10150ae2c2001ce0fc7cb04fe116b8485c70138c79df0bb0d679f3194b537d31e94c01912b03eeb605d8c1164b177dc5c14f27ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5621d20ed12e2a659010e8e52a84bef893456aab84ef1809a0b063992428d9eae821079af50fb4a2eb24096a9a557cc17b20410ef1a05b1b223f7de700365c3ea160158d872317e0f4c02c45314aa766cbe47189dc277d759629d1a57864ac4a26a54d3407a82d8bd9f7ff0dea2b67e85e9f2383f4a346b9390ac287f40cdd74;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdebb8b8f5aa95c70eb419b3c5371e95fb9718da88cd1bc3e6c84372c42b77018aaf7ce766cc97dd6c230852f3eb6399cf5b427e7c121d9441201dd847ea5e0a92cae4ad535e793277a019279d2dd32748c30ad974db1d846c840450bc6f01832e2b2940e05ea2d22adff222fd7d4b6b4cdcc28d1bc5722a8d39ffab610b059f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1048084d3ba5291fd084c4527795015a5aaf9881b59c7995502eac84a156f00057f97e7dd5d930c3fc463f635d99020ae0af36e8a4c9e8265d3bc7103b1d0a54a06554b9415b8d7056d5947ec87ce0c4f60dcad19966092abd7a8cdaeea6988e95baef72ed3da0007c71b2498f08f7f58b8e121d3805a4eff45335408d576177;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68176469ed61be2a25f4e4eb70a82f53140be74ea0f65f0b1b6e5c66bf384c3b2b982dbe7afbd7c20158ba838ada69f5f9f7c15e5a3af460f6e76117a87e0fa3bff797c5dcd2fd652767685bbfee751eaf112ede15bb358c1706387173969a69f45041112b941139edef57fff92a12ef822761e9f0c2ad3f0b3cb9d3f3b13259;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1ada3d4403407a37d4c493052035440ecae0387f5974bb26a14ed7fa80107c094a7fe691421fdb64c908fb49750a4189cd45ee6369af24a49326c28d3646b4d5d1b934e71b8592710840f8152aa54a301965e7d19178046e722a544961e8f3622f306ddb543ce2be1548ea0e51639b131ee23c76528c837c281281a92fa6fce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b0b532eaf0f2df8a12b82ed8193d153e2e6272a5207cff6066729450aea20431df04dce3d4ca10fde9c816f860565c237ea92589620b7b8876cee98672b4046d1dc855dab3391eb06e4afd155820868b10e3dac5a76e9c4d270853853a672693d17906e4529017372c4b2e1a61f44c73941d1705be5e53ba37937cf4c73cc75;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafa67552c4f70ce5f8ebe7aead63ce77df9b7a11ec43c687e3524d970a8ae3902b6427ad64477f3dad9d620bc8ecc7c06f6603cd19efa313590f0e8b86e4a7fb26a26ee2ba593a4c67824ec2feb8438ef71c6c3f6f59b1336798436339cd3bb84d22a05423cacba6e50f711bf16d041af60eab56ec60beb23bf428805ec732c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8a2f644a21a27c6c559a06452f238df9ee7f27d9bef086c37e53377d69cdadc9cb8e1fe561919b5623b94193f7164e3507c06b910cd39ba4fa3f00a5233ac12d68885208d5fc6f072a5c1e6f944bcad837754682251f2766e7edbfdd79019a3352b6e614f93680c5059efc437dce2c549d5cebe39892ab81aaaec1e42b792ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e646a554576f5c8d6bfe3046e8f8639f9bc8b3458014e948d8c5963bdcaf1fe76d2b6f94d17605bed30a45be2169323c62c8d13beb75977cfeb6369336d6379b4ea28c9ae1039b82d8dadcbc2cb87ed712555fb6d5418a8659f44a5ac88504fe65a2ae8c926cad98ba235057370c182b14ac6ce94c61ce1e85f6f75d75edcfa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7219111b8a8c05d010dfd907e33896964e3f6932d4ad19a32bf3d3c7ec5e10e62c40ffedf4837309c5408b830ddfbd0a89dcc3af32d2077efde25648e20e1902ecd7377a06a6078f40830a55a967dc9ca0560a4dc490682ae3c4860c31790030475ba118019e7d08cb887790ea96afcd4bd1d153b73e684567dcd7d7cba7f29e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h756c3e51417b0b8eb17d391d385d70c1a3ad93f8925160a4577342ecb525b19fc75b0434dadebb72afe53569ef3db80eec70ba60c5d384f9a198ecdbaf49c0c5befa7f004286b0969bac9797ecb9fc6ed2d5542b9607440758fe1b313800b8ceb7bb9f5604eb8e60db43846a005d9b5fbe978685236e0bdd469aa87f2c7d2e76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d78bdb2f207b7c2ede680d8dd14accb073b7ce82d5ddd9281f78f2403d93d1bee8060b61795fb0951e377c9c11137479213ac9dfbfe70d6d55c78f1b11ae3f1f9f45914754bd874a51746675d9a21f0bd4b9987fe951c773f6b6616f732b6eef3fe7772dbc90cd4185085506ea5d794f29e71b6890b709ce06b4d05b696faa5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1de42e7e4183a41dbd5af58b5d657084fc327b6e314ae623e35d2c0ec2ffc7c3680a3de602bcebe7517f72b41ec0afbf801733b6c23730e2b04ba3f5e0b76b9897837648396602882d07cda6da0f653acd5e99a295c0ab7e5d83da4d092fba3af6d9b020bd71222ef0e21b15ba010040172baf5f2bec8af7bedb451456f77cae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h427d246b1aea018d4bb77ef0f9f0890ed2d83a3d730edbd6012ba5b351234d40e1bee06e4a9d907b50d12b31f619bf9718b0e8b2a0f51532b91d75af06205cb312a271775c5c2d740eb1aaab266a0345a360b1730e146c4ca0b6e559a231b4298913f36af65519af5c387eb1413d42a50a1706d130c6af4911f0742b7ff55e57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab824d2efe85e8a56d7a8adb589ce25c67c241c84b5da631188be100644c19cabd9e7c33a6ab44645296f19d3c680eee4f3d036315b894dd00a14b66efaccf9c75279c5a3d361e992461f8da559f5c385b7d1293671b620d620614b28743f41fd476027dc83addeef70bad45f52ba904fcc268339c0efcc649def456fc968a31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82d6b4cf527de28e9cd7874b7e25da6541ad269eeb61fafc8b7ac050ee4934a378a216abfa00e6464b902001dacdd2859265aac6fda06200fbef3b04f8e05dac89e1df7a7170e1b58cd36dea3e45a10d88307d37d8187d55e1946cde73db1c3e0f9c6ab48ab1c4fb605d99fe7214fcd1dda3021d689699e12d6cc1f854964e19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55099bf5020679f605df44bff1ce1df38191a11c459b27f255059ecc19599a3388c0fdb0745265eecd434c07dedfcbb654cdb0f62ee64a28cb3a42e793a081f16b5029b42773d7374bcdc12c5171be269a08d8a2388f6ca8ef36624d2eb0246b69c7d2d7eb3da479d9db56a3a7b4b67fef13ba4efe12f70255176e488f91363d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78d420508c0cced82c0598a22d9aca72fc75a8556959b9c53898a7ebc61da242315657110018ccddd35b3037b5183afb0b6257ac9d7860e9c58d2bd5712e1a864780724a927579bacee7b9c4788dcb7d16fee29004bd8365e4e0baf46e1bdc50130b3165dda096d8c0bde45f7a6cf2bac9e50417fd62b515d533df3bf344c92c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6fb6472fa43987869bfe54247e46b346b77ffb2a08ca0ebae1accb5417bb4e7756347ff9010fb9e09e90bd35c5542bf253359aa995e831caad74a9a10aeecc7b7491fc54ee7079a83db1f2afe5e720ae78506f994c8831c89487756c6faf41eaddc98085b214388c028e3608958ee861fa47567650024ea422e3effcf49cd97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30a1614a03996ba02c196e9c04ea6ea8ab602023739249325ab65c0d45106f667a3926bff630704966bfa0f35b9c7169099d3f9677b672b56410185212416931654f74615911191a9ce3380f53fcf4e4e5c00fcf31527a2d2236deecdd1d2e9ded0750ae24f26fbd708a02a59b76b6b49111ccf7d1ae39f0bfaebae39ab0249a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c5f699ae843b39f768797928637b7d20988cc8198e21341ceb97791f08abbf342ae9f5b99338f0efff56227b785ac261365103f8b46d224d339aea8ce320405f12ee18dc21ded54975bfe9ee584031e0645bcfbf0b8a31c8d36c66530ba09bda20b548bef0c09b490acf2bfd6952f44db5ca3b017d37a502407e9dd7189a9d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fec0dabe035a3ca18f1d8476543eeb2c5b57376187b7f1be59b84d75d4b073117e6bc418f2ddb02c572a89bc908fdc787452eb3cf919cb297cea548a7bd981f1bc9638869ee61eef1262536a4d71904e0f9ae2aac676a65bc1219768cd40acb9f54a0a9cd7935f678b605be3e2ccefa35ca5dc8b53f3a062a3a5f60d6c84f78;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87d99c90f23019c2eee2caff1775a8f27890e82cc287ecdee52e0941c5be0c604870f17473caea652c56853792fbeca3e424adc9d9989f1f96eac7dc7b8051f9a0f19c2494b3aa78e6f9062a15a404045157de62be8732fdf778f5fdbc34752030024f6e27aa92aec7df64826d6917049480c4a8bee3c9506f6f854c5fc1566b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c3a6c7946fcfe29182f49f8e54e3e77bcbb336c687e54d76d499b5f53d1e03df0159ddf25eb23c8fe59da55c2f55e52838a4a93ea99f1274c0ffbe666d5f25dd1a3e58e74c8a7eeb4360fc84b07f6322bb71bd719e333aca9e5ea2a58adbd448486c79fc921b87d642cd93cbeb26670232cc2fd3998f933bba1a7cbcea3bb93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he53c64112959269ce54a04a031b347124a09a9063396e71714fbe419e0d5e3b9adb6dfc70331edefd19c2ac88b673833b2b2601c58b05e2a5e9d7b236dee6fd3137c8c0032915835e289cabb53459ba6657f3f7eaf480b59b4941b65a8aaf7be5ec021e037552ee720c676a06d5d3793031d67065bd7ed3af27feb232e74759d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h873f9008e332503cb77a02fb176109849fbde37a799230af3d1815dca6df899f6e1272c36f79218bc70ca0f1adffad188cf1169866000457c9b425c15cbb0071ec431f9190e52c7b2d63ba7eef47ece4c53f99833a60b15a0cb5ecd67e25eacb923a66591822a269f81af44a32bc13d5fb78180c9a377b26a637b6fbcf78f81c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c189e4f0598fd9e31f611f81154e688dd9fc2f64e82075ec243db6fc0c0ec874499470207439bb54600189621fae437af4f4471b29c7300159280673f1caa65cfa6b775ced41ecdd4e5c5a9a99027e9c740c80be5f75831fbc366d61f67767a6a0a40fd5020c70f3be04bcac5b8a01c6caef528c2f58694116f08e80f4b658e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d7f7dc64aa0a42b4a49149a837cd328cde80bb0011ed70f50c8098fb6b679b710ef5437e171dd05daa13d181994386b53b04587887df91c7a8a38435edf448436879ae59a145bf4926d0fd8aa11f0bee448473342f102bd1f74a2bdbe8eaa67e5e151ba98f09614eb0a27f2000bec56d20c61e3e3adccb9bdb697453ade0676;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5b9bcf4d341f4d54933de43efb9f4b72494d683356317b6ff6912438ac70ad6acb24852f03179152f5be9a1ebc87a38bbfde5f3819c4e664e4c88780e6380aae1b3e047d886866561316ae7c8477522f2ff505566b242664da28b9bc3beda43b159b334797f8de393f98658f9f41a1bc2fc5709725cce9ede93e099119c6663;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d91c58b594083a28665e6c08869b3d6507543ec97e8e2446e3eb0ab057266045d5327a778c281a6038d2bd43173dc85c6fc6186ab7fccb1f542ef6b5525cdf656551d9f62ef72d8853fd41c243a30d0568d21b7c032c64c3b44c36f59d5fa8c852c09af06d2aee16abe92243f57d891fc532d3b60d5c1a73fa2404c4a68b97f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfaccc2171af857bd5405afa96b9814fc19eb6f428c2434176d5c63a3d413b9ee20346bb61092a6eaf975375f207fc6fb034da1aa897a75eaeef118d5557ef77f5dad52978fbfe51884b554986684823dd0f3ee56d172f615c9d13f07c8accb1c1125256f50b11462969cb34bf37c9fed1cf2818a4d2d95d2bffd885f7f8a36a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3eb1edaaa24371cd80f746f60a9f5345e499b20e78fb08c75bad7d5a9d0665cee95b487aa4a38f70ab568e57eba873832408a7bcc224f7c2621f6dc12c8b7b3821534b8fbac0788fdf83d41123ef60c759cfe38d6cefd7d327d0f4b01b8f3056e316c25a68b5a9f516f8b119e3c7115fc416b859af31e54e1d30692a751c403;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c4d02b5b56a0e82c36618baec21a98fccadf79b286a8c44393092d8434f7a30f2cd074132d857fbbe7280b1c623769f85fdac25bc8603b1f3c4600ea791ec5fad59ccd8e89824ebf78d0f1796f1efdd1cd1eb8967c39ce7be9d71d2b1e6915ca3e623589bc61d390745528d5ac0b0c4d162d8b654538243f0901b554b8d55b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h716ebd99350f84a449a5824d3ed32a73aa040610a398bcecf212a62c5c7b03a8b2e1ff6860799ec4619dd61befb38f047276b7920a8379f0fecb0470a284abb9044b9ed84bd1f97d36013e573f98953f38881af8e15d2b85d5b4511325f3f6af71f9d4826bc11f87c65a2b1fae630adefd0c9ebcf05f7bc414f87e1853c52ec8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5495fce4ff5c2b6dea4cdadc30a00b5ca76eb522d62738e9ee0354ff84b241b7f0d602cfeca8503728aae861f7d8c492fd93b9738594a6afb48bdde6dd210f8fd036eb6a33c64ff79894e2129c2bcc64210785429f8bfbfba3f0fde34c951014a1525282e814e61b2619c78899dc259c295f85d122ba775a925620d733a8110c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc48d7af34efa2a8f2de2c33fe152b8d4f3edb1d5618359e02844b8dcc9ed03f9cef47df62fdea1f7b014c0dc6f29adf65301b754ecc8e2f28c04ddf9b74cf2cb88c5e0c45a5df5668b18990e08b73c8b1c4fd007815c8860eb2e91b1b9f97ce7c921b425b740612fb7b3f940931c0de396d8226fc2bb4e598d8a962a592db24e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h109159bfb0aaf3206d01dd79977010fccd735cf3cdf768b3fdf3595efb831eef57a9cc21b37ed023e43a6e2f447cfc86bc506d00fca7de9b457cef477b361b27aca8fc4f21dbc26e6dd7517acd72b38b920f295dbdb65a0177efc2e1ec306def7e07280da824576d86da8ce92fe0c0dc33ef0f4b2fcab60561a081a0db1d49;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc14148fce297f69c62d01bfa316bd715682997fff10f6a3904fa11a90e57347ad924a4fe3ed46fd354e029bf25827bed148464a1fda3407c3cb7a49eaf9c1725ad6b27b87b69ad1076cae1f99f36eb3150df1c010494d5234ca0201e1a75cea762a7c231d479c955bb7dfaf3848056adcc1646783ad4f414773d84f73ce79873;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10af1505505df6964010ad3ee5b77deb08c655a6bf3e2073682e9a3762cfb280ef1e2294f6265e640c8f3e8b698bcbe583e9a5d4a0ceb6b511c24a4c15edaaf40f6c740570ca0eca95b23df29bde63e7f3f1b35759f9ad9539a290c23712933773d0f77f5666842eb851c3e94985e3264f023e5fc0586bbf5b24f2a9a7aa04f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a6b87d04fd01ae717b46638fba7185840f2cc5469ff25e57ae1f09dac9389ba9465de6dcc532e45f2b104bc7fb7a6b90c7f928029ecd58580053f8d08d57e4c7d53f37c5cda17037e708b505ed74823b39c2807b9e0b1d084fa8d2e4bd962c0b4d1126652e26975cf78b12f60395e5698bb97cfdbceeb1325b0c058d064d443;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ca6d3564b643d0bc25f13782b7ad79b0077ad0ebc6e0682db5b2a94d3eba18edd3cf7a8f2ea4b7eaacb9037b5701ff88713ccfab5eb133d6ddcbccceb07534f91be2e22414263ad01ad9e97367ca6de5000ba1cda66ea90276994457cc32640763c9becdb05d52eca99136e4f3ef4d91ddc34b2015674a16d546e56e4b35c5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8598f9a79612c8af748cee7c96f5ea8984833d57dac9b9ce99f7f7c6a2cdb3e2a0c605a2a6fd07c6c084d3e9c662de29e1fda81aa313e890a0fd1ab19d560667b442b52b544fbdb5a0c3a84567fefa24a1f4a77810c0eb8388470255ead31a669acb439e5dd42035d9f01aa0d98580e3b84d595b7bd8aff292887e3b702a0786;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0a2257b35582ede010d5a2a520800d25a2e4e463e4c89d0c323f294f07cf13a9d9a6dd2a5ab359569616f9ba49fb9133c580049c7bca664c58e22937d5c5ae72ad38a3a73e35f0d9cbfb4b458f22f72790b788ce69b3fe819af360be46b79832978e9cc1b462fbe762f01023d5a6c453acbd81d5dcc14439cfafe16d9e7559e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75868669d777e34da108a797fad69079a06048df6b87debd775fe10a95ea3f46d6f73016c438354b2fe841b9af62b5666e1cf4607c752c3e31ada56f7154e860c54a87fee0cb4098b5997f711681f2c59b944748366faa2936028f8c5fa72b8787880808c09241838d37b2a8ced395d68809142bc9841d10c7b9efddd79c48dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52baec11e34bba5589462be50097eb922e0fc9539ca5165684482135285a7f94a130c30175dd503b63fb6d49d36b6a20c46a01f7c2cecf176e7549398d3ef98ca8908e4af9b6edb096bef4b085b7fd83c640ff863ba5553fd31ecc84bc31582f5b4d966f8276c6ef156d9e90baac1934df9a252bd6770a1b99deb46d0c259cb4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4633f4c725693ef891005f2972727db9a95485f125cad07de8427027d9d2093237bc9e28a7e47d23774c0d9a798f245d4eac4db709b3cc2d6d1056440253748a38f7c664d70b4ddace03def022267019df6eafb37709264074cfc0f6ed8f69b2806380d2d270b795ce8860b9063da26bc7e3e918ea0ccc166f02c4359aed9a43;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15597b270bac5ae6d6bfec096d95c9e2baac2e0fc57b25a72511a11d10c6a580600290a854784f56215ffa42d96683afeecdf9f2fd9ac4081dee4308a638c0f2ecf278c19f6aeb0809adea661cc3c2d0b04b26a2e93508cf53369369378fe1c96c5cdc517bf3c431d65068578713cbbef996a1cbb76b9291eb21c297dbfd86d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49da009cc755144eb18077f41794f45dc178db180a49ba7108332f098188e578b32742a4d1f6792d69fdc4898243ebcb567e28133336e0a9b492f415d553d5c6bd278acef1c12c2ad1f4c10ce2d39f1909a841a64d8394f4871e3d9dec57f787f7b68f48eef6fe7f06387f6da8eac3114f004ecc494db68be28461e67c696949;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h619618ee63debb1287c25ab475a475ebfeaf45c1b4bbe932cbace940ba84f32948d3bb347c0217ae94d2e164adbf5359469f318c8c6db86d9d8b5e4408bbd76888f1b623429b0d2a2b6578b12b3e559937b022b5bee326c993d0a1a8c65b77f3b414b103007573bca645d2fdfe510ceb30c32d2986b7d57d09aff57fed027a2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b074ec41d509438dcc34d80376633bccf6220818e708f184ca650e55ed1cfe3f15e8457da3b0464bf54e0bbe81aacbbc85e950bf560f20ba175b2ce5eb66d6ba70f275360518b3e01a7e7530aa670099e0097cbec6211cef523ebdadb3b03cff104342bfb127eae2db114354065d275cdb79d874c41a58ec830ab21516ec23e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb296d17462ee144ec092a0b60d38822671c2f4bc32e3169ada4b8d9f7ff2a1023825fb92dd7b29089694d3c43e98404badaf5a568aac1369cf14193876248ca31d5903bdae0f96a56d30d0d30536dc79c9f6aeb6317fcad1a6a96e66204036bb03799b780a04f6197685bf20a0a8be883d6b6adaabcbf6724edbd5f068c9282;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf78178f0a4d7d9625c93a6f1dc71891c899065e2ed7cabc4d9670967b7eb435ae9bba71cefd7ad1244ff37213683e93c1b22c81f74d67fc4673c8a78e7a8ae528c1346cee018135483ab171da8a09d8fc93c69dc8d311e4c61d5966243c8a85db7c981070ffe76f6d8c578633b71a29c18987faab1348629551fe3d505ea5f7d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb59cfb78cde4f818a6b16e78d85ddb616e875f8871e9129748eb27d293aecd74656d323915cb5c112408f4ad2c939fa62afcf1c13aa548150b8329c8d0e28a78dc30efa45cb2f2fe3810a2c9022dad30754bec41ced239006d27df38e2d9554acf5ea6a215c65add54d20d5ea2b03f18b6c9c6ebd62fb1682eedb441783e5cde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11e3baba00792cbec90ef6b5a35dc5853cf19ff4e36764fd0bd7bfa6f501b00ab1bccbdce10663eb609eb0c500a3d861c65a96ca0ca1d7e9997d299903e321d3a59c7501f20a0280a917f01d2d3926d24a336e4a3049dea477b9a3564b5837cdfdf3f6a1588983ad6b8b8c764fb4741202b264b3b7a21c9152a39a430b7bde4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d0da1842c4aafab783866bc7e7b3a3ea03cdf044bddf7f2328aa138b6d8d0f28708176fd1be05fb7fd9a595df327a62c73962717822504b7ef65289082dd04165d9161acdd92bf1fae2d845f7b8fc1466fcce468eaed0d751fed4c0bf4b99f638c0217752aa28a9630fc45e3ec312429b847e05baf0fb05b49cce2aed31ec29;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h573fe0bf6865453a0f93c93683cdbd1b9fef35c7181b05006411ed254bc1f52209beae7225e541ec521ef62b68c93ab1cf2cb69aa049a018a74937a8bd148e0f51f425ed6da5aef85e3137f255c3e80ea55949b92b9c4cf0ef8373e6f11d93a8b92921ed0fcfc3b2e321097dfebb3a297228509a97f67130f65aebc0b7e9fc01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29f184e7c776bf073ae303211629f1d97610aab69f13803985d7110d2122ec7d67f3cad4c9b313d8db006c980768da938d189b9dd7db76cae9f787ac4a621b127f22e6f88d9dd75fd319792abc402993c283accf56e244db313cec4a17cf8bd6779e4fb1e46db9e4672016936531b8e89a9a59f3981908649df6091878cbcadc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45027f739f98c42af5f86340f38c1321c4101e26b54b6d0230b0a582244daca821e950986955084277293376bd9a883fa05cad9c874543e96cc71366c846cc31c727c78ef1357bf412c18c2ead24c15932d1c2e6fb687b908ac589bdb8b9a54a38ffb641d4399bc67fdf71d0880b5112c760406adc11fa6fa90a4bfc5648ee52;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf83f89160222246d056a0e3e07f2b540870e0caf6b7a937a054c77c4cde9a2bbd58ec659dc1ff8355e9c82083ded8d904f78f5019faf71c20128ce512dd8695df7ca2ceb455c562dfb88872c320177f0e5537eb08b3eaa31e7f89d7e469f8b4588bfc692a32b9c3d17d14d095d247ac7fcf5434c1cb366b50b7676c8c80ff24b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f2fc4710779667b03a92283a885c518c6f69c87fd28d546d1b30411842e2dd9e33eb402119c3467f821048083a299840fe814fb4df225ecb454b49e1b945f275e63e788c8823da661facc8d1c24de4643a4e4c8bbab94f5431a1656e0ce89d1a0cd266953f5c4e8bb292c89be24b3c5683596aede91087f7ec6100bd8d353ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9f5ef77af8f5eaa0ffb64d58975109ec5facbc234571c19005a6d1a073e4eed883fe9d3e14d48634bd909593346030c17acbe79944d0d2b087bdd362a2ab8eb07102f30d5801e3faac1a76c99df5b086a6de0fb54d6fa5293186a2a6da33a26a1954a3ac8d2945613441b23f2c4b8b986b7d42b0b17728e4c4d40be4cda1d22;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4b56976baf34699d06d6bc3a9e5054d394ae2af5c4297e9e853c25fe76e0c1d2b7d1453633a255de746c9b0c8625576ec7db8050956e3ad60d46b336551ae0e5fc9b0a3ec4612ecea6eabbb57a7d649dcab782b483de801eeb3675f3ddb4d5d4d80e04032161467d9feaff79ab2cab5c328cf056e24dbb450aaca48333b986e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0cf0c670e5b148671941a958af03135e5557dfb8aeaa3e67e2d3dbfcf1cba06af88467f20fd9977b659bd2cfd0f56d3cd8aedcee0c55a628a9dbcbfccaa860daf5664b89122988707ebd48b57769bfe5a9e6564a0da8714f180dbc754f59d3ac90f442b5346c620708685595e073290991f6fe9614a0362d1595ef434a1d217;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h209fd3acdb44d81f979c2042cc3e34ab30979a8149b9fa0494eef866d7016d2341c82936fa3cbdbd74909a0ef09f901d614e4b25d5bbaa5d09b26d149971cdb8306a7be30f48e119d4cfbf10d7d1ec9f70077ff00d4d2696c579052b3e2b57aa9f16b5275854a5cfbaacd5b6270b462cad9c101209a088a2e28b3abf75dc05c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b6726701455226d7dc413dd3ae234d3dbd46a5cedaff9e95f4cc3d07725ab34856fbc8601f9e559f3e227d341584db8600e33b7ac36ba47a4b14dcf96675f1ba2d7273df11655bd7a5a336d93d63820347717de129f8583553c0982ab75ff21d3b58af6d75aab5d06ab8bb649afd995ed045b983ca4cbfeb6c5d29ca42ff505;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebeedcbce85c06fccb4ab513b199320297aafc52dcc14cebf2753b4a8d8ba371fdfbbb3a19f23abf88a3b3f19d36916ab39445899bc735c3f62adbfd14b51187c1b6fa0d3934283b89a996712ccd0f70fedaaef928277cebd694c1da7c9c922053c73031f10f2755a50537bdde81a274a3fe4e74d170ab68bbbf2a7faaacd011;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9ca22cd637c92d45165d441f72ac96232c09d9354c1b1420f1fa32ab8b1f7dc8078a8ad20ee0c60969362e563b5e69c6256a94ccbc72d4723a66810e73edfb24c7581b430ba964259b4f0a51a87f0877af516ddeb7f87c5ee18ef1bb4c79d8831316185236efbb5c0af500fcc0862aa4390de21d026c252aa1df01a58b9b7a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf878d6aa82af0d0ef44917963b32aa8b1bd8c6a409163924ed3f1c75c38a502743420c2c2117814e72edfcb1d1f427caf0c944ce1fc32809913b193a757143c329bf8e55a09adf40db913d3eb5e0b18cbe8747f2d3e639ae2567b7fc21e27552221998dee53ebbe6b9308ebf75cb0ca9968676fce0526caa3317bc42d9928402;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ff64af2a95af9aab739dafdeb3dc99f3870df6070b921b6b0807c429e8ae9f615cf9304e846eb4a92435dcb5eb412e206b2f3f3400e3b303ce1340ea7d60c96d011e3f1bc967b361f6b9427ff72b4492bf26c8be4385804711d59b3b36e334a039e29afdb12f5877511059ce0fb9cbfeed2308d2a6ed1896afaad61fafc122f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3bab650047a831e0d162ddf38f952322a296163c7b533938e12753dd6560a0e854dfb1c17269fe778e44934d96b6476d3c1aa6360d1893f10cf597d8a19e1ce832533f571860cd0e8530b65d6d1374ab0a5815235289c6f4d27bb63409191b778e2f17240c4e5a96ec15714f25561ceab39293b89e96d999063e0435b658d6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d2ccfa98233047346af85cd892f41e2fad38380b67b24fdd8c885211e0681a654deb0d431cbe1578a791e6325fef7b2a7d99f62ffcbe828760279d1af5e3b84d4020f88e3be7a9310ffc756444f6974846d71779f844901bf85a72274ffde452e686b78850b00458d0cf9bc97943e0a842f612f209e593787a8b65ad0c5f97e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2032a90e084c5564a5d1b9541440b05cae8f19fa5c3f80d8ea83446dd626cd8cac3590a8ff6d52ab4f538c0c487ac256267e63d8febc3d65459cd5ec11ad0808166ae6cf224dc7a40ca1fbae479fb5eee5e94494d371be9f1f0e3c296a494779ce8c08b61b30d3391c6dbf976fc42b165a159a1ff87c4f4c42b7fda7d94c043;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8af0be36e8c652e52db2b4eeaf48f86386a7c75c04734c2c8eef262ac3862d1bd5f6469d46554919f7ded07580e72f7b4735fd3d5d0edf4a1e5f336f8ff3dde26abfd107e0c8750cdad91fded8e8d1ed0afba6ba691eb0fbece53e324ab54f81b95a783067af4b0614f9f1768a068ae890704a1fd6ff97139202483c431372d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12c80573478180096d90b1b7842232d39cc91be65002bfa2fbebfef7ee06e080f9fe6c64bd19c77aa01d51d99c128648ea77119975d35c75772efb0bb821f6d1978589f75cf29a357d8b11c50a94d0f585b47ef1d564de838f09ce6d71dfbe2d106b30499b38a3559f36eeee1731973a1cac4f9473a0806a714ade3bb67bbac3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had6955e8a4901cf8154f7f6bc1da4f7cc9ea2b3baaa4fc9252c7c50639dd3617311fef01bdfca3b163c028e9b0c94d5916037a8344e965be53dc88ee1483ef6b66fb0c8223ef678991caf32625be238375b835352833d985c972b239b30fbd3bb778465631bedbf10b20d5e06f2fb51b5abb537c32ac05f4ee0093cd81e36f4c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc557fdb3aca7160a8a93af7eeabf37eac53f945eb713ac0f02b26fbc4e8eabe91e8db6a8893c8053103120418d7c8ec1bef4e60aad8b5578a272527823a82b38bd3080c7e10d5f2ffdadadbb6c531f5ad922f7f6d1619284eec90b7ec631b1b41a6d3254e061a4985b1df63ef59c492408223063de271d2f9dfb17e1f29f4ce8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce64e8ca5b085d223821cf8465d29e886861904e74e600e5122738d4daf9b5562b57179095f75a4f583877746c45f17a0b7cdbef2a1697b86be033ad9f5fd489f0eccc0a97a37a2c83352453e0ffb68a09dace52628c27f8429ae0041d9a61373f1362f21af40f6ac8e88e8f2ef13d9e489a355f8a72ce95657ef92e0c5a09c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce2e5038369719214741f31e9c1ffe2eb6ee0de1cad40c9d6f86c2c1df560b4e2b4bbdb9d7798ae3f5652a0ead19b3e6138f304afd9bf9be03c42a1df8de00d567e506e8c55d55eeaca50e4e5a8c85f01b7c37f5c02d525e475d25c4d034ac22b0fe4db9491a0ae29add360acf833d29c51224eb8025deaac7dd115518555bea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3dfc495114acc7250d0931231c7263e2102496d76b3cec2ab45e58b4887326d3d6231acca943ae03c2953be8e464efec0f82a71a17783932c7f1be5e8eefac9ff61b10c096275cc10a11913bceebaa41360eedfd9f1eadabc2b45461643ffa8783a3e2fd573e417815cb2b3a632b0f2380f27bd7cc9ce0e89693bfcd51482d10;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h146effe6ec936846ca23b7b342b3aee8a41e6a59bc5b9d8aa62577e00698f577c3f106772b63a22b50a24671f8eb39eaebb5549ec6edd93cd52a92394a10d13c27053e3c29aaeb1db568849f6fd304cf4d8b81ad0e4758c359721d78b628797eab928f2598898f8e97de14d3e825d245dd390b7072a2a4222e5b4e993da2fa55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha49773e2cf6ae2b60b0b581dfb821222571e97d189a23b5f8790450c9a19b116d122f9efcd6e6d8187d10a0c98b1dd531b908bc6d164d174d19e1aadd02ab1293fdd5fd1b75dfbda54f6bf2fa6263f97aa7601220966aa7c618281156388ae57daa9862a4ca0688d3516979f231d5324f5f629e1b071fd02a4fada533038c879;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc43a3293ae592bc649ec7cf3548c755cd61d7bb73c446bb756d0f7696b3479009980cba20cc306999b5ad7a201345fd273d91361a0476e51ad95c4a567151e17e826b924754b2d1667e7c1727c2184e4d8aa2b424f56d328d103956ee77c3eb50b1a7d956f03bbd18f9ee8b08e9f9d2472a7baf036c3db268189c5c6354c9ae4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacc46990dfa213ae3e834672c97c971b3b8354c22985633e75a21089a5b9f516974c956bc57841f10194f7db0cd6fc285710cfc666cb30845d12f3d3f9e3e88791d4e364a7cc1c541237699acd1bcbfb93355323f390387bde5d27dfae1110c233eed488c05ac61aa63fa3cc325e636e9ad6887e0409278bf70ce1510492f3ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h354068680a7251de0d214c575e8412bb7f2dc3f659288b906b586fedcae45b1f3a8c9bd8abbc4dedddec199f55f6d6f39231e3761bb84739601c6e877f6083eca3438738784d9a4f1572a0739da14a5f118b44ee7d35bc671801294e7481187d06a26a4cc08dff3bb8148f2ff407aae983f82c292f7853d03df81a9f5e08b68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13a5fcd956e221abb2735d4d50713cfc3c6bb1de8a603951d8a6b5254b7b2023658634561cf47959d0f830b837d6d11edadcae57ef2d658ae3e1cc31af6e98e23e6c0201374604a3101ecbbe8de109e2c56bea20e9a29acdc48d712be708ae99296e7061676c5ed9bf31b1e5ce1fbb3df496bacff8703549c58def993fc547a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2caa74bb6b2ad6e94225825f4a5738cf944e17f11aa45b29412eb3b007771f2e0dac4035a7132fa39c4abdf9bb0bcbc6f19dbacb7425f5d34b0efbbf711c71d96207c284b0d372e931e9c247abbb6e844ef47df170120400147f1993e5064a2cd835211ea05468074caee19751cbb1680403e79347070b408679492cc4f4942;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h452d98ffaa964c9daae73e4325a17cb1f177795073bba6198ed5fc2118b31956b1e5cbe085edd74972f98e3165d8fe8bb2f6615ca7f98ef937aec0d3381099ee871af1109e12fa8629da5ab3fdbefd58544184eac66aeae73f283ca23f4db849a228150fbcd7464ceb0be29e38f068e35013ebda2b8e71f4bf3ec70c6996478e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h770db8470617916f4b58f0b3253ea52d504d2fb57046c60bbf434292b3a585cfa56fb090064488bf436a80813c0eee7482abff23dc74f34dc58979ec6eb7d9ff5b4d37f561a8fa51cf9307390983688707c69b13f9b281670725e6d4840d27545f819068e5205adb1c87052d62b299a42fb5caadca002dcaa08cf956fc007621;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec7748b266c18a3b7a83bf98dd392bcedd07b9c05f046e773d05121c12089f38d0dcbebe00dec7cf7d2eb9c461dd7dfb42eb8aa9a555aae31ad49d36c701d661f290c63e54771ff5a56a796eae2e8412a086bb68c7bedaaa7b4701407be32c5f526b0c66a18847904f4f86034acffbd4eb27cce8e34f9ff48f44fa8887f908df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2800a0d18deccac75fc09914630e9d7dcba71d68aa751680324c7c0175d5543c38cf60b7142033f52c4e198a2022f3082dc1a4b303f866503e6f2a23e36995454803bbd77c3a4dc97683f6dcf8534617327798d10712bbc70c7d9b3bf2dd1d34ccc4698af6cd564b9b6ba57150425e1dfa4bc4f62d29e6513b3cfa5062b8973f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9071e65fa90f70621e401df578029253629247a388b31c1ab366e5d90414092e0b76e3792c8fe9740f49cf1f2862962cab53227a3b6d1238a2ef7a1be108075e1df5dac2133f4345891359f57614bd2447f43afc63085fb8a8afc6117d1cec503d1c571a47b04e1599650f1987f92fc5d404923875b55ae11040ae3239cdb231;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45757eb46da1dcdd04ffb96a14bd6ea56cadde91888643fa71228539b95b995f3e9f402e65f63f29f55bc760b2f5ebb37560ca5f5233551b0c285b7468cf0caca7377dbda1511987737fae6114241fcefaead922fd07054872242df67223407b38c24c75924f62b11c1fac88a9a3ee0cbac0ab981177da18127e82487d04ae26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdad33ca1d1d7743124c580ecc22b3a0c3a5d108555de0a767e697d775837a0dddf170aed65e11f0c766f457a1fb17419c37b9fe83051d8a78a48c56b542a848352ef2b92ce2f91894019cd0e6892833da7fed3db23c530b23455582d9346d537884ab9b2544facdd361368558b452ddffccc61aa287ff3a81573b8444665bb1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76672253619cb2b3812316b8cf9b086fe898737f9c6541d09d59cb614b30673cd169785e291c2f9e4b0d85aa1d04e3fba2c0c156d1549c630ac0b009a8ba3be3d9cf9a255ec75a47b4000b9497b5ddc1073dbd99c81f133c2b15e532ce9eb66143066971664b1309936805c3c1e1a75fea9cf18b6f015b6b23ec0adf9188fb0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37b19d07a521d82d09d4ab70505298d93256a73c9b94983b6fa56c6ad0319ebec8f829b2abb575800d19157b819352ce7aa30556ef4917211608f5fa965d39dc3f6edc2d39fe094a99da53335772d5d8fbdd9792ccb8bee23986245965c2b75ebb285dd4c797de84f7d9e036d4dd903a36c778e57644e3b35a384623829a0ee5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f99ce00ceac261a49d23ab1f2ad13fa014d1eedb4e743228deee1afe0548a5c785d7ec7856389ae9cb418409d95ed156d0fa1cd65556ff224350c641c20efaaecc211467b739fcb8c564f499f79002b98c9d65ca76f2df0a19f68abfcac27276e9ff94e0e981c57b8a41b8502fdd7c467ba285034e4ffd94b26cd0a3d70c4b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h759c73e251ebd2cb614f237560a0f32c564e8a45bb783f4f974c7e0c04d10daf57911356953ce29faf08c0f88a007fd3181d9ef0c6660d82c5858abb3aaf98b803854c5b4712c804def4265febdb5d8e35b2fcf1d6f1e6defa4f5af89b491bfd3627d80bf6a9deca122e9d3c38d1455476356478e9dac73b7d290fecf7dca55c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55cf4967faf35059295ee57500ffe5425f8b4fe288772a327530af211bd8a25dfb1b061487c25d85a393d3b5a37757504fb98645f21ff5eb4975aa9cb2599acdd8b3819de45193cdf418cccc424b8965df5a5b59f0b8409fac87d37f872722a77adb68633ca55df017d30ef1aa078251510a72d8c9cacb211f8b1be4c1c95e60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h128230863cb7153808eba83622b38dd0b7a002ac227a7613f3d78cc957b666521b6423e0facc7c1636936fcf06b0e60b450357336f803ba65c626c3add8032209a9828a91bcd4d20123fdc1b7f21bb9d9238aca3e94ac069911707989e83da3d6db55074099d6336000bf53e3521168a152baf77ba3e210929b188e9bb9cc934;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ac9670de65477f4dcac4549cb18de143fd9ba132a4284413fd2d541ab0b7935b009dceceb72085a7f42275cbf80998946ac982c98f0c2a680af28fd644285f8afcd18cb2e99804cd43cf8d58a341de4d5aa52aef284685b22dca71b1634e93c674570929fbe47ca8cfd199a3d08d6e063f93666ea97044e02324b489e09a038;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5846e7f6932c74ff3a58ddbbbef52677599a60b2be83af76c5f7ba05e47a3383d8f30c70d3204da73953810697ae04dc720cd3db52a88aba6f56a3d4ae800f83657cdd63ac4db77809aa088308f112846b23780ee543216ba32cdfe62d446ba6d674b8fb14c173da6b72ae60d6078f68ed8b7d2127c6e67b26e9931160cd27c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a5a0e9f3af3d1a8331825b42199d189ec56f360fd9d9d15373a49d7b93a31253c6555d0becd499bf77a937ab6a788afc3404b099aff5cf4c9871175b243bbd4f8132c8e6a82c91bb8fe68222faa2ebe31eaefa9d6b5a7d78179ac630b3fd2b022576a75fcc33e407c9a226aabb62ccb0fc754b94e7a5df2c13167153c3276d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36536aa87213ef31c6451f2879727731f85b7e25f8dfc6f997e7e1630504b6f3820310cfc97bd2063a9514af10c31d9a8790ac060acfffb9c9ad27b91b35ff3bf376dc2332e35f6a718399b50c77818fc04dc0b6a02aa86e859f57c89ba0b730ecdc08614dca9e6e2017e8456b4acba7e43bc7bf820694a215e6a5aa76c4aa15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ef37a6f480b244a37682e1f56f132e9ba0da608be39e02e38cbf41c2923efef9ecb180664483fbc9a535513bb8beeefa2ab14b43481b786c0b7b5b4a3b6bced31fd61dd6b7ce363b2d2e45e3390d94914eda20a2da0e1a94ae08e3319f58b8527cfc7648650f192d054cdbdeeee6ff9c7514a7d13c21f6a9fe66d5217f3feef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9b482581296142f188344975fcbfbe83c042d24da2289f6dba26dabc069e138a01cb09ed908e25dcc66799240119cde13caf9395a6f361f025bc88fcef61d2f5ff4b41e6e3a385efd7c9c1edfbff90d441bc0278791fc6d425cb589c3d435fe4e8cee92e6f982d0ca33c1c3ed3e0d1a697228648b08a23f883a6b8ebf378bb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d26ab918b840e4f99d1018a1dbb3d44077d28ce08e206125b1184b4ec84c69c5aebbd8bbd9c6cbfdfac85cf8e118e8dc8980cab850d76bb8c56d8d311a01b0510c31ae78d7e4b777359c0e3a5da913c03969dee67f5235af1d30f521dedd7ca4e1f4ef95e0a0a9d73a0f37947731c07d81c98343327b1c8a880798e54af23a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d1bce738d9c1d56ef5784534f67cb59caa3de249ac5d13d62881a756ee76cce195b4f9fc7a4531952c72c153112bc817b883e272f29cd2c9f235810cb4997ef2acc7ec5fc09bd8a8dcfde0a6c1f943a4e90d5f03934a068b381375e70efce85cb03c6a01cc3858a3fff3bc395300c883a1917a39cb49cb8b9522133a827e40f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd02fead5e2e9ec258bd8ff4519c0a85859b936ec2c023516e681759965389d1f0c4edd296882ea558cc2e1d64e83f3f316744c933a68efadb1fef601152f5bf6b7195a068f8a634267f11d164b67b9d892c43650ee0827e63fa62a48a17fa3acf0e723fbb6a052dc8db7aa1f733311a130c4e4049231ba31b0f640c2931d3db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63a317873f652b7330c21cb63bd4559500af4301d129eef9218d6b653f01a1333f7e7b014485fd7753dc2fae7d113a5dc1c6bc562648e54ec7eb937ee47e03f8bc480293c953441d1ef37e4e0ada8f194a89b194c12caeee7a2cafa7bbb787fb72f05a364a280cb700be4eae3a47a4cb63f3f4e58a3855fb466e76c694f8173a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf83b59ae0ebd3e9d4b7ceae675ee5f6cf5950cfbdc67480fccd6cf1ccc3d53e34e4dd4c2af7702e6bd0fc7c4031ce2b564189c1f307ad7e0c2ec9b204501b8c8e0917d001e5a97ef61337d219fa31e7917c9ce01c7eef059b04d136bc4fce39e32dcd5d1d2eb4acc129b9acff1ff16a4b0c6bbeaf9f51102e067d625ab7d40a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8303a93ac6df2f6b3b222f5e3688840e1d8ca059ceef03cb79e935e5f3a0aa6f16544defd220fa42f1c5567437d37ddefd2f8050c957e3a7fe20881630d6307061908ed24134dc1b3d79b1468ce24aed3c0fab941a2a9f6162cc5954518275182240d4d2ee7cd1bb9e6c111c3c510624a455409eb32eea46feeb2faad5749d87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66852e7c3c04676bad484ea3df3809e32de036a87cfaa33c5fe5b90c9ab0bac9b8075db4fe5c63b0829a3d647113a978ca4d5635f48f2eee464a6fcb0413814dd6fbbcc1e91d3b5e471e9f8a012158261a9304fa00178d07f435de54be6482519856e358b978cebcc9f6e337f0069b8e0dccdb54aa6efaab616c0114684194cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h409d224742d50769c061d85672ad1201a22366866e83a7958e8129111947af945882f59bb62f0801ae6d97fa41cf237f1cc50b47b617b829475b628525aa190a4f108008184faded059393b884d9c137a1fed777a6d878cfe8d21a313ee21e19f92b6aaefd66f8ecbe676b4e9f2e275c98dfaef831002c2ec82e958e1213e0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8ad7bede2fd6b6bae0e886b9953ad82eb801e58acf9bb0e1ece8c299f71e403fe4ef060421ad29bf8ba9be57c4853f1033108bc5f13caf773437f456f150fc0fd5c8d018edd716ea6dea0138ba3997455367533acce801398bfc8778f354bab0b2185a5d990f1f3b61a2e3db5ec6dc84944cdb9d8622bab85058fe0a74f9673;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a7d99e4f866fdb037fd2b88c1addad4722a677a636ccae25e02983c682a828abb9d2cce9655aa88840b1dfff299c97db87c49815118af03aed36ad07aeacd16cd32fd11c51601bbcbef1101d2170110c6231cb8d78a963ef374f8424b3b263228a1575f05d4f8e2878ac7aaed8bd5e1a0a789ad4d67ea47a589cf10a1bb1728;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab4a764d091c12157b76060089e581f2072157082b30bcdacc765ecfa8838edd814e0001a271d85a9e482f2c727dc760d608d540d42226e4f448f8df37e7fb84851dea98b76102f5d033191bd372d754fa927098e87c6ef1980fcad2237a12d9e2834c8b2eb37a67977f54229f8f9af775e42694692dd8f7fd2460bdb1cfe940;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45d3a399b463eb26e887687eb24ffd060385df53d87cedd3dd716c353a440583ad0d55b753b05fbde3deb91de4721ba576dc4942b84b372e1344bafca7ee90a27549d73003cf38eca2da3eba689f340f0257c6444bfc58cf8000e2321287114246baa70a2aa7e929c386091be35698c05dd3dc5f80ccacda193b308e4f7a47b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1d8ab910053b59dcf53de9e77f38c9ef8caf5da76beed5ed01279794e03e0361ff0ab4a94076dfe772386df7c9c41dc0d82f5ed8e3c74a3df446b37fc9183dd979143583052b8eb45e49bf1e47b556ce39e0448529d1054563161c303af9fa03f5654cf852bfcc498cb02f22789f9c19d909823ca6926d07e67bb8652209fe9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ce8da882eed3070afafcaef782b37c387411484a8c9a7c73c2dbe553eb61a94bee6497c44c3d0232b22bc3862dbafcd64d897b9fefd0940c6668d2e9ab30646e5766744a4e1e913728e170e2a2628c6bc8394c053530ca1aa15ace84b2d8603a753e99765e93f73ee258fd5ab7713763f8f6e1ea9b545f38631c6cee5922a03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8369d5e112e03ef43bca7ac4c3b5542cbed0fc65dfe31b7fc30f10821990f48caf55b72a4e5056d101810f77b3a94a7081751eca1d2c7bbd6918d3cfb22208e123ef8cb58f342aded0f7378589980c8feecb35aae822970c04d90df1a3e13a0b08ea3b402b9eef27cf2b2a441d634ad017d62e281cf8193dadaacd7eda53c37e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h278f82a820f83c0df5362b54f126712c198153f365e647804be3f8d0bab57e05e1f6a25d065c85b63f2d69d77060388f7cf4cd291d2bc51d2a9cefc8c64c19d2f49824c243a0c211044b0b132a9627cbf9f52a1fface61cfe961a95860e644a89df54622b0b0d569cee00ee326fb2c0d383daba30423c18c252327470c9985d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23709b32a3c73795d1d5fb5927c4189d85fd11868097a5ca0b4a94128bf6bac4734977434a9ed34c6c75106c8fbc14facf01ba9fdf2d9c43a9453a4cbf6c55fecd50103b04f19ec5302e526a8bcacaa3b893cc329e246fa359369dce245ad70075921cad2092bb6e2ead00610f6b9f14b81306a4583029ad2a4c7035fe4cd5f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47a1cf27b54b623e613a2c0e1f0d872ad8871dbbd61cef29d6a878e25cacab9f1c68d3effeda9e3604899c50e5928051998cb268f15d234d395dd44b943a1e295ce35af8115bc703a3969f05ccfe75ed4b93c7cab0203e15c17661d991b529b56454f231dfddf278a0b9f01b9ef2d44b610c3df8fe2e9e17a003c30a48af2a90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff481604334349b0b3be6a5b9fb5fc9bfe3c878dcdacbeccfaabd298168d9085c0479157dc60b586ea913617e5a0527ed39801a06d85ee5d2741e7428d17dc524d65c2e7d721af51ce6261d438038ecf437e142d9bab39267d606825ada5a3e10b6ecf87df2f0546b0a3dea4fdb472dc1833a604930151813ab917ba244fdcf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h177c8371eef4aea2b5c5dc7ff5b7f1868a27afe82eabe3732c36e1a968cf3274cfea8d7cd92979e2dfcd29df70cf2dfd2007a9184c6b063c30b86817d3362eeb0af59dd88544615f5717d169c8486458e3c4b8f7206db2874928e0d093d0b15487b31831540b57ee4a17b7e0cfb0178789c32c90fa25e1c7e60149c6d5eee918;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3f1b8e3b54263dcec526dd736b966368e32051fd3fbd747597e778832d2300e99465750710ddcf050dca8292a79fee75400028c4c14a56944484c1491a4bd51ab52f5c4529293ceea22066e7598679575666c588a184dc9772daed79f641002c89bdfe1baeb973708463b54aaed869a1e85d5139a27acc8fad8565888eb9c3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cf6300f22fea24ac43f9697c0bfd2e8d235694ea6c3c847714f3bb8ba9fb49258a86247f41e29946381065915e536e7f67ce3d3bdd9709de1010a5cbb1209ceb76e2ea23812c943ec03a387b71fa3086efb2e3f4f3ebfde93bb337159d1495314d9d2cc37e0b5f572bd8fceb9cfb8cbda76e0c5236686604c777fe159a21bcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cdf98f9d0e18ff915e009de4ffeb3c9590e2652a556057a930602f153af17c8d3adb5190d7126d65a4de5617dad83acf078fd8273bd531a718cead2faf6f7b019292557b6a7d1662cdf02ebe68cea4671759c984b8f663449146547adb0890cf95c9d6c0a2b5b89bf1b91c76e9b53be38666e8df6bf7c0dc4d9981b4722d610;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cccd29edf16a8e40ac18146fe4b4412258300e01bd4e54ee18f3b62f0dc3429dd141438005c2b46d09fe8c15bd49bb702b687bedefa73a90a0dce37071ee28d0fe6abd11df89f0412111b58cffba842cb7c21e580146e484e5952ec02c4ae0b9f0aaefa14a29992dc8ec7a293b573d82bf2b8fcd14aa5a75efe52926344a8a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cd35bc27f17d018f92d96d200e35c7793cb65972074095c6f09eb24cf371d2db042c23ead38accfc9f8085705897ccae576e6ce8c668f5ccaba26fb63de0a7a9d504adebd1bfbbc0d169cf9c37dbe929728b1cd33e11964735d903c0473d156e1dd8ba8f83acff871ebf1c83349846cb6e6a97318bd30e542938b8199d68fcc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h229f7f429bce715558a46aae683df5e9705e9c7621871e6615f0b89bbc3183d2e727dbf078bf277873f50246117bc30fdb0ab0dad9ece7a077bc86fe9c65ff31718e662a658eef4bee7e69e63a77eb402fda0074478aa3f15ef7b44569ebd3aa2dfba6615b702ec264a7a9da35f3deafe3ace1c79d7f007a9cd77e6e0d6da168;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47cd3fddc9d4e853d56343890c2c973a04ea33915cc19a28d178c2fdc9eecdbff1b2e2748c1b3c15f84de53774424b2e77f4d91f1b6f4901d9ce738fb56f735ef5a845b59b5a68816e3c3300b15514719c5671fa5c6b9ee907f778286e93523f6a50dda95b7f10b6b51b068d897daa3715eb632ee5506db552aa158f6d9d582f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd922815d2c2e2266031b5f12f7fac4414ec5d27d927ebc90f2048bb2c4343efb4e853ab9c939d13b6a349f066b8661ebab96cb2cb7374cbafd1075c324cf4c1f03c5c399f9c463560f01c6603554bdd4ad3b38e5356186186fd0c5407aa10ce57ffe0573949e068cfa7cfd8cbf2c5c46e16593bab3095854a925dc5823a789c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65a8cf2754ffee569ef8cbd38100a9b06a75a05f677af899ebc73725d4b01dd00c5853fdefb3795b07e8827735c6d33fc7e77c523e2c6fde542cdb6174d436adefe463c208db1e148d5c9d9e83006b921f4d1e487cb370586b22c27e3071a8110e00d8e51d19e07622a49bd34312102e5723a51241e01a8c62223385c11c4b8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28f56601d045309b444b0c2d073535f389310318ab7abaa40fcb4b53f1103f1879ccfc86b23ba6d0cfdeb72afdcb82b6eb60f395a2cc54538837d3713d99c0ade30f21cabf4e8c3579d91f703d857be511793f8db754cdfdd6bba5bec536dc08d9492a95f089145a079482070739e8aa5a2a1c814e60d7cc5950792958079580;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee91718dd90aa19d5bac907a42aa4774cc2a77f34edbe6dfdb6f2c44c3ba8f23eb43b68bb195941889e8888b11c58b1f25037cd200a5d0ee40a84d1828d4b56c37d4a892310455c1e401b7e9a6a0a677b27637f9e3368254fda109f8a6beff670242c2b57dddbb83d6b8c4ff07636a9363b9c33486446ac70d36563d1362730c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95d5649d6b296ff060b0f8b8b67710467317e47be6573c0cb6776e8898055056c9197dd331d1b921acf5d02c0543ae3b17cb23a3a7497f7cc5a20ebf32a0b5645d1fead4ad582f77a8ae6980e32f154c44235ab65d3d6da8441232adc2708f649fe0de02e01972d5934e95b6d2ebbffa6efe9c7dccb74091078845787c29c32b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fc0e5c1c91e4d32459cc7d47bde98bc01158511c70782927ee49151e68e50f0d78aa4487e5186a10d1710ed4d48dbf4cd9ab5b282506caa9a91f37c934106d171e22ff59abab1cea9a9780ec09548b88ecf067456accea31609a3813ddb47ca3e0f19d1d39229d8111a12ff874d96c4f9287252e24577ae4e55e4565b61f16e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71e185a4e366c61fd80ab0834d339bf58362a6f390acbdac2a4ca37b523914e4070c92fe5060c719bc7789a4da6ac257aaefacc9b36b8410828c4eccbc5bc3b3d69db91be039f42f32e7cd3a046e2d50a2f19715c0ceff9f53b713edf2701ad4384253fa1326acf3e10a16efa6e2914d8a21bd50acb6cbb9ecb2210b5c3280f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae48f2de399009866e855a856b3b344ed15ae9cd0ea9c9c06cd8aa2bd4d34c79e1397336e2ba999d3fcdaac883cf4e2370d4f20f8423ec82cef992310dcb929eac98b13ece84a1cfd8fff7c6506a347d22a53c214bc09ae020b2dde7baf78800d02a6f8dcee451f4df0b4063f5bcd1609c54c4010ae380de62f3a9a83fd6b4f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h382380b15c0c949f324887becc6094d4b843f04b9f37aee7f357db7045b8ad82d0bdfc7ad89d4cc38bc4754807883ea655d19eb15dfb6f6553bc154b61c1af5e6259d4158bb271ff79e5981d5bde09b3f811068a5d598e5eb8960b8461d25c421a5d392fd16e7bd80d61e84995c68104df93167ec056d42cd5ab49c89e75bbbc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46512b4f925bccb23f1fc0670bc27c3cfacc39e981a232b5bbbfcb3ec25247e1927b05d28b7557a4792d49e46d2cc26c1bcb37f0d54d83866c8c002fe9ad43d451ae19338f56c75010f5d1c97d797bdd154a7bcd008607b45dba761ba73527657151e960a1f0bd5530fef123b126be5df3d49c69465e8b766ae2e4cd7787aa37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b981ca0b5883a6145f87b5e9b83a07ac3c46a0d6063da3ca43facb9930ed4eeb6465c54fbd6ca4e451bc56a6635c1cb2991705ec28ea5f0bb92592e6382f9dfd616e61b9d5a42cc6f06385d8c2086f15809f92a4910f323ea394ca089645a1f5c9a015f33dfb4b63ca228ce4cebcb3f8834956e183c22eb16aba743dbea6c21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc3f5ceb098823be7720fc6858d6e181431f6ba999609acd40b47c665d66119366fde7e4b921c84541f7bea65e7ef41ad6a4ae814ee029d2c6e3149cba734db906cec0cd5b5e57791b64417eb35324653fd08e2c8c469c24495cc6a8d55f6bfb287905bf576072f45850bce8c59c528e28d731d926d1b8010495eb31fe50ef01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7602369aa8edd7acc68e059d0a2f493e7dace7367b644eb44e7c5ec053359bbb53838e94f303d39fa337cfbf710c1a3f02f311a846f229a6a358eafbcc746e1a1695adccfe9ad40e4843c800b6e1a7892a5d2c675202c6ebc3515ccb0c63c111f8a8b03d9c60930a7df3d628d35834b979b0d46511a9cf5444cd0f06208ba954;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44d87142e29ce8a6a3820799f19364a17b649ce6b0309cf9ac8475a3468bc41543869cbfc76f80b7935a389f00dd761ecc9a76e3f2d68d1328cdf1eafb83fe054b42c929cbb6ee12229fdf59eb8e072973104ec23cb25eb10005d94d5de22d64874510af12c7327fa7681c069e542e9be330a70e0a8f11c4307006c590f3b1dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35431e86b2a5590a63d349e1170f046505a351bea677aae40461a3e067f2bb7f25b5f8fc1723459357547d125dad8765a8ec35e13b33c09fbe30af1df36f9ee2aab2817f3645389df686b0d04d5cc243a40b08617c0556fd10ae3b13a67e4c2a9bd1c66743583f00b63e7006dfb11b69fe6182bdba7bddb424297ef61c7207c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49349691629e9562b5461bfa76ecf034dffabff0ec45dba2183762b9def369fdaf81cbcf54800c9ec1d4c6c603b4aac44efa77c5dba0da50281717256333889c8c0bbe52bf95dfb5a3a7816d9b028c9cd7a378aa11c4d3a2c6690ec61f9dc67aaa4026ee7853439df60f2ed775ad6ceb690218fb63f06877978f6f317b7eb0a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h365aea3175f34e67b81ec6351b724896a11c1d6b76948f5e401058e4168c2e8350cb01a74cd8dbe3667bed21010a959ca50c500171e7d9869ff60f2909a5ecda885dc4f177a987d3b2169cf92a3b7b2be2856e97284bc55da85a4ddaf8646f94ad016f2c5c49be42bfeed03faf374dc6578ebb34a71689dcfa410c506287afe4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he613aca1ca871baacda5f00a31b5290143e5436235a64385595fba3c3e97d6333f0ad59c333cd68aa7e09195e1c63f2c15f36ad281c399639baa5464d2b3fd23f472ee968ce88d55367a9db9c881ec5013d6b9f378b96f7d6d0994a3e51666aef0a8ac57ffaedab20cb50a50168cb9cbce8d5dc7fd064a28b3ac709dd8310038;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha65e0ba094d3d1118c8a8b03964725c33bb5125e039e23ba03aaeb7094b488b97d5fd5b95139f03e0f1d16f356fbb78fcb1e9f73c299a4e82d51897018cd816315b83a48e249ee4e2e21b7dcfe6f296244290822921422f98ef4d6bd6c38727c09e2a4cbc8b5805a2b3d3c07a226c7c0a1bc54e1b8b92ba938244bace4538f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65e85ee1e84be69ae509d65ff00d6d7037816d0c8b3ebe86344a07d29e17b4a31d5c00cb444c3703bfdf9e5ccca1b4403191b472708e76eb70dd3a050e270fec21e3b49184af759cc12ad103fac132ff75493bbd75e4da3c24a214ab2716b40bf5e133dff695cab8c88ff0925b6dc4a97e7382c0d6a2f7e7b8d573b2109a8f46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd90fb89dfb2cfb2a72eafa4bc76287a56cc666801555e7c9c059b5073d3d0d1fe51d08f0c87d0ff99bbdf45f59a334ca4030d16f48cdb52f502d41b939a95bf5af4f8a3fc21bd2b9f6f9aa12a17804b68ba2cd81293d750f022735fbd929c9713bbc297cae128482151afae655b3382291244e01f457ccd34e27e6ca801ba366;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63d1ecd124775a5472fa57d42ad8a10096ec5c798c9c72c9be616ebc92c0908788a983dbd72b17b1c4570cf4eeaf05976c1becca0d900a39b10426bb3d86ecc76a46d1b4635487b56c53c763b33023dba4b1ce48e27a8092321db4afd8094e17c9674a4b973147d33a51afed98895690125b9817a90639bd494bb49b3678ac21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9f23bd686625c04e25d2664b6c0ac59485b1a0575f90cd79e411d6020f4626b4f11954babe7f06c68c76f9f97de59c1e7ad2d27d8d184a20a38eb62352060e91ddba7faa6288bb9808ff0d2797dfbd9a000022e7307c48aaf48d6f4a6c5162c27e1330bfc92872b12272cd0593cf20c3ff1616a1a4b00a3342dc2e3191ee2b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53f7443eb537716e2c76f7d6b6dd4a1a733c50c676973581d6a263109451cbec092123643fee21bee0b4b1de9148af068922c26033bf2a126104c89262ebcf34370a1e99d496daa541f9f8462ea16ad6fec6c42498804a5c70a8efe8610a4fb7f8a5d74874c1bed10962223dfdd2ebcd735d70544004a000c5ef5a088e98782f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55d64afa9312b91e65269f44f9dbb80ea4fa433aab86debe624fd2960c680652e8e55b88b32ea7239bd6499d2ac93698ff2c5abdd9271606ab52ca68a2b5c11a18ba4aaf4167731dc30c123cd4b414b8c9ff366aea0bce0042df34c737ae322cbd422f80d854cba217285d5270c254f0b864314ae3f48c746b2b51bf540d0515;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd14a31e2d3f8789ef544b5e22fca2266d0f44d1652d2f4d52f1f0ea01655f2abf25ccc8c97da317afa8794562ab62a921c3f12d9dfc1f0fece758d1b839c5c119ab572520180146086f553d2755f004c788affe950eeaa2615c1018c4b19bfe1344c7600c997b88dc66e380c3d180467846e6ce0fe9ef0a6a58c6051d3645a48;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17fe0b644d7caaabb5d279b66e715381fde99d61077a5d07fdaabcd5a021c90cd1ab1ac494cb544ebac457b58d8745c62df7f214437fdc482c160efcbd8c4a4f46cbc3258e6cc7857f781a4cbab6d02012cdda5777977f47aa63d6be06014975995f5407de327433f46f738acda40748ede2454a95de4ce6db88eedc6b456176;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89ab9efdd9717cf6142397ca3c6b4f52efd2e44bf8292cea719dceec7363700d0ac1ad6c109ad3b57c7423b2cfd7a7ae2fdf6243810249e298cc7d25dfd39638bb5d297412f691c8f7d0a883faeba2a3d666ea3266a45f6e4d598a01c914890acd20c49fddab2c28fb1be99c82023ad2fcfafb2c69a3156d5676c14ed09e5534;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4577d97b063acfdda5ab9a9b7863d499d526930cc2e64738ed641e331013b5b56cf8832423b70efc15c606352fe3d3ad8f43886c06a7fe1df3e084e1b2dfa4e5250ea076135669ff673470b5d7db8023febb7a338cc72887cb0c33b083f67d4554669502e42fa08ad258087c0f68682e7e82a10f6d05410450ff11e768312816;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95b5df5b09a2ac13c5cb63636013b12caa3ff746b1cf4c63a07d01e8eedd9eb8bc6a142915cadd957e14a0e1373c9b10e7fb9be84615184dbc4590a50dc0228004e4a7ffaba897932dea377e3619a5b02fd400f9c7ecc2557c291c2a00799cd832a478ff9e011824c2d0cdcff502ecff313ac69730700e251873e471731b6977;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he31b0f46f800ad28070c8b1917de6bed41bba9515ac28c7458310d73cbd3502f836ad2b771362f955cf54a6a378f3fe4dddfda226249b3c044b6a4fbc2d116413ea38a82119ffa94066897a349f5e8be85b50142b43a053fff54edb7c3c986916c4f11281c5e099311add1cf28f5c89a868718227f248dd593ee750a3b07c75b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe6d629d57ca8c65f39894fe05fbfe9f6e0ca55c0bf837e31134f96502d3496e689a4d3e86b2528cbb08d9349ea112a18ce82a49d91121fd60c425d9b3fd3f307c9651257ca41bb9138398bef1b6ce3a5bd4b60098e2e549a959578c9a3b729672d189592aec918b903bb09e39d67bdbf1e3bfae9a5a91a76f52b09b332cee0f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7440b114f84a266f1248b4ac2eb43d3504ecd9af9972deddb6a8862dabac70f9adee61d75f354a26a7f3771a32a8b2b18379dfdb4c3b98297bc8bf428c65ba70c81388020c77128cab7558b6fb72cc8c539314d188635e5b141fb7a75092de206ccf1fa206f835cb7dc76d8c6764d38c5ba65be41295a5bfdb91de3d59233d40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49f2366ecfd784e8507b362ce41c55531a934ab9645d79e885a468cc6a5de967b397f28df0f4fa185d14c4dcc319d0fb5b260750434df350c24fdbdb1c92537c847641820072457a6706d373a2f3bfb6f0794f28c554ebfbf0bbea74216f6bbd02c9af9b0a50e3e370fbb78f92e0e5bbdc576634086440d7b90d5317df153bdc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb11da133d6690f0dde50cfae720cd78005972deb192714ffd292f4a8f7e103bc6a35ed0a40d5cae23e2467335694c5b1401ce3874526a488815e42aaf81aa357f069df1c5487fdf3ee6b3779927d3cc61966e6e0071a52d981d488cc26c5f00399e433abca63c05f0c67cfa383ea4f7f0eda5bd4e7d2a7c292bb13c70e0c61c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50f8f6fe5bc188dce2f3a5b2002315b448a58618bcf5bb2bcd76d643f9c59d2cb3d9c53d4a76e82bad6e13a7ad7e09bd0bb3100e31cfe960906df4cb3c120f4e2f30c6e1d0c049567069fef0ce527e36b59c78e8101d8c951a01363be366c5659abe8ae9c0becc09745d454691da23daa2b96890c87c3ea00b62f7efae5e3b01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8d7c4ac016d833706caaf1ec042603607e8086114aa4b4981f48ee370585ec482c88347733f2d81dab7d4e7c5b2fb449b93482db3cc5230be0b9639315d8e2dc7b22b98a8d6cf5882ce76aae6279790e275f2838b814163445e0e60e03c78726efce0c5d110280455e781d58bb36968a81423e9513d5b206075729833dbdc1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b708006459e44ee2aaf12ab039a43d51798811184b9d535e1187cb84b9139f2f3cc3fe9158f51e2883ccf986c5a064c41ca97a689da222d065c768ba3db70460bf3d71a5489a149f8af775bba0db82ff7494120274fc3b8875efd86b0082469de2d10839ce982105ad132a3080f316288bc92c504f25622a574dc7f51d9364e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d3efd3243124e13c14aa1c43f01f71dd0109f8c7127b206628e63803395490488e672b9dedc6f55d6ce46903154d40b81cac3295550c15566579353a8d8df50296e2d67bed75705f8b4e69cb87bcbede75afb35183139bc6603bfb7f9075b5e2789f0fb07902459547112da989f4f32125edbbbf4bec784ff252cad3571cc02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd69c635edac0155fa3b36bdb7e33348b59cef8dd38d3ce4a75d4305abe08582dfe3dc02df303c32e4113b73061a36fa38fdc4c5eb054c5aa2a029ce2ce5235864d51b697b65b1a67c4341bf42ebfcc3bd739ee7a3821aba126462d2f9fe8d77f2cb8b557ed8ed29df72c8864f4dd0a6ae3649fc0952bbc8aa17b32d13a2d03d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc95595bd0fdc8b2578cc0d735e597a3736876cbdd6409aec673ec4fb63330b8fe12366cb34b48d1f62db9a52ddb01c03b4b68205a7085503d1dd962b2a54de093940962f98150214f8f5e188a1baf4165d9d872e0f2caf85adfacce942fe713f63988c592bacceec40fd77b732625d2573ef97f86d53950982a7b93c7499c7e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha47ee5cf577745ce5b335ecb15ab206835575f57f36202a59bbae151a4fa594efef0cd3f370d2478afaeb28add080f14f4f3a173a4cb6cde4c945ccdb4135ff070e186dc164897da86f81d67c19a4c447f32b6ab5a1f8090b449218be6fbf000bce6a191c362b18020d1506d9a6f291ad3187b37f1aa4df5f309928f69bde19e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8998825215e2c5b71684d52330296f629e7df84aa4d2b35f749d609562fc3ff0ab34e5fbbae455998ff2078a8c4d83f6f573568062418ac8ea1fc668b8635282fba562dfcdc7a72a159928b9105acf8240cf124c593d28bc6b0466d205c4f52190b6772f9f398e80b29bbde96776805980e35e936af210085815132e5e071d67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbd829b65fb2facd8dabb3df6f473d33b5972c9e44e5d6e1096dc1bacfc2f2f277286f67eff08782eb5cd6b2871faaa807f627404f7ccf4db596c9ab328900a49dd40357b7b26800bdf285c60fcd645cd82c9a02af5305e415c6ae7ded2d44be80fa8399c14dce524d4613f65c8d56ede1e4d5413aefc03f21e5cca173dfae89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6df97a06270f996d452148f5624d1e4b1c4978d7dd5dd3f094094fa1bf2bc48f94864e3ceec67df2ab90e2311b72fe516b06c4f6602ae6f65ccb10dd9ceb94b9646e2fcb1e432794680f3eb692a664febfa663a3a60912358e28afed8dd02f2130af25a7f773acb64f6d79fe860e0e4ea4ff91ebeb6c0782e0e91b2202fe115a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e824cdb3eb4ee0b1c49005385b6293501a6eeae31b15428f7d29debbf4549f8014568434123fbb18c653fadca079bec3577786846d1923f59862acaf632f06306eaa6ef3752952c0692043cafd86d84d77f0ca361424ce2eb4689bf3ce5a9882e77a0b717e2a20d22e82cb51277b5dd71383125924eb0375bf198271d38e848;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5effae3f797273fba705b261d3b573d8a1ad41be6547bbccdf5f1a59ac384ab693bef17ad43905f94bfb71c50b8a2e2da2b0438ca62951ccc9fa84cc4b2ad407fd2bffcea06a93d7f76c68d67960b8583628ffb25a8a953ad098024891e6ff56300b3fde263d3b7e5f64e09b29cb93640f71b4733eeac919d2c3923151f29ad9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h995c122f49624c3152629bf8a2f6719594a33e8266b74b4e0e951540c68f59ce965f29c142bc3625be8e27dd7aa1e520a78a50466fff64ddbd65cb29162518f1ecb7564c80c8597b33ef9e92f8c08aa63e3e231779b4bfcd3c64c2afe50846b4458867e789f3d0d7ce180c3b1ad90bba9e1be3bc586b8241186fe0c20be1c1bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he044069b614a1ea667e5842f1a88a5ada7b20ae9e85d34535a313c8620b63c1255bcce6cccd18d97f85fcb59c9bfaef6d29e54f54eb839ef8cc26ed55bdac634d0764445ea51f35f5ce90a3b3ab03539164f2911c800efe98249905b3fa632eb06959421926483f32e2593750034a4bac79d0201ed0fc32864a9cf4622bf6825;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67a06989d47258025ee1a77846d57b7325dbb5342a4441136a4bc98fac50db0d01b9012a3a63e00a2d36a1438fd623427b661f15fc924fb45677c24cf3a7783809e7e951c35fe5fce575d3f72028b0618d66bc10aac44af00258021246c2241e4b14e89420346d46dcc2cc8c80d1bde9a4aafd27263abaeb3a669afefe8d6605;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd570fd2f880c0db0bd9fa6b88bffbddeed905171705e4af1f5719b6b7a0b8dcc249258ff4fe6895f15f3fc6c44ea1dac8094b5f8a4e1f30329e5b6c5cdee71abcad6ea50de5a0c90092e962a919bdb8b6dfcc088cf9149eb63e72aef8e07be0aa42f5dbcae78aa30a9ab6c4eec3bc89977dac1e82bfd3bbfd95850282567e03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had9840b6dbcadcef35c73da6aec666b8493f72f0c1ac0f06fdd8ce9d13d90042d308df2cb0eea66991589b6455b6b32f3c4c8401c375003982d7e5e855b4d13d299bd2999b807fa50a115d6deac15de654256661df8e4e002c3b9ed2fb914e22e2457b262ac14cbf49d3e2d2c1f3e92c7b6423d2d2dbfaf50ca69f84d86dc327;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h155e1892ca9cb860ebc446ce9cb391a2c6bdb3f616b571d4819deee4f28ebbe1e8b0353eafc755614fac826f13309cb0e8fbf55e97e179c9b2142ae8f325af1453a1f6c4eedf50f78c07f52103499fcba27b2e8bef0c979ffcb205684fc4b3c586ec89a96bc3c9f16110b143e6540228af39530a2a4cf89e08331972780d3b52;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4a1fb2719cdf71e428fc80dbbc3ac8c09a4563d17959c51676a9cb8600d876841bab940685a1f4e8a6452932981eafdac7fc8e7f5c1f5d68b83a3928a943b0bb34ee2d010c2f3ffd9a60da881b71a530967bfe11f02fdf6d3d700d9c5f8589b280a33c97ad59b7d2912ba5eb2de757124d1ca9ccb0c8637b33b6d4f11afac64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7e9596113d89e12331fb7e929134b376f88dfbc31ed06e3885a6af1f8fa939a2878c580b579014bff5106b91a27f10e71f6966ba9208508e2a076277c1cbd3f550acd24037e3b4d5f3e0b2931b35dc4da2214b1e12bcbecf3793a65c9c5386883942bfd29a0fcd49ff487ef8d2630243068548b20899474b92d031fea460c05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b214af277f07a28beade957c95bc0e871d557dfc64cdfb3a41a7d16220a9f3b31257b747fe52d7ed901265f38719ac8e9e146ef8ebe47bfa79830d562ec1f538ef863ad3ca0a12a49123b426567bdc54ded6a8d9c3b8fb05739efa68be1fbebcfd25440acb81300cc203ccbae4aad2590e7d6add3ed51f6af38ffa8574f5ca0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6c9cbe883dce37362c6809380dfd1c8cdd4e9d69cd623d349d80de671a89bef8a81b0c4254954822d1795d06eb73d6cc4bfcd5261bec69330c02206f47b6a976f88b60eed2146a4dcbcb118b386ec2c707a8a3ad14361b964f70a2180bed70b72a5e9e06cc7f29b0173913f9e47d1922792ad7b5d3ee61c4ef6767d25acee5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27a3d63e07f92a932f26a850f10790079624a97d7ec686eac4588d0a413dda038b5d98fbaeee4dc1904c4d067e7c923a597e0f54d4c46c09febbe21ab965316e797be72240650f8b56b32cb36056e6f0d90e122512ea394d994d3c244901d3f73104e178a6133f1eb09c84150dbadb1b36b4e6f738594b80325d294a4d268855;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67c670dcd62f2178da2932371c0d6805a1a90624d6d62deb22b5ea97f8956e305b713cd272f070a10764cece121f37ecc625d94d49e5897402a0a410488f677827d9ebe0d5587e7a0f9a923b1e32a5dd8cd786f03803ebde024fd12c50287798f07b068719f6b0b15f6770215c7e0484a231e5bae339d16819fed325c8279bf8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25c5553a65a7f93615fa8624451e2a4e7c8ec0aed7e85cc593b5198d707b7c8ce6bfe99a6e00053887b65968accb1410b16f050a82c5f4c5d71357346dd82abbe603f74e4298543b1cca9e3fdaa1edf8947d9737dc19453ada66cc07a29257cadd054f971abeaa8981581fc0993d919749e2587ed6e5c9e4c837f6c874a3e6e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68660959a5d24f7f212c28c09d64fc80b41d0d18c4ad5afc09984b2900f00cc816fdb49ea7410cfbba669a1c903767c8d8c12dbf2bb0f6d03e1b12442da2097488fbf447b280d1057f054c5dd4fe68f224a363dae8b4a9d2ae796a6790046554b3deee6c97be59d15292d606df647be97e73e01aaa8e5a6564b8fcacd01165cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d979e72fc53f8f4dbe113b2c49c1c80c76a31fe5e7ee36f2914b75af47c28afb14d45129441c9b8d5660825ee0f3dbd86fe6222e9001874c515bcb34a28ea0c34b9396874aff3835a0b5abe546e711102352932a003b19e2df085086ce57941861facb87356865617ee03417376a07966c3c461693d1844c056ac330fffbe32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heef3e50c67189eeaded79d57db497912674d83f07a60a2b50e8a956592580c19ed69b29eb95ffe473b241c8c9e1bcecaa6d1162227333e5096691aaddfef6da126ccf3c37905dab5a41ff398ae7294334121a6fb0870dd2ab651f5003435e25ad6685e7c39da4ae75839f2c3347660f9b9238fa85fa6fd323a3196921e98ba94;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had7efce646da7bbef2ac9188f6cf0df1a493c85fa09500da0c9f923a2ee51b72fb32110c3927c5d6e89042d5f1da9997d66b923f4575098158b6115239dd2624b976a8d53202cbdee067ba21c1de390487fcafbdc7e345c8b43a2fbde4f126b20aefcb25c5fe20edf64bda2e598437cbdff1877c32754124d3e42a5b56eda379;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4794118ca0bc0a0ae9f4c823c088e2ddfd49f8c55c8704a203dd1f5a633c5f759bf98e52707202250757d45b9ebd7acab98dfc9f5272d67f4927aa8185d0f589023359682b73fe5e5e5e96c1099021ce688138d4da27f9c286f0cd800219a22b5c2dac2ecb4327a757bdde22b3460e5aaea46ac6eb649980ef4f74007fe3641;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d79a85ead55bd646fef4703976310dca0d4c5b90642ce04cc1213e4cfe1482c8b63c839dec15588ad63bd7bca4b888492999ef49e577bf16ea2d39f4cd5d78e99e4a153e6bbe7279be2ccff43e5672bc72b3e21d4860172c620d0c701109daf4ef2faee427a1093ecff373fb61447a43b02e82cdd358658b0a0f58281396633;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd883623475a058bc5fe02248a336169bceaa8477280f2ae20ee82806a00c2705010a3841ebb12e2b09016507a47122748ef5910b2d4d63b2a924e64ac41a8da9b54e8d57b573e768cc894eb970e465d14fc3c1409b2d59a688d8f1e068d8b0b50ca57de9fc7e553fed484ad6ca052ed4ac92b765f13e80af33774c17741bcae4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he31caff859154a180b1025e63a5d2c43c9447a1891061a5d5d74ce289ac09754ba84be00d43707a78a0d18189b31b36ebaa8c47fb16bad3574fde280b3b22ed2d7b312370ee5901886efa692f7a5e92cd8dbe52cfccbb421706200ca26931f0595781aafe7fd46766285492c6433506adc5a6487accee3d5b8b8c3482977830;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha54a58213ea7e180e0921e6e1694723fcc64479b636d5d86784d3438ea3b43cae508d325152880121348da3a10cc40c4af275f1a0c9f0a5ff65f709b8fa9f3744b9d036137a9be01e7cdf474ffd89d19095ffa309d0b573ab7f7ae7dacced00f7202d3ba46b9ebf81a99c2cda19d4b99e3e79dcd2769d6cc4b8d3a54b0f9a16d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b749ab445ba83e085dbe10930bbf131bfd97827f53f17336857bbd583a0b9b3dc7596e64ed148039d360cd115c92d320b5c9b7af78b605f58f8ff8264c14e5a38a34aeaa6df148a3e0b4bd63e8d9e9d77977c09d952a7f3c4137d6ccb2fdf19d690eceab048018a8b26f9aeca442703c717a579bea09bfc4dddfea2e277079e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hddbeb77e09c439f1316899209540c974e579e3dc908e7e9398777e25b85029f7beb72fce5735a800f2abc1815fa64efabc321ceb9f140037d49f27ddb954f2ded16b5c2a7eb955b1f1c72fe8692ea2d19ee73960b9cbb523c7c4045d3426f4a849672f595ecf3df60c6aa505574d2afb6b240c0606ccbf05772ddf8f8744e308;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50b7c4833e96b1a53d4992181d4a21931913362edc5f6f0433c1c7692dd1df6075ae77463820e59e49e40f752e6f4d1d199ca43d0a95a29f8483540ac2914e324c0445a307f334085e2be36805d0651f2489e989aaee2f8d03ffd5f42962d7c159edf83368356fc85d7b5030157776b0a91c3320d44b93f8bce0cb51a244667d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ad8271cac9b974552a5a8810ab78b93e138f1941b9d4a2e7ef039c98eabd0341a18a6e3ecf7b73f896107f9ff9eea6d8ceb391f5e923a8c40947eef8a63045b630f2c03dda2fcbcbdfec831ada16ff7b63e8d658fb3d48b8aaf4b49b1e398a6f8e7854ad05625a45bcba6128a97192488539ad11b3d3fa337765fd8b3c80816;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0915cda2b5e200a1bc0345e91c4031f827d1a40e406c78eed1cdd69dd813d3eed27b404d841ff5bef0202120aeaef37b96dd42f3016aa0164bf2f8c79638dbefd917e167c5f341c63e50dc4a2f364cd705fdb7693d8b01363842de99529eb44a7d6d5cf6e1adfe0fd9c316177cb55b09cef61eab99a5eeacfdd589ea1883139;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd05e3e45d4c5ebb35bf11375adaa5388a1df34073b7e4b1c90d8d8f7db8e159c3e65b6fd8343907c3be35c373f716bee70985fc5e3d8e08729cc7790973bb16de2c38c3b94fc3c082537920a84a2fb3431f5d18c9c8ca7ec88593ce4569cf2bff44f8563f0f9ce4dbe90c3bc420cf15960ea762c1503f3f9422746ec0ff7d3e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3731de3ce0699887d9e6f97c9475e15da867ec516291eaa207d01f59b69d32830646bcd36cb26c4a9c639c7c32832fbda3064aed8b6aa673bcba28f15ee8608a58e0d37d134304545ce1561d467ad1d26c7d028468331b09064770e7440f2e31d04dc651ddc223fbdf948d535c1de260829d647d3ce179ec0863f027435686af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc2be0b935ab25db9448be9b1a514ae0b664e2e6c164b93e0789839bde8fe375b80abeec602f0834a49d77d5a926943bd233f3092d24f20d0480d1f05d6c1d2875c0488e0b8843ed3a85cb5d38445d723b2c594ffb5ec32ce3f6c7e68d0fcaecabaadda1d841a226025e64ec5b77990db2c0c3c5115d79af5f6339e626ba9f33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4a22927b3cf43cf048e534fcdef9f822751a42fddfa1d7afc733030998bfe7a97952974e6d9702e718a1e765b429465a2b9923df53ae5ed91de0ff9244ed3807938b80e3406b8a3f857e4235dbb86bc18d8901e70906906884334c5392290acadd7fdf566a70a93af2b61c892bfeb243b2bd2b100eabbcff311542a0c55813d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36daa0885b63c1c24fb26a5ee61ed39e469a3d91aec8e6374f06665a1a632f3d1183fc302e3f2283e73222db35c91a8fff0c5dbe84aa8034ed43e153b420180e89d0c4e073ae0ddd82015ff835caa540bd9cb049350f1c05596882edb26daf8355b7d87046d07ef1cb62d3fe977428afa759f5c598bec30f9d69af5cf2cb69a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9bbe2b388cbcc6d7d25664ede0ebfb0cdba973ce1b105633aa19ace907b938f5e88018cdb3c3fb45cf16a518fc574081e4a0c0426388d335c86f4ac584abcce2014edf520b505fff5e3de6e363257b03ac6df50ddf5248d8caa1bb3825ae24f441747e3568e0cb3251a48fed66f8e8260587f63a5e091f01c013b5f6fa2cdf3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha596fe96de5555797d2feef68e6892edc94779d8c4907a1b99fa64c2b68c25b5760ede89082989bc51ccf3d5a19bb204695f1e593d545c6ffcbe7e966c0b257b8d52136eb504ee63acc395d2a93a30e6a4559967f77f860f90281596c6c15f13a88599628ddb6a6b39653c89ef71d0dbe8bc8b1b6be452c7220105f379c14cdc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h822fea780347d9daca4465f6950b62c1205a333a5cdc2509868df22b553d63bc1ea81d5e7d60ec29c0a5bc302dec7e677c4c3af6c6943240a662f302ac063ec41c8e0214dfeb43f932d95505e9fd95d31ed52fe069ab2fbbcf43ef26981d6b3b2d845cc26791e10e477e39fc7b239306733f72682aaeb5565b4be7d6e99478;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69f42105d4556be5f8fa7e901b068be58c4f46cf1c8c41f56662a3ebdf9dc0c614dbb9ec2d503703f504093b98ac1fc2b09457b3bd3a7cda9f46cce990d03b8470b25789e651071954aa9613d7b2f1b58b376f050fae8ef6d73bce1d997b04afb81b64cb84315e5d43715b938a4401911e268fef11ed6c40fad209c3c2c35c3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e668260357cbe0e5d5231bca789a6714003a6246589a5a065661b3b871b7f1da4ab568d5a1e991a275032d2e429f01dc79819e2425fbf8f4495d4aa265196d5a65a7f79f0d6cce3a3703892069586deddc269157f4bd2ed49795ad05f55093649804efd74139b33971fb3e70aa2e72d83b4b405a79e313c068e4108531f94db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f8bb59386c2ac2cf30b742d3a41705f847b21eebced6d6a6d2c0d0f3829900b38ba158cc99a01e53477047f403317de4242a374bc7b3b9b3d96ff30b6c35dedc99c3f6c983880c903dd8dc7625cdba9477ffe45de1eef368f26fbf501dac20a55e809a601b87b81aa7815f16c3c58f486a7dae69422fa680f8768380989be2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd065a9ad096475f6dd9f5fddcb5cad9767093fef75a22f939d3f252008ef79e29397015007dde0f22233b405b5f7facba1843ee1f806d323943c4e76179986d0e072220836f44bbaa8bd4cea13eb3c874f326d87690b0a14ac151142520b25532c92962a8990dd6e174627dc79c90662f6340c32af05627f2f265fd0c443525;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fb60b75903a0440b6fc2671a74f10ad33b071cc71e0d71279ba86992a381f8908130161f21d60ac8b36c07699f8a5e8941e465fe20227259a15a4099f78fc65c3640cfe1635511c2413465a54caf1c106c094a54118c4fbdbdbe67ec10a6d868a67d09dda6670d8a0fa10451a06fbd21fe2325b4fb331981b878bf0c2e85d2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8568bd0a5d3dfb502c82d445523e946e1b3460ac9ea083cfd3991465a0b28bc99adb519e47a8e805ec799968f0efaece85e862fe065502c066e088d75964bed0c2a63f3c915e6feaae6df481bcc01de90535944d9f788359a9c1f10c0323c518a7ee7283fab0aac8137623134a11fe09216ff588bd12540cb3438eb49aac41f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a49026229e9f3d1163daa42d93af6ee24a7079a3a11d871bec44e02c7ed627ccc2b6b18622d7e697020b70ce23656701ea1f1726e0169397c3453b80ed5f835a43a11ca5e7ede5d915aa657cbe3678ac2740e8aa53dd795e9c09447daf9fd998c0b9dcec67f9a03b0ccd9a0e9fb90aaa322a44dea0cdbeb5d5d227d8b81f5cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedcbadc3095a962216cf075bcb9f32930deeb3595895f1233c82772f722479e5e097c3b097e66b6d29084319fd223e6fe9a722771c9d9bae4f82775e48a6bbf280680ea18be44762979546dd8b2cd4852bd3832aeb19bf313b2f6f0648c6f8321e3b4babc26b14917824c7351b1a7231c92f196ff0829a1d33ac1ab38c18182a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e5d29d4b386e0c38448d4d8532e2446156dd01372d2afa22b9dff849a148e7fa61fb9ce4eb857efe6a53dddc0c97d32556264de989ecb8958c2a984ac6ac38a0882123238f53e78a725ba699bae1b7ba6036c8d39c65fe56b01c35c14862635c89aa44e9554dce113107c38af0b33719e4947e7a38d7118a68acf59ad5298eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a4256e7076afb82f9a1e709c35678b7c30188a458e9a15db892fe0ad2a41cd01da432d3fb0ca4782f4d07a53bfa249ad392b716fddb72fd36371684218788dd290670f37c349e1817208c90ae3eb2d70735357e7f458778530fa190ed4334e0a71a45d55db5dec55bdf8fb29c9d6bc44f12e5ee5096ef0c3b4119e916f6ad58;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd72045acded42b37009b33cf50a27a4a036d306a83c6d1a677ffc64b1000952ff10117496241b2fc6a3c7ef6a5f9c726a5e7e42e696ee222ffd3b088dbedb6d16584c613b2c5b1e955e01494bd4c846c409398777115f52eb3b642aa7bca8f68b2d7465a7bc8de473fcedf747514c1e77da7eac736b352749be335e2675c55e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h333bf5011b4d6bfb2a095eef8c74fd00134211aaca8576f5d64275c4246f1ced807c10d3a4ddd27e34cdf40e7f8263d8ebe08bb4fdfbd364b30a32e5e57974a64d9b342e5ef74a478421f2209ef16c502f70da1a110f1d170a09a39a19811ea459da428b9a780bab62b769b6289c96a20137ea0d4da9fe590e9ed6330b475b68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2894a64841ed15b5d6ef92582ba3f5b4eef6c3aa8784f69e6c19682a7510837ad526ab52a8cc69eb99d269a0313c1577f7d1c8d8c56ef413b05cfde55cec7b8f852b5f52e09d416444bfe749c9fd105c0a06f42d08805125d62be64f52733440323bff49a2a0128a42fc47245c5f8f0e26e80e01988808378c4156b1eb445c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4ef0198303dec42960b4551c797e199e16a8bd86ae0cd08d4b8c73b5f4309f22fa9619cff7f6659ab76360ba5486fcf5e9d014759135b3847ae419eb889850d45c252c92152d653742ca505b70ac7d79f45ba9d1592c99ae7467c677b9fed8b5ec8e03a9c98e1991b47e30c8a83baa17d7a8d0a19d6f44f93f87eabb1555334;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c10a5ab982e51a0e0413a79e85e44866f448433c5da396386bf824784217cef7718570d3d64f8134358a711c8b51145c2a6898822dd18f6e8f3ffac8b7443d1386904ab355de0a4fe74c92183b181cd3530f29420472a927948fe05443283aaca2dd2f6c37c1e4919486f98e32e18c16082aa35c69f26235217408eb05aa013;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc54a0270c478d1a650c36dead6225dc7ba2945ee7af8d08b01ea50368c47162a11720827994e4f87ece09647380c6836cce0e7e0b36cdea93e9a3cc1b377e81912f455f38af4a2faccfdb32bd332380a39fba9a3c8df0b3e5c3b0b99656885aee9178f87abd1d4e0d6dc18d91fa93a89cb5677bbef3ecf4ef8216f4ffa32bb20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h244c225c5c4efde33231a5a22b18b78c98c2475bef9b3261a5e7b3dd128ac6f58867997dd18e38eefa157d9b382f09edc3bb3b3ce137bcba9cea43bda5d4051582691d7125fec8bc09692bd7b72ef1ff1de769a5c208c2beeda17b89f58f8d43fea2f321860575a2841c08bb10fdfead26e31689c1d9c0efc950d4a7d3c1f25c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bf1c1b24761243036a6b39eeb76d16c2ade2e2b1e61ba47bc03fb9f3546da97a869e610ebd585e6c2a3f21b7990ca61bfd7f33381b9d5a8308b184a34746349be2d74260bd2221a4075a18d2ec43bd74fd7c1c6610ced673fe85762cc6914f61cc7d3f616b623bb88e4029aff47dfd3b11cceb9fbbc893683133cc0512b99fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd55dc80b3494479c0575e6ef2999dcd164918066019b5bf3656773ef72a1d5d2b973f23311fb1a8c0c81a60d8717571a8e8964f978bc8080512997a62236a8900ec54c12b8977c0e3ecfb8558dad0d45c54f7e63ee314ce92831c69b046b91c7475a9a1578d49f01f2c1f0c81a51a1723525a9f5d2a2368414e0e19b727fd14e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb189ab38ab51c8d406a3d57103778142478ff62d4eefb5bc54b4ed12a6a1bd318d363f9fa678e2dcdecb27762a83b72bcfb16f088d651101f261e4fef5a0cffbd5cb5b3ce37537e37cd8325377d7e57cc0e8ede6b96a0a7c5b4f90b718ac112a4680bc06ae463e832f052c796502e35d65f4de787d8bfb3b845b2784587b7b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd22ca2fdfe9270d9b031f384288ebee9d28cb1915428a12775efbcf6d41b7cb6686b002cbfccc34c7a449444896b1c5b7d7cea5698206057055fe0ed9cd7b6bf72cf87074ab77e8f0f7fa6e01433aaa44b809ee7d29561ba4de7050b02612709e8b66c7e36ae762d8419791d939809590c9d6a93346022bf01c9c50ee483048d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h455c9b322fea26be441de247864d47d97b9db225339682ff2b6b3be69c0fac71af66073956e5fb558239ca88465ca31f19207be9b2d2446e07c0f6d5c25edf7bb6261674d5d4d8bbcfb52a3bbf6939631a757c432bbaa69a57268a8cc16bbff1ea4d6890640e44361ece129131f8bfa6543f93c5277ab6f77422b89b632292e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heff83c912bffe11b960eb279ab316f7fe8f025949c7d1b779f01413c02178f4737eb6af099c5665fb8b7f31d41e77bb32702f31ab9993cb5453644f2cf31c479349dccfe105efa2803a2679a4beb27bf29dd18dbe24ffe88ee48c8f3014cc262b51eaaacf1c12da7b5267ed08a3eb0846112562025f095780440c827e8c7070b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc65b35b68ae389ea828dea33f558e1ff9735377d1e18fd87d3e539134087073d38792fa58867a852b0339d853ef73abe80a37a88461d6874de9c4f896c8ab67885f8b94e40990b26bb4943205998570ec24c34f089f6bb28eb607802e0570c47ab098fb9b2e46a7cc389eee2cd2aa2b992c1fec8839c4e83781dc78e4abdebe4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b8a5e45893a3844f5a3b7e532b549f45923d53d8ab4ac6b8740fce7fa624c340d950c38f7682e33e90e5319914bf52e357292f93db0da6e219e9b0bae24cbbc209ce4e0e03a053081bd9cba5e6d0577d328c7455d96ddab11fa61037c98cf8cf5b6074bd2c3d74233e32a43cccfae920e21c2d7583a3d309ac699aa43676254;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebd71cd8c3df270cf931f839fd6a3933c27d284e370eff0f529813e2a5cd01830cd16ba0e535a0a22a9a9399193afc8c4cd7c5ca23cdbbb00c003cedc2f5b16bc10cdd7dcc936ef1d96e28838bdb50a4671c036bbccce16df478569afc9604d369055e29b116bd77217b45bc435f737f4594d09df201dd9d6735a97d0f56ebe9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86c3cdcfb41e1eff657a0095fe21293493d2052f859c85c0f7645f2f7111173c22d5ac8f37fe1c0f6092162decf4dbaee890d4eeb76ef11e8135fea675f07eeac2ce90e413c7808aba1853e4d3f79d8983a72f222718e9785e31840ecd6f8fcb1ffe926e898d7830a1a94a70aeb33e6598ff8e367c361a048a4ff38b200b61e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8586bd61faf6114ec8f4e26fa929e65ad02895815532a0df739bd5b934988c8e59be1bf863ee594158ddb9523fd80035418f454237903fb8ffb870de983a7b7071bda490b6ae9daaf2542f174e798a10bcab9889e5875aa75148bd27db72ae1fe8fe193ef28937784024d9ebcea4bb6478b6c0bf534fdc8454b48f03d8a9b6b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc9c6141386ee7a26539b9fb6ae46bf92dba861c20e2b52270d2e2ce28db2dda179dd9a4873e6dd88c75b7e84260497dd7e2496427d78b98794878481814a99da2e64ba98179682c683b450d522ca406d79f79562a76f31bbcf090ac564fa8da67384b70d8056f29156d77ffae5a50d8df7f6a08a31a957f89c69b532b81bf7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb339b901ad10f6e70987122c35b4e3607e628618c5458d6e67b8cda2bd960e5c09995f9c3d1ce5530acad278b0d6b46af53be56e1dc87c3737c16f23979905d2fd95685bb89de350de4717398161b5810657d462fffa07688380460f61fc9681ed491009eab8343671f1cd86b5862b324a3ff55971ca30a8eeb20917a22590b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13b9300ffc53092cca127bb7177e6efb88b4e174c8619cc20dbc12750597ab61b619fc1c8314c816cf84d182b0566333d07130df04b0603abf441830db7bc35cc074e06c0a7f05b37532b2a2740e97196667e17e4d7fbb97260905301fa5e6d384d5ac67635497b0bf9c937f0402c223249151118855cea48a4dd13814f599c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee79450e94ef3c63001c189957cd224b495257d3812cc0844be7b46621b8f51348d352e84db1d8b6d77ca9a0a5e0bacf6a86e1b45b670e1b8bedd6b0fadbb3769c5831c0139882f3b1e387079b1cabaee7aadcb03a4c215fb8945d708ad6ef9a317dbc7b379e3385fdb164976b307805cfd5c386b58dad0fb53c702a7adf278f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15a0ecf3346b30e639065159d4cbc401b226cc1fa7fc3aa38e0defa286dbca2100566373ae7210c308f9bbbfdc5e329c024a4d73d19f8f7c4d7b4f863e26c7c6337df1ca24ce9062e2697a195565a5743d49b314e23aa7730e68f122ec9f9c1db17001907833cb07f8c585ae3f74a1769209b02bf8d701b064b7aa01a94957b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13fef74e50a8a09f7bf015b7dd063887e308465902551a46bf2cf77fd1de537af0375f8b1f91a80f412b2e889dd780f712fe8f1df3823f0ed20c55f1e4966a847edaad9ce24b4de44cddfd836a3fd89be89aa04a55b7e914d755124f687cfa2f698dee27ddf7f5eb38d21b53c268d9caf1021297d5470339becc44a71359b5d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3fc3a4e32544bdb0cb6c14cb66589e539e1d4313ae7ae5e407666d5afba7b0868cdf343beae062f0a60d9c2299ab19a1e2c14da68ff8fc6dd8ba3666760ee25432888f511efec89c0039d4657e7a4af97f13d695072fd8e41b759c4e34bf91372410259976915e5613716c24c7f6874bfffaf785b4f1c20b9e16a535f5efe3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa104e87313bf36a2a75ec9eae204b47e8b1cd0160479558a3592beb8671a3b826b4785fbc7367d3e4daf9ec6cc2fc52b7cf4541983969a97c2a81cf0be7a6b2b6482796d2bbf0973a2c70affeb3a3a8c3e7a807b1d94bda76a8ec51c8310b9b3fe7b1d3006c17702db785dd7e2197b3e39cceea26b3454ef5453343938d50ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h620b372221e8172a07eb3caf52526bd1ad0843ba893dddc3e86998b1a633110bf45c5389100000da7e06565a441d8b979690d0605c8af494e3e17d81ed51cbf7fb2ea2f0a94725916451c6b7eacbcf6569d4bca90e33dbf3d687b254d3c78eeb88072b7cf80ad751f251e7bd0e07bf10a66aac1e18cd35c8368204b602ae6994;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7528a39fd3514be3e850111e9f5682aede260b4ae68a4b644063d0888971e24b5a2dd4590e47ca10ae226f212331c172a2e266103cc4b28ac034250d99a397ff652e5f8b7f765095edbc61667bf938a5cad6cb773376d39bd9b89e6325d24677f1e503cdf92d1ff26aa6f878b02216a8f490a1abc1cbb4811aff4fecb472fc7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d735d76e8e24b969685ad9330a60e34d3d85ab4897e08b3e0b2a72ebee061e952417800f1e8f073355771a4fd7147bba98b60e8b8af5fbe40e1dd45f81d4a84f7e34745fd50c0dbf3eb630e5d4f2df31330b852400e508a344894edba5ac9865c9f346293518ddb9ea7653d25bc34930b07a965f587b5726d5e99edf399fbf5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84f1e8df37636092b8546119c68fffa3589bf47a952d76b0737cd2a9e1b1f5bd7ec90b64e7d7771c9d88c7f405e6b3a1e94982d6da5a2f14d34b1ea8e2119c54f3ded95516eb5df94bb8cf40a685f0c7ba5a4e1dd2594fc735f8676449320158a0b4588b2a8534042bb86e4d5ff6e42863a763ed39722e160cd7edb9ab80404c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85848cf69559bb8cd94b5921faaf347c02f6df74556cb802e6048ae9dd7c8d6a6f00d7d5dee5760c5b9105a7d11c0fc813be2d15e1135f41c3a3d3631f0bcaeef70fcd1f789d3348ea82f63218284511d80bac4b37943341af8ef51a21bf3c28e122b9febf9c19e1e7844ef3362bc0bf0c09c99d425c8d40b6469cb626cc9ae9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7311773335bd45ef4a595ce435333d448966e6ac13ed5a7085f0fcc9e26e6efd0cea2630aacb5db9ba4231f4da724b884089da5fccb31dd4749ea4da1c789891a21f9982b4f7bacc70030a21a0f062e5e635a3bf85735bbba2e093a650c1d0b28b469c69866fe640ea46a60d89d97bc9e54dc9270c28571567ec673606fa42ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8f609c7a8ea567c0ce8475ed9c95ed98f4e6ed61d44084665b6cd8334cb2741f85c1420fd9d35c979e83bab218114f2f5e7cb71bb455ad6e4ed6eb64531d7ce74702160ca97e571e82a30661b7d0df2dece13b5f1174d683fa82778795849334aed8c29af8fca828268437a2ca14e890a998753d640b03ee61d9d2ee076de4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1bdc7a74f713f9ab2d0daee8009db6ee2132624c67be49f194c5ec0af602789a48be9601449b3d966234f7b9f7568441e670006ea2875a7cb0d89ff7cc5bae2314af75b7a76e7818e602312b70baf3e2f1362a03d44382230cbe5d8671e27efc3252e0e41dc542ddaf845a7bd1fc813689d2ebe62c2caa384cb5323765a5c83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6dd5689fe1e1ce8d6fea1ce4e7972d6334e6ff1aed8e0452dfe0d03bd241639ead229d4e266d60cfb66f46c4f2ea69cf0279be3fcebc9ff8838894dc2b4578d35134135e6dc97f7a9d2d06316861689e9e71ff849bc8a5571dd0e9dd0777f4ebe788a0c07c4f9cd908b717f6dc4ac6917b47f47e5cdae125ee11ffd1986b56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd895172f7bb789b089b727f782ef4e593bb699b6ee51ebb8412f3f7bbd5fa2a61b62d4c9eec7a0c693728d383aa904911e5340f8967283fe1b3dcac2ce2869f23a8026f8d05631b15e09d3a664353814352d7ad8d9d707d57028dbb707b5c92925dc7fd5c7cf94b12c7aa2cca8074a0a82a00fd76083bb895dd2c600d1f8da84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a2a5e378389aff9273683d372e6b3b5dbd8f38592fa4a553d5202f3febce82356e7046e5c88c326c4f1017455fb5dca9fe02b5584fdde82b7ee509eb3837c83a79a9f49df80fd65d2973c83df90862c5655be9bbd0457780179ea46513d0d30097572961d900f3bdd62a85f7442fc3cafb4d5c77b188112881abf1ceb1f880c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2611527919d513e22af059b5371690e5adc25c47370bf9b7f74546557f6060b45591bbc75c936128e3fdbc571d9d740ab089dc8d89c78763ff897b0bf2f19dbc4a2015e808cd4973f9de3705ebd034b9476f417d949b2a673dbdae299f4df15c878a296c0f02d50f75f1865740000f1ba354f5da35e1a9c289853b7bd848ded;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66e8d8a2badbb3d6d08ccbf90a591fcde1b7a556c0dc414fb0864f3d8d8d7fc8464662e4ccbb163fb6e678329c0ecd13aa7b4764429e34e4ab6c03bdbcce48641d7b683920321766605e5da717a36cb1baaf1ca26c765711999ee514f19b7d058967b006e96a175b628aee9203a984a40270b2a4b031ca1531d69f368cfebad7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a265caafd3f3e4b3697686dac7ae97dd0e49178efd8db8c3f7694f634f0d150575364b5e825350f0d7a7c320bebd87c793928a1a506a0fc8c1afc82a131a3a7f861bba7d049e1819674f8bec6375caa2c84f9e0015845b8b1cac2ad1346a6128a65ad7a1fd7d9a5c14a91050906589e58b9e1fe04db95ec25b0d5621bfe6949;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0f6ed3649a4ec190c43a75e436d71a40073e3e1ebf86103d75326d44c5e2b27a43d25d81267507be85e701b1be0b01da5f660dd911937f5b338f8ac1eab45d29529fa3daa03635a73f935b57e86536ec737199cd9992da5cd129d1a9972a2bc34c9215c5ab0a40a171d65a6b665aa5b32ab6430127f0370bdc175cb58b28007;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9379fda6acdb0a893198f9f155d681a8e249c997ebb07983a58eac3f5bdcf7b08b7d1788af51a59c933c541c4cf89dacea06d7759d3bcb1df514f49d19dc65bec57a15c3c8849ba76fc37db454661b01b0ca5f387442dc6cc4dbd09671be01939fcaa7649d45625a947064cd3cafb183ffb847c2750a2376f5571c362925bcf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a5007697909b9ed58ebc8e9914d1cfcbfcdb46729d5965c120fdb4bd18503196e355a414bc47fe655317020b296b2cd22bfe0790133f0de188082c99b12ea1e2872d81e01c097364956e735b130ac18178d2884f4987e02f711f871126334966b8ced197f3741f71aef098915f25eb85b4ccb3e0bd81674bfda484cadf7fbba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1575b6f2a1564caecb91919c8977198c22af025805648de84127c8b11c9f9666e63516e686169343c9202757079734d124f6a354f35efa43bf3d3d9f2b5b3f67ec5782d0fb8889247b1c56f9d42d413b60cf670483215bca730fbe11e66b88b1ebe08b5a78b15cb8515f28ed5398b8c2cd2cb53d7267f292e91fc4749f36208;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85d3e401a6a97ae13d44d6e66e198c6184423aa0bb507dc43cda25f463f0debf370b1f199c70ac31de030b1a1ea65174f093bf556a2452290ab39c41c3a72d0397aa367dd6572858ec38e6eff9973a01e4053f946a3c386c6eff27d53209f6edbb59853d9a83a523e5bb67977261b22bc8ebd6975383ac6d8907480c04d96919;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25f2761c959593c7a5456e1743492eb30749bd6aa83d846c5b05f03c161824a557b0e841e7617b3ee3035dfdaa3f490583bbd046841b76c5725b96750279831d8b58511d7d35347c5973fb781daaf3078be0bbfca602567765302f2a14d44b3100695535d7d7cade29219b4ef98023081fcca1b7770e5fa4f139d6b0c69cf199;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6515691e77c73fd75b7c8166b54d77ea8061ae9b9fe76623e8f53231c78807aea3907dbbc80bc1c8007446557f8d461aacd02e58ca46198cab323a504be1263db55a07b26f05c31a87f92cc7be74ed43f64b30c9edc2a95b3bab1daf4b17621bb79dc7a71f1967fd3921dafddff38e16ce0e1572768c8ad5533c8d71d0b7759;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ea724eb085540ba182ae5a296fc8923939d4d8b2a487f78e5ff04992ade562a1a18a3508d9f6bcff019fd1cd1cfbd1cbe2a0dc0678fa77f90e81087ebeafdb22aab7f09fb7dd1de78649e9b66ae09f85e5175b3b86c27746abfe8ee93bab196e0501eab6e8be36824f7e85373ae874d3f9a68b8bbf04563514639c3ae881291;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7dc195527d9348c5e4a0e6bbfbf009f3206450cab6daa2bd9f2b93ddac2451691899f88ca50d274ef72abdc736d91d12883e5bb336fdf3625ba5e6a67e4e67f56574f76870f33d83827be247558864f84f54cfefc263c377c64cb70b36fd006e98ef0da02ab4af82e00fc2a29b54b1e359e758735517e9df2a82c1b3d486ddb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3eb7b3270f0553f14f135ce82c35fd9805e7cea553d341d3c122f620c866c7501a18e9493bd17ebd7d77f38e057c45764132018242631f7099ca73bae9b2f68118e68710a5fe8301bc736d99e46f6e44056e6b41fcd18975426fe198e95fecf262de3b9600b20a60847d2859994d7a0ff6a09d7eb3a773a77eb5c831a27fd785;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fe79e98721dd7ffb147bbc70778a98f782b64bbcc834400e43969e5999441f59a0bb8daa2323f1bcfdb2517405346011c993a7b4da742c5072d024084965b25e84e480c5d889c76d5d5b154d63cfe7028b223b11dda57078cb41d1104722a229ab2d688dfc71371ad0a7f8ba228f2666f11d1da108a00213979ba330a63f216;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9490a5bef76e6f2bf7a03e00be1ed976725482e9e4c2358e443ef6f893b32e2302ac9f629f3bebe1a3a429357d08a4691f731e54683785176bcc2169a74900b85e0db4ac357840c013be608bb5eb6e3d39600c849d289a13d108d8df1be1ca4d847183a7c7b2a56aea7b36160b588e4b020720328f96157a6adea9a22a83ca72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20b96ccf19d08a7b3dbe80c037c1a6f4fa5744696b288140829978a9dc491594c2427abd26bedc6b93e3ff8cccc24ef6c2b0e605ab9124bf950b9bfe602381f3fec905ddc00ecf621fdf004e1b0bc5690d31091d5a10f2ac3c713db2ff6c670456ecf2cd39c5e2f63ed991f5c02d67db6b1a698b409f18e2b05df9ab7fde070b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habd9a2385698e14e8d12deab4c2583cd0d1745a5355614abf3f084e92c8536fea7a5aea5ef60effa04f3c9173f29806656e8e7f3718e8cb88addfd38d6807c9e39330e315a05014e1625eb83971f2e5f0151729ae2f0f8a21752b9cb3cd46155625768ced344c16d8f2c342fd8a2b6932f48b32f13c2adc31ba3974542059bce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6353ba446ead00028f5290203a5ae6d478697f902d6f7f011ebf40bdb03c03b2942e0f40ad1f136853f42e0d5870a6d35285be4ed4c135d9fd5321befc4a7227f4d88cc33372559f2d5d518008d02b6771f2c55d43a2cca70ffdbc172ddd40bd47d6fb4df875965fcfb17ffa1983354cb06bccef73d42b7b6e09a9925576ef64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haaa7014619ce1657f2788c3f56235202a65751780a9a9b10136cf1d5bb7cdff4930d6151f2b7d457039fa3d3e66862c475bc267f73e147fb984bd4eb8bb34d567afe1302e9b41bb4cd6e14b384ef873e2ac1f7722a7fcfb720b1f5e48db5515e549cd6a3ec086d74e0e10177ac36263ba953e6a4d0790415c6a8b31b30afc308;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d4213dae555688f4f6e43b924f2bff0f67095523727d9deb53e4735bee035d7d298c34d311b245d5a534b2df4608c5d52e5c6c2f885d7d1927357a85aedbbb0b4287f181a875fcfa9094343b565b75edb424331e61cb9ee7236926819a24c4e70a7fa8573121b0c292673cbac3cfcb3d47f01e01aed246982a19505f09e5f5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h546f41542dc7bf517480d717409f5ebf8ef5d8a6095b8275d1439ae4be8c1694e157f6382c0b2849e19990c1e5d14813c62be60a20222453241c68becf2c7023e8da842e18a104233246b152f80a518c43f16698c48e11e43846ea51ec49638b281e865cfe6ed20298cc9228b40bb12aaf0a4181004c6d95ba2dd6bdb453a15d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4af32b5a39151e36a6b22b1950d6e42aeb3d3585058628202b4d8a0085ae14825f2e5366fef7700242be10b46becc768f919e5581e519a3679c9654164bca6d50cd896b353b377a13ddcc83d2b1c6553468b53e0845411780849e14ebd520bc921c4becc1e8a25bc698e23e4031540023a06ac6698e6e20bc84557aac4bf2398;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6970aa4546d9c8fee9ca3651ad755d0c375bbe54ef47eb32ffa8c5c7324f4821ade7afd00f5ac2bfb21f6dfcce981d8a9476c5cb91645e0f238c41c396c4b74bf48ea5246d0905bb72e9a96e56fc4c52cee8c35757c56029b599c841ae94ce102c96c234a1287b386558cd3b3a3144176a39bdc00c03cc56899f44c106609a3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd74b64b91355f8fb0b506ad05f3fc8d363d9d95dcd911f60106498e6580406ca74328d3d5163823a9ba57ea9fc300e6d9556209cf27698d25723ec7c1fe3de830e38d05094d5368b69bdab0c3a3f45694f85b3e2b3843706d0633dd833717f7bbe2bc2b8fde6172ea856b8d9fddb63ecb77d00a54095db08a73b2c322338fb21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7b9011b169d2dcfd0d27a08954942a22b6caf0c0e6d75863703974b435140bd8cda68e2d7f149a73a9f42ba2f0462a5dbc15de8df2b5cf13e1f3a69eb0dcda10623b04c3d9b46c2c2583badf802b6e2df033c69e76543569873bfc00e07908ab1f1bc39de585b4ece5c85a3a2699b2d21d0387a187a8f67581b640123029dd8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff6e194ec1d1ea809166fa5e33b669444a238e7c506bfc976106325ba1fc24f8ea5e8b545d12e85af2c4209fa0b68322a81c4fc2bf8445a9e5c36d9878daf735fbadfbc6d04a30a242d9ecda0f3f14b42825c12018f91570b1dee929a87be1d42595eece9824ffc2dd60d40312a1b8ca6e76beeb7433219d320aa5e70970a19b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2f250d5e443ca812b732ba333465e96d13ce6587400e8fad1602646ebec5f60a5014ce1f7d08b56b138cedbd373cc26ee89a71e0a234340e5dc986006bc97ccd103d85a2b6122b2aec86588132382f05808ccf567d5f6c9d22aa7ef2ca235bdf0259be6add9a36e1e98bf312d208cf1e9e087ada111e15097171953333b3299;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h234624a5e27c80d4c5b9fdbc12b28559769109ffc44e8e468c179f4796dd6e6cd8d8ddd885a6f342ed5b0dde9ee369b77321c5ba1aa6cd2a009355a5808be79075953f197d2828dcca22a9610a8d4997edb0e29feef0a83f2aaf235c863348a20cc2807e6ff7d1b435b23a36927f98a4841e3daf4dff6879886c33941bfcf9d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc31a674ca5b086507a2ce91219e2cce551fb9d952bc34bb8663f6bbd970a2d21ac3d20d96dcdc5a91a00ed79f7213597f5d923d38f8dc6d714d62f423184ef7662b37f19350e76d1c2c0f4b516f3664ae9bac9fa3ba5962914fc3119ad5220cdd3d1be1be3fc53bd4df135c66759423e24eda969e4d010e9b1d6a55f5297630;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56016744f5d62ab74089aaee8507438cf26443b25af0aabb4a9eac30c0c25ea5bd859b880c3a4bfc44a6f64167a51c13f8029b2520ae2cf74ec76539622f00a4f844345739fba78916fdb2d769ca32350b8d9483e7db12f3bdfedb06e0f08017b843926e578465a990cd46fbed2a0d4f83720c3343f3c7725acc37e8fb6c337a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e9e0fc3bfdd71e23dcff4cb0f37dd35e8ef6e68490a8063ac8f064613c00b787177cc26d659a48cb71d3e399f9300cbce277d3efd5c63ea2e24189894d3f7c79ee5c643dece05630ae1a7bfc1bc857149f920af09ae3faea0c98064ee82ef5225956233b5eee331cdacd1e90339fc1c505d30af6b518643ac231bd525db3f6c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd3542668f3a09490c6c0c3023567c6381fcc43244128a0d228986d8e89787cd8aa4e4459e6609baf48bb57c686d442a006801173d9ccb95cdeffd2099228f26646f1e8b8d80957d12b294f99f21495729269aaba413bfd0aed251a5c4924e5b2262ac31d3a92833e52420e14a903df4381dd11c501aad23e32d2a947677af5e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75ebeecaf5aea8c6e8e875f818a06cc007a671f6ec5c54bbd9664cbb1141f8283c73b754a09d8ee080891ec2cbe65778e1ff8b632ccdc90ffd202c99baa4e40dc4e322a75aaeabca61933609399959db9bb40c426d4c926eee865c12e14b11aa4afceffaafe0507f2a266a2bfbd0086d659756bfbcb3b90da238aae19e9c396a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfee16db924c6c60d803b8adbf69f903dedf8ce80c10d7efcec77abcf798fb356fc00924993c306b9fd4a99092c6af5fb38d03f7ed91b21100c66673fb8ab932b7bf44a5431f5f1fcddae77dd64d9a228f3534a39429574807f1014b88e117732ec39b5b38b1ab54463cf802d7f9cdbc03e824abcd61192e9d051d58f6ec46ce6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cb85410eee88eb16753e4b10f9cbad7baec4cc32df776f1e638af2bb0750b0a4cc87034904c2c95ede9969ab0cf6dbd82264bf2a5ae7c25d45b11387e1d8d5c79686dc8eb6a18de87e807bde9adf187ee45c0d7ed8347a900d8ef763e7f0408c1a141e12174f8bb7515070add3ca4d80ef07538374685183bab37cc52f27cdd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4dcf862b9d0886ef6040222aeae298e06e91a0c44a6aeeb09c367c1d2bf828edbc8a383da497c7627b8fcf577c54b42cf90a15432429767f120f9d120c2bf4a3afde356795f1aa655be60c2c8fa4a885fc3539e8459c17b37c890b98af01d1c475dc4b286148d312787a9adb7480d5aa5fbac2d2ffe681ca6ced1be591247743;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92cb1aa0611795cd8138e7319614f33a22bc6d305bcc5e38af018e24b63c30828e21e3e85d938019ad0f895cb427e3615348aa5e3e579d2aaab4bfe410898d44873e7c3d64a20f50c8536c76970501983bf322d5a1befa8a8db53165a9bac6ac9a0988ef5da9fe6219ed161141e956c62ef08c317d2e83842635f62d20d2d99a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c3d7c618a915f714c405352397acfaea516190ae4b53d3dab2dc4991c2f19039431924b4221114ac19e43daab7e922c9aa4a73569f32d7f9062385211dc06a92ebe75bafc6ace40f41cb7cb0a66fca1b0361ed26779b95fb87f6aea7f021705c200ec6c910a98332cfaee8650d48d0aad9b6c7d07b96456b8d7abf241ab145d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h813c4b30a7c59c9f9623077908da16b4bbcd77c83a1578156fa963d6074bb1f2657b8704eb0a8bde16018ebacb976efd9eb853d9bf6f990ec25f2d8899478b3e00a154120a0de59d6e9f950120bdef3ec13be8d98b8b74617aaa9ee1ed17bd88144a968f6d32a32166370e83c94c4ebb2926419a4fdc845818dad1c551c2f7c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf99c9d06d62a21d9e813cdf10e227479d3914dd1c0298e12261726482a4841e61e2789aad6886a6762474e4e8c29761911e1c4b50fe0348515345c9de98c30fa956094ba4a757605350d6e356f72274bc6562dfe079c4cc42c13f9e41840772e4f68e67caddf0abf778420382631244a173b3c890b9a959c840b0ed68205a56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b1e1c4fbb0fb50e3946916f908b640193a926075c3bb388f61c8ed591b26f46702735491f65af6136140c52e8f162396f5f8e4da387cb60937e3c96809b55d87e2070f70b553099ef5eb28e1913b4041d7631ee843748ca539a1e94f2fa6556ac697a0e6a462133366a12e63167cbcace6da4c58af80fb42da7c805d716c2d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf75e93e4ff6b3733b215627643402bc9017d63663404fbe8756f3642d42e43928c5bc4955358f6976a1e30a149ea3d7d04eb036ed060bb9cb9e4a7d2411ef51b3b6f5ecc04226190177f0bd2a64d0522275740841f9098a70f9a0b790eacd758751de25ed357c7bbd7e6618d7f27529714cf68e1a473e83003a391e6057aa8e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d81334587f5897116c791ee437f0121b4a9c618529282eab1de36476fbd2e7725afa105956d487c03e9b3e38c71447b9ce7ab6e6b4b3a91c9cac842d0604a01a8fa28d0befebc8c27e3e639767a2659f448a324f40bb6c14545fddb3c89d59ddc4bd0d39c7191ae4ad3283e579e79a2c5db2064c86edd019b40db68a45753a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c1d2e12e22fc7a8bffa10516916a395e6f6c3f109770c1cb0b4bc46ae38ba3523610e384c7c9aa69b9ab2f86a303452906eab09a0108fa8a01ee75606ac03c4f3605444bff53119d5ed4218196a17dbed376f6416bcee67909ab2495cd9174c385c2e636157f71e2834e5ee86f2f8535fc9a5c64872b2c5305e500e3594bb5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6bbb18cc246581c1d9376f5f238be253202df97a5d77862ba0eaff0a1286ede461a6a91ceca063991a088854e776ccc6ae1a484af0a0c63da70ad5c517e9924897c85a452cbaa66b94c7921c2228e15a82b14651a5553364de6bc5fafb855254f8ef3a6611de378af33e8a851abbdb19ba9aea12a5475502fe687ea61d4237f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96d59b26ae40dbdad75dd20bfdacef01cbac40f72961e6f42dfb7c96655a1789fd24bb865003e47d9c8b28c4fa60b5a9a4a5a9a6eaa404f8f7ff98082aa301980e48fd249f6f76a84ae541bad2c51846569314962a0c769c5aea7057aa1c2f6bfacb710e15a623500b2aa879fa3dd1591fb6796fc26ab4e214432ae7ab09f50d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd626aa79b37a4db48262aa778c1c3eec4a2e35f808bf20585d104cd4c1d1b92042cc74f5ed62b2678e88f452425eddd45261d5ff0f2940ef45475c9a48455a26d55caa6f162854258a9145d574f146a0e83a9d44e6c2e7a884d2f7ab6a46ae2fb5d0135a5b4cc78ba282adc8355e8b36eb91daaa989d2b41d3414c022b1fd903;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae47699b2d01487b92bc24c5671e5e04747a986757fd2ad2ed986b8ee314315362024d2ac85a3760df8e34afd51a6c7df9154a70816b5172c9b33421647e2c78c9a3e1794968e2e915ad8d4d48faf3e8b7967e4781a5d69b4b920f545fa9dd1bf0792c09943bcceb88a74e9e935978c89b09b948181c844b19e4cdf921a03879;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf9c08b01dda11749fe331b2b5f862bc9e459280dede874bbf82cc287c49ce4ab9835628474c858a4a585a5fcba5056c88824bb17414cbebf8ba351d2f4018b65394d7461d7731a59303661ec1b82fb8824a8b138f218f0d38445e9fe3ff6c5299c9875f0e24cd7fd27d6ca0dd2233903cd98b198191b67c27c87d733f8182b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12aa5a601324b60ed6bf9a974afda9e3f204dd91580a9f5874d87cf662dbac73e4f4c4f7c2ae6ecf1e6077af7caf522535874ab5b879a55f3e91d4075bc9a11c5dccd436db0b57e58d6bfcbae475de99e5a6c14e19dd0020c9231b9f9d8be178c57a2b1ec4a67be2c5e1afe297a32b51e18d0fdafa6fcca5aebab99690f1872e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h407bf633a52a26d50f003d5e9de3e528083f09294a6540b5ef38038ca85d1247e34e486a755964a0c04231a5e7d5d4948299597e854dad94fe0238d0b51fbe2f9b7ae828903a0af008f122994ef44aa077ff61197759abaebcd8c72f26346a791565c2cb321568cd6fe9a7be7173749a3bcdaf5eef418d626c9a1c869925fae6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1411d1af8b25bf77e5c2ab92f287dd440bcb238f2861ffb11c7dccb2b8da2df10eaad9dd1d45aa2ce143a6721bc4ddc94943d000f8c71ae3e65b0f847a9c94ff3b5dcc930695a4124ef592c325737bdeabbbb216fb51c9a6bd36282f17c65ae8a1bfd84c0fac9562f90a0a477b21a5c91077caa332d65c5a97c5e1a006741fd1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64a79e0a3e6187620e1f124ba2f2e7beaff611a36d76aecd5e8b2f9dd9395a91929847c8a1ae4229b288393d059365b0b2685cfbf4177aac98448fc9de6a340a2005aeb9cbfb3f2191e3a3cc007f8c68016d9ef4f22dd6d5362ea135d395c6e41c6482d1fd8ca0a4ca8a1d89d147f6e108a5422265b3b0c6dbb3f8140396fd98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b458e540aba483d99a0b78ef099433bdd0c9bba6b698a1b59185b78e3d90020ba4a954d8cc64e8215be03a07bf40252e1ba12f73a646cf5768c9fa8063247f2448c886a103f305f3622f734163d798c6a6331ba83075dde0b43d6bdd75c4bfd6913617ad00b93caa87aa03007902d2fd3c5d990e393baa499ec3dc4fd085eb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he34d5b880b844fdcc456c4981bf81e7faf5b13e420ae3cd0fd0bf4ffe5206fdb5d475709e69224cc1724197f0d16803d6755da19f37372bc5d6ac7d23fdddb8dfb655141e58ad3bbdb359210d0597d2791e25cf7fe0b727c6cc269de779cb3056d5e406916046604c3e98cd38f44e03c4d35df6b589668c48df5c1d848e490f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec4c6186d19cad9600e553deecba675a435f2d738fe5918ad0ab8c5abd459db473fc2bd7fa4166a38e6dd82d561f3f78859d0279b46244d937fcf239d54c24a34482a97ff4099aad1ca75a0b3f57806cff867685f249c6158acbcb56a7f1fb5a7c7aafe1b91083f37e8b08c43594c02ee030e0098acdacee8f2d135fe82ad0a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h691bc846db926b6bf5f068c6c2a2a10e20a81e059994ea3d323cd95804e0ac20f9f7a6c31a76b05d778783e890a4ac309541ae8e5ca45d074464b6a4e8c63d46ffd4b36219923405bc029f948261b0202420fe5ada34b78bf43801d06b2ff6d5d480ce850d2b8176dcbe05cc761604e84ad9ddd240df299f51e748ccc4c02e1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdeb919690b9a30caaab7416d7d7bf8c5e1f82c55813cc79e2ce4dd2f7858041cc41b8d56d0a66dac218b2274180bbad9f3228a327ea343ff52cb880c397173d259e26d558d0a3085d4c173376986b02f1e23a7cab598b1636ddb3b3b3dd4d4f0343d94d38c0e140eeec04ce89f662cef2db8261b8085ded014e48518b958532e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef4381bc633e388c27868501debfcb540e21141fd6d7609c0148ed6ac3875b41aeda2d780adc15d37e78111ea6dd1e6f7731ca88c2eda7a1d26278889755e6f0fa45bf4ee2c9530f4eb5a40afe3388859187137863f553f4ef1f87c0c4e97d60515ef8c0c7026e8ebab53e9b29c988e1833fd63a87153abbf5d2ef8f44bf794d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc53bc7eaa0a49bd54ef14bf2bc98446556d01d637995e9e642c6eb922d6af5ecf921a6559ff68cfc73a9d1dd387cbf932951e4a38c3f53e6779ed1a1fa189ee44c146de4e62afbb0e0ac1d2381bd60fc42d3427447c3c05348a3bab911ac3eacaad2befee1d56705c5fa06e061221e83bfb0ccbc3b5eb96cdc2ddef6d23e0b05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafcc06733543b7ccd8f15b8afb849d87084429f05b7c66e3057a67e2a85d2a0af2a5a76f22ebd372e2a5d1594eb1f668a01938239f1d1dbcd0b2836073815b0e9c592d9d82097f422eac87f1221885fa780a86c974eece5560b82fd01395de738e985a7299ae1e07c90de6f0ced62026c871f99a2d02a1ba48cf5c00ec318bde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h463f771475bcb48d3541abee06526ec9c950b5fe056a8961f7b3fbd548ba64e874077b6e9c45b0b03f961517a3440bbf56d503d991aedcadffd2c491ee3a198183bd2927c2461f64c4905fb3e1d2798a536a39630ba7a7edd7fa855e2495b3a3854232d5c78905239614df184ece0f6565fef8c89f38e7e886bdddec8c884be9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81e7e22b2b1d9ca316f5ac99f2c765ad1e321dc6b2d0a25753fec70856e900a126e923487b9b9b1c7ddb79f76b4726d60c16ca8757323f176f0739600548d81382905191d5cf42ef33a4ee80e75a48b97c2237929cbc5eda607811d48805bd9d634480d0447f5f7da771d819f256b9b719ff84b2d003d7efbf2a39ce75d26aca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3887ac80f7735d33a196d944a571bc9b9fffa350881c1e7596600238b2060f66f06e46f077549011dd6a8718284b41fdb2cb070a12782f523d38b3cfd8610b5cb2664438400d68c87a7b87c613c2e5d5fa5269aa2720b2d9833498ce4df275adfb90d343316542c3f725b37f44d27097f8fb05fbca8fd5543000475bb4ac2f54;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h781c01ab9c6e344230adbbb043f1d9aea202a71b841132a8fcd5dfd6694d811420c278042809255c41f0e96eb4ec4971f5b46f9412e6f87883efd54de820792a4cbd6065d63834960f7a336c238454957e1055c7f480e6ec3893c8b063febd5df50e3fd307dca5f0ff99a4a9f262a0d8bc8edd7dc6b9c9712babf1c69c5e4e37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4651f70de4808fd039c80034559aa4be52b86dfae36063e05fb8ac2fcf72f28e633619bebb1a4e52a9772deb92b598a5cefbbb7dcec17191051f01f001329dbc5219360083fd6a0c30b2e52a1ca9bb3fc5509a7917e7d04c1a1efc8e2b6305eb4c919180f6461ec1144ed1233a18fc56a9211c776b8ebf80e848fb10ca2477c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe381b2eb8881903fdb93cb498fd1a0362ed1edfe7cd5a3fdface0bfa6d1475ca947fe103d3b4379bd64c6321d88cfa93a7516887b6b1cdbff42ab581e1dd46c89b7514dfebf4f3081a820c329c35be32f683a89de9cb8a5edbf4b1589643dbba2ea2aa5f2d355cc1b04f0c8262f24ba9334cf47e3badde2bd6e5b055c6982f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb878bf907dfbda4fb8f796294adead773d980c2948e4ff111e8f5596246602b27b0266c5055c7e440734641a957eaccd5db6719e80e076c8473de960bcbe5733a6ecdb1d3cb636a62618af524998b0bc371c96e72058639c104c4b373d6ad1f811cb758ee34c551dbd3a1b178ef31c664db8a5ca5196d9c412536ca54d8031c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87655d1788867d379f5c6ee2b1f0c5c40f355fd80b1444e9619b714ed1b68c56762cdf5c95b416451cd97679fbb3464feab3e04552e8caa2674dea787add21fbdd587035ea8e260f52b17c14f186bbbcf5697f187802aa6f78254165f8d7d74dd97a2c3a311d67ba4415e11c1f3d78a868a8da2d54d1866050b76af37734a06d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha906bc92718cd9c69634e7fcebe7852b0604cd37f3da753836ce68b40b3023d376b1f7c22d63fdde4fb1ab24e8fa9c7743c1f83e8fd511b8dfde479105514f6911f1f2acea845e7f0f940a056760223e62fed93ab799fb7fe691022d02fee9c4ad6e525b46e0b0f3a8008dc49ac9e2b90d161175cb6a73625d3072cf6f382fa7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h674634f6d91b4e55cc0b1c88e967a9b0c954790fd6090431e1b2e39ac6b4fb8b0ca10c6b78ff31ba0b8a7f64ee8486168a187e048918841234dd6b2a8daf99d17612b7cc662d479f2732b46e4e5ab9e5e36e9b5c1dc95ae60d4da94f0d7c4e8898dd30868f9b5392f54d63afee70953a2ae40d13fe29e5a8866b3a5b847f929e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2321d10475f72143af08bdeb3c73d2b989e9014ab233d5fe365673a33135a98fd483b08e5f02f03187b826b5718da94182490d715e598cbd573ebdd3d1dc384a508c5cd4c3df5a6f3fdd589d448b286d023424b3aceb4a37ef98a63b70c5752c219c1cee36f5ab102489a3733e34f4db069ec132c0515fb3736d6e2ae9d30f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5342eccfa9a459dd22e2d8cfcdc1efce9f564db7f794b3b74f95a631cd259a51df6dd963cee134dfe14059f7a79238525b5f462821537a00f4634df2c9df001a810251dc00ad5d241a43cbed5cf20e800a209cfa60c12e264bec815e32c09670a3b1c210da37b2a6bbb5c1efc7089b4070cecf25c3b518e48a551b0dc5dc1482;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3e1e596b1a51405a72f194e86a1938b6201cd2cf0a093279c7e19ed6087ba0d88e8867bb69fa957b87c97651481f5114c28fa66314ac47d5802ac6ddad3424a19d195a0937fd4e5bcde3a170127e8fd6b1741c7383eb5a24fff06911f5ef8f1b7b16d1dcc27864a7280050de52960b06fa4ef26fec29f10ea1fcc51265eafec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd65ea62ad6e17da6e8ff6f6bac2c8279d4234c30b6abc40b47fc33d1051b4b9e68218b121534841a1520cda602bed683579707a7189be802d294bdc56f8792fb24cb1a92f6d62e8aaad1c4fa90940cd16b350697725af38a6aa59c07d5f337f8f87362376d59fbbe2519779dc53418b69d790b18ea38838a81c63c2c1b9da65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5414457ecaede7002aa6d05e36ee9244c59ffc99a14088a762ddce51dcaf07e475de00708ba464111b0c8cd11c8310152ca69c3aef14d71b78f75509a924ba345497bd701be80d2b61decf9a648795edf54949e190ecf34c0cd115fd49cc2ec2c5f6971b3f414520a142b42960adf8d827d6e12a8cef77154ef780e6d2557f0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h266124e411c325b92ef9a29c56e778144211db4e58efcb8be9934ef12512fe1b2ff60abd06762c09afd5604839456fefda0ed409f5c33d03941e9b1d23be5ef34bc8f8ba0bb0164bb431a9063e9167d7d92e529ea3abd8c20f82d7ef7906c358a682b47de4fc24df07066308356ce12f5cfc0e7de6c00c4b510bd2309eec7a15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6ca421f33afa6f2c667c2b058bc105996b4662c16e5585afba6975dd7cbbaeb88c220497fe97456378efd4a1e53e5667ff1757c1cf831561a94d913c9d5f48aba1ab4f9b9707c12e57c56a5133e51b9c06b78ea6b26d68187f051b89324dc8917a48874bb81a7cb16b848f6626f16130143174352aa6c35e25c8f7875542a3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd610dcc747a36dd161de88dcc1227c57c225561ac6227d9cf89d0dd0ec987d66339da59f3d3d80f42909afc719776ad1f58fa41b67487e4408fcfdf69f3a073d7a7bde96b687388272072667c83566a9025a8d569aecb4783642309b351829e52e49d0f08ed5f4ff12b504b82ff3b1493bd51f0f682ad44feced6edb58d8760a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f6a61c00c794a3d145569ef79bdba4eedafb4abbfaea8c57419b11018c87984f59c6381233b8dd7eebe2c80c3aae21bfea3ef429445f075575965cb9a35b7648f7ceace5a08b5a12b6bd4eb56b6aff5db3dfe6af18beb0e19a88b168769dfc0e56406b33b5903c5b0691a8b868b7638808774e28909aaf6f2392c2658f489b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1148eaf32661aa745e6a9c17fc6ed79b59531986d73acbe7060753475d54f68a46d29791dcd917ef5273913948f582f4a66a0d6343d48cceaac64cc77b466a80e39abf5bbeef6b032e56b45b5514da2f886b45271658dce198268d1488d31fc28930a2348c3c1b747b2400cdd1cad5f77fd3c512e94150c57fc474236aa1389e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4053585388cb487d247c72b8cbfdc225899bf4e5cf079c560e4a371914b2e5bbc33ebc43dd8b9a9af6157ec2b8e945294faf806ad4be4a401cc10657ccfd3a5409bee2d3bd3d6c7f6c53e8cb68ee6cf887a8be1fcc96aaf3ae182df8aa091cf92f43eabcecf3059f67eb4d0e7bfa270993cc812622f7c945eb3f5a96a96e26f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2035d16595b44ae893b1ffb362fb0b166aebe2063fac4c78720d9cbed7114e6362bf4c3be22e0d25d7488882489a8b3d2c205fdf11b8fd7282fc36c9d893312e4c3242bc3522b2e7ac3fc6180a0a9ac836d1d9310e621991b00a0c3905f39602cc0373dfc38badfdf850d7c2d2eefaa3ab23efac411ebc1f4255eae3ea5bf663;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f4959f87b2a2887d5e24c6ba42ac4a6973547a88a1b5ac83e5640cc97126b1a27f85ddb24e1cb10fcfa604194059a11fa54228b57c3b7984f35be3a4985f8f4cba9c7115efee50d7e5bc8f150552f801da250554e9aa9635df1b825b2dff6b0c253a9c1191841bf6c0dc4ae3f4e94a1d0c2f9f03cc4474390b5454c611e9d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce3f4633bdb462b1123a92d044e4f4403983cb297427381b7b6911f529b0c9f9003a85fad1d0430b8b847806b8067c1962b269899c0c6d4bd8390b73eb3210036da610fadc3d630e5bb9beee395ee97b9687d421024611f5e4a432d7e9e5e3349999836f08750605616b79063cd8ca656369256d8f46bf1d7d44e57e38c79258;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c7f0ffe9d78000bd97558b47429c2e7bb2d19616d19067ec68b8b4b2a4440533fb398c494c721a62ecef96f04fa9ba34b0c420fffc99d39cde88a88f2860b734b781f394fe43649331ac75a5745b68e9b6afe71e7856877df8fe9c25ac8f8cac6e003e27be5f22bec9664f0fc2ee0de736e2d591706a822eb8d0a76b31f77d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4eed909dd49e630bcc70af290ba9a3372b8b3e9f3231c0621840da0a7b44b001f94cf0c22f8fa95b451204194e16a7160b6057ee687381c55af201ba5a3ff3ed8dfe11fe3f71ab5bba704597a9f0690f7d337a0d00113610697ba0c517a92fa8fa54330373762560cf2aaf9c5b502429c9faf58cda46c58d8391a7ea5aff4e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9673559654b4387cccbb383996aded2b1814abcdf33630a2dd52a3b09fff9c196baeb6cff71f9c6e2b701843bf2c9e0da6faa858aa180d5cda1706dffd228b80ca7694c114ba34daf4671922bc7fc369227532a5b56a31c19b5631c85650541f27b31299c062beeed2a78a6da1407ed3a40e9503723d3cdc90a6502a05cf34d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc495759cbf3e6a477c674b8bc16f501b874271f0baa4ad38edf8644d9709811031ec7f3307ba1c7172cbf6d5e991ef08809d86e0177372ff0c8fde898816c55820efcf578b6b231a7737dd74fe3be836c078f6243e113e905ee032d96127e74f8e25a81bb6892d3de8262c6d5853ced18f178ff18da99f12e2a89b0c5a9258ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e162f35a3fdd65c84d48e3d8a1d66457e3b5fb2000dad3a616f4236a0802f7df79f1bc6600757d1e940a5c3980c61d904da52dc2758d666f4c421d65c3c1b5e59a3edb68d974cd0a6dc9caf9714280e23099c53ca58bea9cb80e2a5e20757b32d7687be287fa4599b8f8c14d38d16b97764952661f64dac90767a02e61428ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h862eeec746b2ebe26e633acfad6f5606410e20e3e88546de24f67639211f0c2a5801504914e54e14a90071689f7be9b359a2dd0aaf442084d3a4235c3089b9e4f0ad344d378c6c4e2a26c3a01c919ad03abb20e57d30c3204d044e1c67670b472639f445ebf61f0d431f1965fc970c1a293c6dc5bbf1379bf9ff17c1795209ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9c3aedc6d9c969eb7d8f72880fc7cb086967e5ba0f9ce588af84fea7cfb2678aa2a8ebbcc97a2ddb9e032c4ff8be5a5107090837cb37472e2add6303bbde5177d844c2cc9fe0ec1e15d3dd13f332a7d6a237c8d6908fb9f747e2f8ce1a7bf085d9eb8cb6530022cd80c316b8ef16381d114a2a905821f859a11c4fd7dc51769;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9941f9693bcd35f3778a5123947aff1e3abbef2649eeb41753cc87c9c9a62d93cfdc6a387fb683737d9ea2d407a131917af20eafa2c366dcfcdb33c179fb12ffb46b3d061773330823c6f08bec07ba58a871864e52d9ed21a05c968125dc4b5f7653aff2ba0bf6087b6f4a8a7ea49f0f6df36f16a84b6c01bdaa4b7169b302bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f7036adaba8350a1608ece83e69caf2eeef85837edf697f922b4090725db05bf0bf2e86bc45a5fbe5c9ee07aff2f0dcb795f99751e106949c6bb0eebf3ed122a8830e647fe239f77ccb715659d86a2711d8817e8557313d2e81aa36288754aadba30758bd0cf758fea66245d7b956435e3001eac314cc476abfcc1f08e0033a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7eadb11af26cc024b38ee50cf6b469cc175e114b533dffdc085077fe2e6434e91bef7f198ce4d28a45a86c430b24fb27505333b1bf8eecd97c0a4fd0fb79ac97c34068607e8860105b980d4d499d43bfb153202ac73873a85857135d22e48967754c1fc38130d993cd1bc685cef5dfe011357305f41b31c6b8678692e4e696e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bff4b87cd09c8073c86b58141d8e907a96eaa2fac6d9979a113fc536bdcfe5d653e66352ea51468b6cf4054b1b53805548d192372da3c2cfa8cda183e9049d0d25e821604cc0e89229d7faa35df2543491dfe80a2c8edcd8f50f6bf542c3e1be1d6db57385acd5ea403bee4796e8884115102763eee1033a38f90982a09eac7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89b87ce175370c2eaecba149dacdc30e31fe26a926dc7571ebddb9ed0dc993afec5549383cb856e7b7147fd38bf7d61960d81df236a5d35b2ff25ab3ce73237dc873cf63e48f2cbfb0e43274034d698ef7e61d62a8313a103381e1de725ad952c8edd3859b39b39179ec7cbe71effa72b5771bbcaa408bcf7149aa7d27d28602;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6068327530e58ec93ddc38fac7f3141306b40221e157cb1a87a3a3eec7fafa7a540bd33716e592eee05f6cc27c173fa65ace5657bb9d84345724fe97e5921d9091431cd2275e1e761099af19cacdeb93c51211cd00570e2460db576ad3a70a55097ede87eb1d11e499cede036268a036778573601e7957f421358ac99d59d92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fbd41cb53f2bae60e3e0c75ff8090d817e42abb174105929817190a6695767997c149ed109c6e73685812566610ed488db368442b2bcab328e03f1776d2569e2306844d58f6f9b87782b2a2315ccf75a56cf8d275675ce37c835ab8c95b0ae370b689e5c87b28b89b2077b3eec6438094ec06fa1c0944de990a88fef5644354;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd34d862c21010b85a80a5b0df93009fe61fc1b4b2eabd159935225c23f87fa0b82927bf50dcf07ccb6ff2afb352cb11fbddd7b35b6a386012930eb959921d5b0801d2c72043708bf0f0f932050eb90cfa3b55416d795c4e331ceec9ba84b696fb07d260c63ecc67a6e322cf4553b6e205c8ed4563761aaaffaf5e04a0b2133c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2623acdabc9ad3cd41e4c939aa00fad0b4f46a28f6469e959255b4dd58e3ab1ebc2820fdabfa101bc2a4be2007a2e412b6c85b4262f1ea9b1690b9e6e535c082adea02f3175919f397ae981b57184ed461e69c48419a596ce727fa64773b0b1e157456d74eee34015ece36d5ac710a6813582a33e67f4b311d2194bf79900b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha11a66ae8b7e4e1fcd48dc94851bb9f4264905421ee4210b052892c0afba60cbbc735cc73838b77b2f26f80e9a9df42ec5d07bcfe051e9658e309f76d8f8ab07c14f910054972871648861b750ddcc3af6141c316f59c867daa3f7c245af6112020880fe00b85df09588adf598f63947e4e955f9f02343d4825e0d9d73ffb17a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34b19fd5b24faaa508b3374339128a9f3767f7aa283a0d40f26b4a45a6207ea27e092bc330e7a5c47370d61ed47e8f0db47a3827c2c44b98c3808a2378f8a85827888069da14b806f809ee63d0fa91521d667c40a9d99e275b39bd0220712a7451035ad4d626d7f8a6158609e96aa594163bf1c3189ed0c2d9bf6a2664c0d20a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31c4b4d2cfa9687d7f56f1da7ff25a4862d5ee35baabe74012383fc11dfe1454c6511e5486f6adc11b59f734cd40dfd2699a967edb915eb8336064fbd886d93fef6bf79e6117a6418da6f2063fd56c549a6546d45342311c041ad7ed855c4a9993dabf70e71acae0f7c87b16d8656075befec351477e420c38e70f6214878f99;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13488e38f79c1e3be93949048b49e18bbd1ebdd0ecec7ec7c5dcb36a1ad1a1528e23b58a83e28d386bae3c5f0a0127bf05c4d6ff3ad17725ec9bb9a8b7ba0c9403e0f736b93d1de7954d91a11b4242190c14dcd981a3a4ab0f2e4381f951be541d6dbde44237ff443d5a3daefe57e8e31225e8019ef0fa56a5ffd9691b3e9499;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd67e6f2ce583e6bdb3566e6289f1e6709d1ef204b47f4a4e9158a9f0a36a90eb335ccd24b10540a00f82904c54131e2668c7c50ce60dee17ae00f111c15e9b42f60b68de619e23d6484a6073a616709dbf4c607bc4a96cb7146b422a600485d7e60424dd4fb45f51c094295cdc6914c1b46d207cae428a79f3f1b795eca82339;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c2e9eaa21295ca8f07ea776a5e3b9501f2ab2eca6aa6052d0e30243aeffd1da84d6d847677ee5c77a3ddd4198c465734650f219f0c12ca861f1c7308aef3340db850fb8f14d3edb7208f91f49feca3ffd0ec8262efa0c6dd97ea5e58ee3ef12799cfe17fa44602ec5839e5c020b6319dc3b2a2d5cce20cbc0d84dcaaea1e796;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h679a6fa55acc4d07d72d17095cf3618737319a55e9440d0e7c9275ae6e536092129fd94f06d7be45f33fd12ba34f5065dc9f040804aa110f2a9ed869774e39d40de2c027f33a74b462668ce773463ff67159663c838f9dbf3ff2afc4ed45f27b5901cb5731ec0e07785f36fa8226104dc706a241b2c32cd0bf0d3e6a8e0b5724;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h489b5116ccd2ca3ac4179d252dcd065bbd9020a36f4221352b9634af3366f33d051f44b62a182b44118fe17f86f069fa4c557a0e991c889cf77bc0c5d0591c521ec474fd7730bf4a19f8413e1a6267e9e4456357af0ef1a5462a3f81ca5a01e87f0c3c4c5d9476f493fef49574f3ae5473cf93d73bb798573c2c8b784bd6f171;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7f49db365e3e84f678ecaff4eb3a60ddf31d07b17495e2fc4ad1fd33572bd20608ecb17b887d695ee689eeb6298b3dae0f4d761993573625ad8a502b9490a30be502b6f749c6aa713ecd8828e4f6bd05fdb94f3c76f7a0140f1476201814705279ae4eb7b544bce5923f24199d8f92dfca5a2f62046181010a236ae288d4655;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a329b6e9328ec8704a38d7dd105b394ccb9d18f529c98f74fb72a27608012f9a6a6bbcbdd0015f936887e437707671e0c2484fdd7c3ac7264a49ea55a8583ac261bee6612abda0b8321890e98ede03bb61b1f9cb57e206c28feaa36655fbc172775bbb80ef6927df311687149061e8d5a58e467d6e5089f8cd7bb781b13e00e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5aa52a322423f196894bda35419ec1083e1b80bfff4965864c796a701b803c1cfb56d857a3e6e68291c2511ae71f71b6fb5dfb52b38595d4d5ee6e14ec1a052afef8c3f16c68607238bf1456c021e3664c7243d678999eb3692a10b625441db6c5133042c5c006af2aec9e0bf1a9ee5d2b11c53d3221ef30be8fc7df624ab79d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed9a66e1fe67d01dab3c5abfb1f9af35fa049ba77e0af9d69dcf984910f63a4007beadb941b8dd8fa355893cd2857348b3954fbe262502d65995a112894c05d18af895ba32e861567731e339e13d0e25a35eb4e2478bc9eedd9a5cbff72510f6009907e3314acca1aadd4770605faa1fd2cc3f316804acb75437af1a50cf9297;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcf0e5d3aa474e127bf9c50a397ab206f42edfc171c9c12cb4c925c0d5f606c5da4639ad25358c487edec073a9be7a573855fde06dcf73d9003b06e138b6052432f1d9f747b62b3d0c33fde9f5cb41b80ebe681a4366db07dd6ab4c50420630e954cc0459ce7d58adc18d09f399aad9b38c4519dacde06311a19d4e89fb17497;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fc96f263dad1b2c1a8a917981f28902afd394ce086920048cf6230bdde062003bb48e7b114f60774df6c1899324d86735d4e62505acd8251e2a8ad8efc67989d262f2598331e11b0b9ed3aedb9ce5102b03aa5200cf69505008243899957629e373134aba40159b5250fbff494d040369bbaa5d116f0a2f7c376fc6ae6da7fd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bb46f65d2ebd2c6d3dd864788f87dd4c731cabaca8e39c70d382168c62cbb9c39de23954e72092a27a1fb00676a8f73c22bd6c60112fe38761137df9eea6fda1506a123435b23ff2cb2b182da39d8043669277f3148b253ae9ed4326dc9da7d9aadd783bd92da7d0f5cba99087d5b72f1de57867a12e7699344b3b4c855818c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82c3ab9124309f663350868daaa99e8c5dc3ae7d59c6458e67986e80fc3c832c8aa78e80359a7784b7538a1ff6ab79e99f218767ed462579e036afd748814ae6d1723ac37cf86a3c00e933ce38c24d3c1ab62880bdaf4ff89f8fc12433d9a32158b2610541c1fb739c6b327df6b1767c8881658e141d1c9326a1a91461b4fb30;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h400cca30b9e327e0fa49829c496fedbdc174a71e681513a8a6dc5942710584ac864ce43b31ccae11b3631199224db22f2c29a98ff6aa87684853071a0955d51afa4e92bede2a323dd1e7a22d6e5a082c092bbb05fb85689fba0ffd864048a89fd43868fbd09e56e74cd36673cb38c75f8a3350363e0bf1d43f608e77cb1ace39;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34789064eb00b3060b322b179e0db646ec6d7439680cf988762def310b9bc2bd6d99071350740ee543c72f381b5bdbc393054db5299d0172824708fc3876557bddf2342a0b3d87c8475bb67926ac58982a8ba3234d42a6143eb250fe7087d84be5d47929f23c813e30198386a5dd6462c8d5dba641235312f2358908f9dad78f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he83c80014cda44fbd668525b2c035925817c612fc653fd2141b17cf6da9be27c82cd4a7e2274efe3feca2b07d1746024b0ea490b5976ab062c54be1337eb61b0c92eaee4bd4dfe72e06b82dcace9bfe043100e725c2c8b298188450c5125f167199897c6dc5c7f4d49cb3af7c91daea010378845ffb725988f35282ba9ad360c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cefb96599fb834f3a90b12c5ff2e3c58f9f549005851d215706fe1be12160c3ce068854de2a8d01e5f24d64d77aa0e6395a70a77f19728a44c4da7581ecf2367593caf73d111bdbcde78540611087aef23ab461a6df987728b9a21d89cf12a731cc11ae77b9e44d3ea51e95950a6006805e0115f0d04b356d150e5fbafcb2c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3480bbe34d07ae997e5300656dd7d68de0ee88bd86c7d23b013d992f8e942e0b1c227195f814d32d7b26e84b0e44645f444bf82147d0c9e293086603669239523e381012f08504675b3331b90e5ba4eaf19d37313245cd89f3f5988f40ad97df5528aeaf88655b2be4b56e42cdab10b3aa1fcec53031cde47aa98a37f98f8c53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbca3ce36f4780afd1d30ac3ad72aa1798aa7b75ea33df8980790ad50e9d601ad78cf22ac18aeb7ac22b39d6e6ef2a32f222f9ee21746290764c5930c4f4431151c01d34ec55f3a4fb7f8b9ce4f4407c1ffc609728e04438204262621f7339e41b0fa8d9417cc9687902dcf70e51447329278b8682d84f2c718b91531991ec244;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a7fb378edd1c859445be723dac57eeab628a8e70752e6d8a14d2a0d6c011a6d2dbab8eb260c61dd0d473ece754dabc67776a741cd6fb8630b7724585bcee69f59ef261b8c416686b147233780ae9cea43458cc8791ce8582dd3b59b171a66d999e52f86b97aabe8e8c98d316338cbc4a044d9868b7448abac42410f1fe302d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c74271f3b60eb75f0ffa074e74b2dcac59d3123f1fd283956ea56434f8ff0a3571f4fa4a9eb80e572b8e329fbe81d173f6af3f5112d08ccb7ff64b7920e8b4ee1f34d69253b447add7cf16bd8352906caec61dfea8d713de27bb52b5a3f01e0b89f868251cdb01ef16cedd0c3e02e8967fd5afde0b2d986eedef411db05a66b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30bc863d3371a9dafbe3db5641b9217f497f68829d13f6a44c02a918b2ad7d451aebf1b258be786182e0af56ca7dcfb5a12ed3e90331c00a26e66fea2a23db8fca68de0561a798f732703e70d3db957ada34d59df6cda0cef1298fc7b2af2a97da2fb5e3b5b849081d911635d0f4a70c85c419d213f2e1a5bea4c6ff0ed09769;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f84266d492e06094cfb120150ed2ca444cf80c58a888ea6ee407682055417e327049fd821be9bf8a4368657f9c18aea952f42bec20afb01c5962b112a7937bdb52be2070d8100c3024d502667d25d06c168e1886a482ec482b7bba55de4f06dd92d1617cc747532ea913a17559c5e020be5a8b83434703f581937334a21d80b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebcb36614a76d3dc32b049d6807a766b74bc973163c7d7521688d91b8ae22ccec0bcabb49ce46c3b4e29f1223280d27e0b5d5a344d4741ac94ccb7646fc4a0fbe40e2a6e7bb7659aa5df372915d6886161915dd774b6c829d3ba11ca5f7b77921d9cc6a375758aa377bd776e600d5d02162390205bcea990eb934eb642241061;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5adcf0edd447cde86c1ba263622b26b3fcf0cdb7a801dcb3c2e271339e8cc521e3b22abe359a7df08997fa4e42c9378d90022d5c85994ad9c616e807d1778edff1f71e486418ded4d4b6b95a81086ca6643ef71f4d1c3c919639f39850bc006cdcfcea7921e6218dbd377e634a0c9694716119ad06ad25c5a97dc87d048243f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2af85ab668f909e64dbec3a08d44d3adb9378b9f764394717da300b654d9e711a2c9ba60faa81ba491ef8764c78d3d4638f89aa15e746800efd3ad32ef0f157870bbbe7a67cc010b8ca9aeb70df5c44fdee6b785ef308b7b8399b930a9080c5269da01f37199e70990d82b05fd0b31e3a01d078c1987eb6d2d0affa3f1dbba3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81d453cba9309ac002c2b6327b89c3f1ee3c3339dcf686eb67c2793a780442563356aa4e3de247d83bb1d476ce4030208e51af5658f0c8f27e5ce75580d9bef346d0fe77b368da80b3578350f10356c2d5c0b5d22b78d47af738d171d13b9c9bf2b8efd78328199704d68b7894b8ab426ab8fabcd425f9774bf72a3ee576daa2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e2674cb48bd742b254a2c783e70a7643a7ebe5cf30f6520c1a0ab3bec579b23c3c195293ad6eadb302737967e929028f50353d1e38ba280ee7659447cd8db029bf97744a97c0841f087a0837449958c15ee271375a4e801db4e823ed1277fed5403ce687f87bfe762c69d809944727e89c049998aa13392282f87a5febc9f12;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f195445834e829b96ed16578434fda392d4894ec35a62c3fc9455f897d15478c156bb1dd1aa5b9c52c914c06abd977a241e255b083d9944c55367f7f5825838a35e6c9be30e3af741aaf8c88854602518d44ece20869719672dae0f4b1705d60a20e9fa089d5c344438dce8b16853aabbfc22424b8acb0f49b3447cdd7576e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha32877dacec1b6e7d58dff422995c87fa70329cf40440f5471bb3410b38d2575a105f12743081cfe890d6ce44a872926e9ac3cc93a3495de1808831b32cf94f002bfb7dba22c9dd0573f11b40c63d9919672441e715d34540d8d24ebbce6b40bf37aa6153a26d40a94a2cb21c88020c7d730a421bf4d7d96e27d15117b15b8d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5232c2af2c4df68a233feefdd8bc462d8633a1bdaa2b7b2571d5f9d94a44afb5b50e8cea94db2124baf8fef69787b2e3493e4319979b420ad0f7de9bd5038cc6e0c20c42ef52a159248211b4059224fc3b5e573c1cbf8406b92092c4805686f3a090fbb4b659f84a4f5021c650124d85fed37e6aa97e30b73da7c3950d747ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd8fb620175ee26865e034f11142eda46831ac7ab106721299d0bb5a653f9f1907f3986843deefcb8d94eb5a2c7bf6e9461b22ec61d88059552124986c02854f2198063af89ab2220e310fea00ca4d189aac16a2a8f5e2b420431cc67e4b9a5525382c177f59013da1824f456c6294f308e3d91afbffecd4b6af5aaa14c96d6f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heffb9d5d79ee7cc17a75ea6662a522a40fc792eef5a6955b4f67caeaa627cea6c8ea1967d7c03e67b3a8cb034f35420d8a66cae8409eed40d396a11e60f75778b9c715e0682c0a716ace561d7f4b802ae37527fc68fb6943f807ca8c1335a5ddee934ad40217b17393aa5bc9b0d80b503331addeb94c8fd06da15a27cd6a415d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha12c5d308a297d180e1c5b12e72835ea07432d84b883d2a4611c4ce6ee72ab29411e8ab89195133c1041bafa90fc75845134ef6e59dd2ee14d7aaf94d06cd392450ee197a7f07af38cc6219bb504bbec28d45acb40a2953367f8f1ef9c9dbf5656f58c68d29f142f5cdd974297a55265dbc74b620f65ae358f5720ec8fa7c777;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he82371e0ac9fcdd4ee2318212170cf667c7e0b58c453b3926bc34bf99b26af98907819cd2bf25557a1714423dcbe5488b5ff1b8b3d7fcc4a26892a9ed10c9bdc1677690b56b2c59d9657bc2f780979cf98a9a1e14cf3c1668c62144d76e49d33734ba5b27a020f96216e125d4cac5d93ac96657688cc2f76b9e0b04caa3cbf6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdac6df0a78b025634c28b232e04999a2aa0560ba3b68f58bea6017344e6de15a10b5cc1bf3fe9f18579d2c2594be633659127def52976e8885bcec1f4449cf3a647dcd338600d41b07015c804bf20a28e0aa06ca329e4e5754bfbec127b54d3003c8f77e237da773bb34dc47c60ac9017bf4f9dc06c7b2e357d87e472ae3bf51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd82028d4a87a1b5f05592e4c9ea91bf84d14d0f4e57403634517306da5819ef099a559b4b5f36d4554a7e03eebe542064f5f78ad31e027af5943d9c7e9a0f77f13c8dfced95153b13c7154f51c16f0184aeae916251152eaa887ed5d05b272ed9aebfac7f8fdd2c7f300264d8532eff4b55bc0406488a4e6349420982d4a3912;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf540e787c7a714bb1b86e7416d1b28ae73ef0aa1f166d1c9dfe6e030c69180b1e12b89f65569c8a66cb276e43f2b97adf96df74174909483cb228164df2640b49e9cbac5996d1e35d66a793556a24872b99e1aee919cb6aee45fdd6cf5e89f51083c8e8cca40953fb24152fe96a5710a7ad9e79e60bde924980a88afdf46438a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf905d3fb89a513554e65bf29d54db818a0a7b77d9afec1f72cf002fe25cf7a9f23a33041dc038ce8eb4e43360b03f4fcc93b7884a3fa21fb2ffcfebe55a64c2de14368937f0757925ad3ef8a320e4763e4e7fe1d40bfcb95c95f6f4f53d803e22623f5c78073ffa335e0066093aea89fa9a30ee8fc96ac46a4a50761752fed08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10602f28330a457de2c2af581ae01cf3ec4248b0410762df836ce38462219865105a1a6c277b87122c29af64ebe76a6e4d793b29e4c82ce2acce0ebcef701e98d8e8d6a9141b7b76ee476e75dc59fe25b7d6a70ce4b8e5053b48cbb987a0be7489b59d1b858125efb07a64e00824b88339ba4b7ee802a0df6e311ef95fa1cfe1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb57a09b25a91b8eb63ce1996714788f207335da2db102f7fa9a78ae154c2ac15bdc009089ac20bec4a75f6cc7135068863b7bb3a94fc3d5cb2a49758f401c853ea64399a08e13c0a808a71d16a57d068f3432dcabc185427b5cc99819221df3385a4bce2c48f484901c17fa338469fd87c5544ad718332ff3a41170cb63c0b75;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6d1c15456c0ca78f80d08f1161c26bd7642f3af3934fc70e66b827af1f803f2dbb3e6edbbe8c4526c815af9222e308c94ce389bd09d71d1b097c4f5f1ff8ebbf17eeb19a0f9ce1aaa5ad47d76486fcc65728775eb6f4e04df9e368d9f070ac0f2d8af05672b2c85f157d6709a15a8df94e9e7b28840df2844cfdb67bceaa599;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf993489bae934ba0fc5a4e111e91179a897435c3caf3bb27ac8c7679a32491bb82466e30c4394b080f79f019d6243a87f9e3dffccd870db3647b26731d72cdb3ef4ce1f229e01d300b2a69e07c90a786b35e4f7edd4b2f6570f27b59c7ca0d935df05920aa85dba7a4a9822f6988d71878ed6a156ef2525a69cf6fe81fec9893;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbca3eb284c554c3da6167aa9b7b5dad5c215a6b4d128323857e6cd0fdcd7815a1071cdde92f531d02781b63c7c186267892178c63b52eb4bd39ba2aab837fc46f8015395e539d79de4e74afa0d6cce71a50edf7ce5abf3f665f666e4f561993128413f80189316ec7af334609907a53d7727d0532cf618f892d8b84b911796a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had25eb0ebeba7f96523201dcddfb5cd48cad0c4caf76f78f20ab4ad93724f55b43fd56b15802d61d855f6862cd355309d2a569b5678840cb180c3e738cb554e1b697b09315d7454f6662a0bb2454551165f3629d8cec420241a8a8b2cb4dd761e13b02db397550bf443e6c1f30051aaec5da2858bd2c5dca1ce4608a72c8ac0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha432cc206ee2e120d656d3ccbdb5eaddb941ad359a2beb143b0f3c3b768569393e51a7c6ef0c3cf568e266e1c89a0078bbde546e81eebe0e38a0b91abedc6f20eb8dc22ce2b443ddb394ebb14fb1e972029709103cba92c30ee0f48d132bdcbb9c542afa024a2a969d4c615472eb9fd64a390522b85a104a54edaee1aeccc85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdca5a3e1dff3adb5f0a90d4bc88a3d6d2b0d8256b1a82be8efe3d5a64e81a3e7a419a372354172b381c91cc2a8093ee8e5bfed8474303a85c46cb9f9e10eb11308bd6caf14b9d349d2b751120e2306d217859593d953db2487bbc8e71e7593ea0f31cef99931398df4c10f6fda94d6b1482ecead1d71d5c832b60af2dbf97503;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde067a9e62cf58fc9c4e8aabf65afc681bd34c60d152f0594deeb9e3da67fdd03b2ce05d770ecc0ebf822ce7083381cec23b025406124b1300a19dfe1e258fc498911993b5fe436a507cc298273e7da37e5506f1c7f4fe12448a0a11a194ad0e370d264490e2bf89e7567f43dce78593f68103598ac85816685e86866a84e74e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8593b81d8b9621728553a6fba6140024237cd88dcae4b47aec3062dfb41a1d1576fc59912521cff346f061ae5c3d28e0cda341ba086821883b66fa419b8105805e8dd561e5c95b000f74b572b4fa81973480efa31880bb409a40aa7f1fcfe37fcd7103e1501293bcc432b01f0b4c1788b3955dcf5d84d3a366392745c71843e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf19e514663741dcf9783c408acd33c1a9f479765c3bd5d1ff5d1821ee6d4c1ecf94b818eb98cdafa1e89e1b1933d2d0e514df590b5c9acc4d37368dfad96b0c5b61dc36440c4c8ef20b50336a3d7b8248b21f16d54542004fee9a5efdcf4d2ec8435aa4ee21f23ea31df9fb33378fcd4ab5c700f6254ddca53d7830a785afee7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9e25dfc4b168ea98071f7b098401b16a5cd1c5a5fb1f220a0e16a43f56e9847de9cd8f97da923d96cb896bb7e2134884873eda1a252cb013c23f70f0305267438027a7bffd62567c4a4f9c5a1681c3254bf07116f6e922e4577ba553c7d5274ecf8009de42bbb05bdfc4c6fde3b04309a2ad23c6e2a83ec1fd27c15661d683c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2de6bef7b1d134a76ba66838cd635263cf73c1609a8037d8700e0d18b63c81f8aff66efebb036a03c15450a21a389216ff3062e0609581023efe09086ae6c1f2b1cc1ec1c0e30dc9bd6c48a0624473a7219f7cb687e9d3e53b51b1f45007c4b3dd1f0b71dbf16a7b0310d02e37b6c36a9c660fc6e6d87f4792fef6dc1759b6c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b867790d1cf5404140e364be78b1989c2e67800dbda03ee3037eac6eebf4e247fe262b6149fd5fcb0bd544daab3b7f80d3c84d089ab174142f04d8c5e9107bff2d6df9e27487bcb787defb3af1f1ee4207013bca3c8478f00323df87589f9a3a48bbf11d39731398e5c48a9b3f5ea4ffbeed2352d2c5cc6ee4f2ff1f9e8dd4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12ec358fe717fccebce105c782d94854e0689769fd733786dddf421bcb332920c6e92a2cac6eef988ee3fadae9797ff34dc509ca77aad4a03218b7186bf6c3d69a71a14ca9721963a02377d823eddd4c0212183f01038b10f4f4a6639295daaaf8f031aeaa5ac67e17143ec7f8832ac5c891c85df78810c249b16681ecceb88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cf82562cf7c700951aa97f743fc1d5c6be46675fb5008cbe48de7105ca4b2f12cd7593c72c26b8560108341507fa208f8a36ac8d408dbd2473cf68949c8f9cf9a3654af9062e88fb511026c542e6212d7f6617fcecdb40b31e157d444f36e60d30a6752a87b2314db37e8ab4d6a7495e3670a112c3ddd43477fc083b6dc8078;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bc6fc09a9a866e472128a6044b5587da961c0807f122027aa2042fbb83759c299fca014df1a97bb90110fd1eb96d7c3b833cd40161e50ec6b532a103251fe5b28fa2635967d2187ed76d65dfad22da21181e98d68a89e2844e661ef03c0f04780855645bc653442a79169699244101a1591c5f1919f4ceb768400afe4127364;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88e5356e31d69721dc5a68a777059759cc9a7121e63c405db2920ce9aff015a3d8a49a70688d185609b3b3586976fb1534b0765190db5c51774fa0239e6902c8334fcd9c9b0f7b8afed450f48fde819ec693ee4a1350c321d94d7549b7efe9b4d222f3e7bb0ae4d078207c4d34b25ac6902b86b33d49792d60d37399804b06ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h661f83adf0c480a1716395196d3391466480c3980b932c6931bfe128949463fa5699d5a6d126b828e6dc9fa7cf328d20198a39d9f92cfb51e817e8d2b1dc4dfbd014f2c6a183ccbc820a0bb64237c3f813834ab849acfb905f31678180d45c9fe144744f5e64d3a4bea0f5d7a430cc151894b482a3d21633d53689e3bc92d5cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f20f94d1a8008bd5b31c43cc78b67dfb24d69ce6c804dfe8ff819ceced32ac62ffe6bf80d6af566defa96806bd068d20af9326ea057f03cbda05a0686469f58da15f9c0fac0bfa5e497245f1ddfe489dc2a66f24f3e1bd3aacebed6088a9ffb42224e71508b513c8f70c87452c22f969eefb9fd18bd5a03e120d1672b2cb571;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1ad80f34a48acc1ba1d5006da985212eebd743ae36121f3a963f73f0466d4826064a8ca967a0ae3ebae875b9775d945bc0a743d31a849cff4775aea41fbf1ffee16f26681f0b9d836bd6d9c06cebafbc21d227c5a85b768538526d6f6f548a9ec0160718e68fdd54654c70bbc0ce8708f3cb1b17479e282f155fed158c560cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h738e5c56112d9ba08fcce5354632a2f95a5754151adf489bdf541cb3a2419a51c3ea98bda61a1fab4c1122ed26477eef89cd25b369df5b25275b52589313391082737641688ce965dd4b490cc2abc225037de823f2fe86f975b1a442be701d71923ff2783cb14de28c3925633e3a90981b24d4b035b5ec9087345291568c3ab9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92866ea09289096b7ab53c75268fce50b3da906ab8a31107be32ecaff067f8b792bb954fc497fb3d5dd602477131f67e4d5d44412bc9321aa92e3fc27d2d536548938882b6438b9eac1629054579b3975493be8c17506223d2b8d81939a1278503c1cd537d03c4fa7bfecbcc1ce1604904b6e10a9771a860e8b4ab25ae6e0ee1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8d5bad1ec594ded0e70c2c9e19c49cb10dd477c4676fb8fbf3d4f980fb7ef0f5b5e2daf3f19e037fa8f487e7610327424fbc02f8364e4da57dd2aece39fa7a445d29570c121d34eb41534b221bb2de764b50b57aa70bb018fe59526f08aca45d0039b460351aacd0c15be872ad694fcde117f90f62285fa3f52d211040b041e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heaa36ad7cf9d9a09ea6b87b806e2b41ab153daff045b5b600669d7e4c61f29abe203b7d28c7d4b0e6dd0e29de802d0d7bb15c7861e8ea74545c18cacdc1abbeb809757cc4f5588946d474c1c5cbd91788ad6dc61652efbd5ee822c07b7db448d243152350a44a551b88aabd8ca6c45ecf39cfa9fb27cad84008fc8717d11930c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55cf2663de9bde00831ed378986b84a60f64957e228ee158aa419e9cda39dcad0a3863472c81d8f1495f7489facdfc4e8d6f31328c068a249593078e62b49a26116a1388f98da4c319b000867b0f6ff998603c2832cda398af0771f5b1b912832aefe6291163516b84b9d1c59684b42f68a0b2977246d4edd43c4cddc6951245;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h477eda09c9dfdab48148c9c93c54dbd8377c5d654df6dc6759c44c347e5a275ed53a9840abd7cf342db1623355c6d9c569ebb43cd64f1e23b253c7777c88a2cf6e0c91ea464ba751c344826ae89f551d0d0d2599fb382af9366f97f809662eabba440f49cbf4de584a60a59e7d114cfaef9bc6b52597c037a28a473744e1c9fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b265010b330a233973261819dd0f633c41e45c4214722b414871d0858e33c5749c7d73b67312388d65efd40da99074ff66eb93da0e126105f70ff6bc32d35a1d999f53c8aca9fbf609f98b5a54cf94e0b85b9b42588e7612fb6f6f1bfb6e03962b78ab9069996b8dec5485a6ab811536b8280683e67bca7442ea2b75fd22e69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h798e689ab6e01542d904820fb44d4537f378cfff84f0f10b380b2d355112f55b106f6838b5e99d6cbd34b317465d79cd49cd66831caff31de1fd004a20fa178eba24e0393a3693c4e1d1fa6ee0d6c212b9bd2f62b8effaf9992b61a938d39fe205fb6f87bf0988e43be179cd02429ec8e62e9fef485aece60ecaad2b4d8f742f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e1d4ca701b04b0138f3869c0c2fc6ad6cceed716bbdf820b247e6f500c243e0b84ee4d614de3f2552acb66021cea7f0223e65e9071b67e12652925062fe86c6dfec2fd978e7cfcea3732a08cd21c40c2bc8f41e1b4a60bc96168213f683440b0d1af377f127b09c0525cc51554e9963f0ba0fd4644987eb22461556eff5b963;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6fa2ac7179bec8811a370225515af07a60c721de3e9ab1e4aadee6e66e0db97424b7f30c98c9a1d8f57baeabe00a1efcd141b10d19fdf5f3f74b7914d0141f5468e64ec16c39bab32b8a20c66430c53ee5b689737136ee6e8ff02775aa37b3ef77e63c39948fe676e67c54945eb60855f93ce368c71f67aaa5955226f89c0f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f7704a69b0779f48e08ce2070b428ccc794e5a8bac3a3da721505cbc487baaa49c8bda3295b663e93dc299b609419b8f59a2b2e7895e614d18ac1e5e85ef96aedb34790c5f536e0216358244153dbda00e667b5592dbd075ca386bcf07859e222d4e44906bb1f450cfd937ab1a1e4ed12476a46c0f177c6cc38bb67f4f05d9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc45bde3c0c4013f23f80bf70f9a73d1c15196b2f2525a7f4b3968c03d2e01288162c20eb03d2526207242bca173806df8ea8c39d23ffa563563baa83c3589866a6b77ddb3fce991bc80ffed956ec59bf05b9fc3c6dcf6949e8165741f6ea67e941ec8bf82ec5b76d9891dc8d3e19979487a1973333675af5272c6745a7692e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95ad20fd45b905b1bd47b0752c9049311b16402aeaa18c37ac044202182d83885d2f61d46211edfe51be23364030f22b9801c8c367c09d4443636601e07bd1f05631852815a856b9d5c756e6f860845e98ff4b7a888f6ab6a47bac9e2cefb2fb9ebce1541243ae5bb19549655163125ddb018011f2ff3ecc40a59a071ad7a45b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cedb363e2290f574164f7f373bf2ebf5a1e0911172de3d1b22c323ae386cf16d320e456604f4a678699c8341ad915399c3eabaae071470f5456936aac8f3142cbd6dbf2271ad35bd232c1ef2aef1ebdff17c4531be8bfa43f51d7e65095c0c3c0bb51e1df87d00995b6c0e8753779d22d0c3aaed1159b709c2b01269535ef06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a74525a826bc84c80e9613337107d33d90629f991155078fcf17f6956bd53b39a68eade6be774693a33fc06929e3b59e46f361df3d029227f1d001767ecbee355338c6db927f8a35cd2d3c4ac1b383660c712177c17644e1b8f46fd2310e91af56d6f42ad982258937469c6eecb055b8058798af33522a12b6334bdc667bc68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68772229f26f0fe49d30fabbf6affc834816229f28f52d4ad72f1afb911a6e8ceeac04cfe1e2dde4712086d2e08adb5534e09005e1a5377b4030fc48889610ade81915ad7a8fdc970cbf0790362bdc6b4f024b548dd0ea14105377ae33335ca749cd3e11dba31e7fb38db7d8254dcc37f715005757073d2f03730946c7161c6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h315b965fc5251fd8450fc5f94bc7c7465aff6828bb8c901b8b7fe7f9af1b4292a6aea5eca052c2cd84e8ff60fd1b489b37ee88c17a314ece97821eeb3f1f6742860cf853104545dc438cde8875eb41c47bdbc69c74bd32cee784d8ac01e5adf795a62e560b7a923c0e72af8f2e3ab8c120e8298822c5fd738799ed79620538f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b55e13a6a28e80f6fe4809bb8c307bdea9cfd3ef0bdceedd42624a0b50a76619336585ef0c9f0b26364c350c143b5c9c23d8ad546d390a8509ac7590b6394da3c97fa060a90d3c6ac70ab96635cfc239ca86b7a4effd4fcf631624a944e600777169e569724c8a4abc2c079137ce1d1eecc31ba683a3fe4c48bb34b733d6b46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32275022f3efa2ee1cad0a28a00b8fe65346b76b273c604581198ecc801ff1e89c5d6db9fac492360ebd96eba6fdc09eaac33fabc9b4ceda7caca1433c52fda1f87728f2c347a6832eb685e08d69fa81a2edee5e94e46b8f313c61d058ee7631c4821197b62e89a45262e1d10c41832d5f38d0f87906ed24b9aa16a655f091f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d7d4a9a0b8f53a49765f85c4e021789c7d33f68c29c94ab9daae96aadf46ce952cdbb2f829c7320d20e4f1ea7d160a56b781cdf8fe595758fc0b7c6c3d8ac0268735d034ea86cf27724a609c827b483529df08e6dd3e7eb3456cc70d6b36a445ee5de27b3c4494cd25fa33aa30e241a80b6898a927b954eea417f9316bff58d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1224dbe51b0abb67c77c4a3053208b27d3ade6dae0f927864d7015ca74255749cdcf1a5708b061ca69f2d30b0a0b3467ee4eafffc165e5517ce9d8607b9d9f91b9f32840c1087129ff19ce9045e72d5907972d0378dd7ddebd3f422aad11aaaa9d05b01a52ec5fa9e1996acaacdaa9ec0a029a76d1671017960103845459c31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb0e8213287a25205e6ce7c7a29c93f62a4dfb3d1976c833b5f2b03770b4c9ddbd12d11151864acbe6cb6fa904f287758effac892b3cbe5ee1017961facf7f3014a3f02af0382d7c119775e491bf2692fa51b3c134af3a888ef168c457520ac0291c2f33e95f5c1bc8c09bc40c6dbfd769dfc23a13cb4674d116d9d806ac177b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbecba69b43afe1382b22959c7dec379a368f26df8982fe5525281ccbe32a7c6340f462dd121d9616014c85e23ebcbd16d142777a122c7d750fc3e66fa1748b2249a293a3ccb4ac0c3cfdfd1628b707d099340432c75cb1549ad89f987315b72092efdc369f13ef1519f10173484782e31ae78eeab5c50a5c59f1290a04dd872;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ba55875a40408139e424beb588af4187e2b019c0e947d6e8900d8e69d54ce4acc6d1e71a4f32502137e7cb8e74f5d016be5d7888dc503251a68050ab6db853e62b8db3558cdb14a2cb77faa813175cbd4fed23645802e7c7d29e6e6ba638a0c3e97121648f1de2e09cb1c97ccefbaf4169f9ce8a361a913bf7438011386776f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha303d425dbc7991765224bdf10ce9b51a06fb5846e7baa43d45621e0e3e4408707307347916724175ddaf42f853e11c15edee646171db3ab1722c929508e82bbcd1efc96c50830183c2e904360d51bf83bafb550a600892231f477ccd575430c5137948189899af602a68b35a71ea20fc4a358bc6f3b40a51944313aa8a9b715;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h132cd34e184710e2387480a836b2af52d373a457acad5a2e02595c4dd434844d1ddab0b9a2f503f7a9bf4aa94195a29a72f16a887a2824060a41fe06ed962fbbea1978dd1009bfaf30963b08cc59b7aed4798398b0cc08526d4fc89a69d2db4e61c05ee2bcc0371c03017a2d9722fae7417d5db80736e43dfe1065a09a0c5014;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5433afa8278018423c1f6c5d8f2db97915821de39d039161deae8fdc8396814a1081b71d9bfc9d76dd480fc785583ba5fcdcf265a5dec7048d2aba29fdc3deebbcce456c929cb95df48afe0da73aca616632fd892318d64177d65625306ccaeabbd618241a7ecd1fe68715539f7317fbd8a5e5b6550791be9279f64f5842695;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4be4b04f17109c3f95ce4b2915ff0e486d2d6ddae6275eda029e7f48f42bad624da3b7f5464c0c2457d9910ac5d1ec8895c97ffb224c65819b7c25153a7f84e37c69093f6e8583543b737009d970fe9fcfb0e89f5649960410132f76d5bc367ea3e93b46316b29bfc0551d166d5dddcd159b708a0794bd062b9bb383809454c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc4c65dfab7a5cc78baaaff9dec9132fc9fac2e9e9e1ea2a75465352c41045db601c778bc0c92cfe8532ffba119dfe0543df6024323998732ab2b9e06d6c3f2c42f7c5a5a6af1fc931d51fb18169608e9acc8eb9e8287f7a5517e24a92f5a7569309e94d43be6d065b39c35b349579c44f4ba87fb4380d13f595335749af64e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92ed914fe549b1199a655e2b6d05da0e71dd67c5254a67a3b3e4b77d427867e68221978f2f2466649cea3b753d7bfb4f66204187b70415822b1f4785b82fcf312e16615514736f57e57604fdc4503b02772d1888ed39b0d223f65f152ef2c07efdac6e8c785ba916f93c33e57cf76cc4298f49f8047116c60e7a0c77ca720bfd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2de0086c4da1b7a4d2103af7cc1eaee7dd1b96d90566713b6646b04aa39fdffce1e28c8f85d553f89f2d4e7008434114458d18be5a40eeb93c882363bb938af74e3eb8132bc8a43a776f8e82f9d4531223743d4100281cb48ebe651290893ec376f43c463089337679dc98cf95357217b2242a2212cab8ff94fcee78d2a5e47f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h637c4298cd9e2ace2fc0a950fbbd4c446787148e5e445b6a12c1ef5f8308ad62e89d280c36747fd9be0a6337c177d5b71d0a1251901e28ab22cefd54c6220ad23bf6634902b0814a9bb1e977e56353f3841f58a666f1007698149be184bb9aa84b4033f1217ba7550ec85ba15c2023a3652567d568c63938c6a8653eed899799;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cf9a4364fc283691b1135c0c7c77cca3a0c68b5911e7a80b47d6c72053f1c6e8099ee3d7fa6d2df337e0f747b54c3503e0c3790a3a558526a27d2c33505376dd3210623afdc9c75156a871803e462a106e39e90a467ea60394455a44ecf3a13351b9978f697b62d943f07a2fc9a4e01ced4c3f423ac89b89355369b3a5aef97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd679f90ef14a472f20df00cf99cd65f5d0324f45d79e8e0fba505f0b89432761bf1ee19759da8fdfff489ac02aa9e7883700e8b516a519c793225e7c41c2f58a877c26ee302da1ca7465422f026ba9017f184c563a72cb32cf05cbc40174d100e8c300bf8f69c62bc8bf96133457f05008bf47c32e7cbe0c7df4d7a52af5b660;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1bd56c13c569556b5ac7f1a99a27aafc58fb0e5cad687b44c2541ab756903776d29bb74866874263f7d4f8a2d1e9944bcc2c11e50b4e5e2ddb075a60644cb653d5ffdbbb97fe563e3088e5c00143f1f431c18120c55ccb1a8b7a9f315d0be964dcbc2675752624a34d7304cab9ed19107717dbb0c8a3513b4eab04c9944c36a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h825b80e4a3ea4326cb26292d91fdc88fcff92373bd5f130fcb6de1d7a32fb8d4e2e52d7006cd7eb619cdbe8f80809d79ffa49b8c8f8135ccb7a4518fc1a472d33348cd4b3c5674bc51982d11264f1050cbecd5e6b4917ea3e09f86c68a7b812dd85d1f214f2dfbb72a61dd8f192db40759ee2942ca5b6c4d0371eaf8b10607c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h158a4192e4880533e333cbff8ff440aebc9b94db14e2cfc0b6803776fee8b97be78827ba135f5fd8ee7219da89d90593cd5939f42f22bf3469a6e462af7d62de538418eb572976b8f426c8f7fb272b76b22ebc3fb4391db6cd8b904ee2fa3aa9dccf5e4f6025838bfaff8e2c6d64dca3ea824482d3a5d7bb14093e3d1bcee46e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47dcd0918e893a77bc6c7db7f75197f2b34987908c716dbd152905c07351b35524c1c54bc99c7e34a40de0e1e0d07c5fdbb5db1494f2c43449d5dc17f2bf13984981915a553c15932c68962780a58c8ec18708f3ae94213458cb7267ed76367c04f044652f9da5f533e94a80b858d467b7625582e87616e49befd0a1f9c1499f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h636ab0ba153c4aa8fac2eebccd724bf30198d409db9db278a308aa9b46242531c86a705cd4752f738f06dc1d59e8a7c7e8186b37602edd66bd7301a4a53c1a5ac2b460358d4443798597967d6c56448c9c5f3ffd2cc5682e054388867ccc834ca6f75642b2405a29f1766eec4db975a581d0a68128a0c42a8982541f1a9d5168;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40e7e2f6aa15fc206651d006071a3cb4deb2d29ee3e812814932a688b004c4f51582f2152012f46bb8ea277cc7a4e8e442cb5c088c37df39d2472822978a28471e216b7e6d56dc41c5e731d70273e126e2a3b247715d23f127303f5f6d154005bcd29f4ac505b08fac34df4e8a124965a406629ab31e559c5bfb7313fa7d02dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b05fcb5c399dbfe8d12ea7b1cc78b18348ac4829d8658b0923af8d34d8b7ef5cb788633fe6b99610b666fd2d8d8cc0d1e70c1be2f4982a116b69ded112879aa79c838de356b4259418cf69e9fc7ff282fba8f5619e1e05b60187d77fec690efd616cff49f058c5ce0c56e0e59bdfc6bcb2c5aca259e9448b9ae12f90f81d778;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c99c57531eff97b3caca08a9f3e55893ada1cf9c13f114ca378616fb361cf51b6a14c5c0b37f3dea63b780a2d96e2b0596ce405f1e6f024767fa65c56e4e87c034073296e9810ac7d415764582e18994d317200cdd11bf88ac78c6e9cdad9f5c944cdf6e4cfe9fdf4ef173e2d4e53bd143d016efbfcd038089a0e9ee1464e22;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee43f6497693a610ca4c55bcdb0cdcff92e0a9e28f7a8e127acb94d17c52cdd2e08b7ca862bee8eacdb3858d8e768b8c6f097106b1e38a1c0c5fdf02dfaa9a7a5b97a747b696b60ff58735101235d1e8cc47b18892bfabe721378bf7576cbdf1e00c896e97ac3c7fb192a8bad97c880b437f0173f4f5c4b3804a4d01de1ce2e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbfdd6de0b9569c733d30c8ce099b7c2a3cf9792f389e6b29f849ad872f5a4519f03be4bc7c8909979ca346d3611d7e4b1c4c8565e1a097c32513008cb59e833b922a5ca1ca080bb3f453173f419006eb61e12c7d9cf05b2ddfa627d05adceffff60bfb3063d69c778ea4aae905ba587987dc567397703155f8c9a4c0bae3e8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c3888b9eccc1bbb687ca736b773f20cb79f6ef36ea1fbe054c8690e51ec3cdb2aea1f09a56a5ffe0cf56c1d962f7820f2ae868913d13e29484b95087408a14dec544da29a6b870432e6e3d99b1a74005d9df66be74275161b3d882144bf8f468f866b2af16f32dd646c632af87b90ba0880089c60ac429440635486f49e6277;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6b5584f0a384824cdc88ed3820ec9efcb18bfed0c3c24f3936e85c48e9e7d9322c2d26316c5b91a7e1ad28959dd832c72379310656e587281b6679192613dcb78d9242f8a507f9745dc234cd1f379ab768d45a616e33527fa967f398f3ba645f6bc00628d3f8c24c62fb5e5d69851107fd38f48b020c7718c414bd4156d3c17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6ac874e110f75feab9763459f7c1a2e386544c568a741db33a5503913767347880302e8c8a8887a4608cf3419dbc05b88eb6a7c4083f2b5b5ad617d3abcfb766079693fb62cb6adbeeabea8cad3d46e46cb04f4345cf01ccbe576f1887ac2327247da7de534594bd2b34c5f68f1b6c6761c2f4b064fc8b1293c2915479bc02c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e8645f16e12831f3a8896a96fe052c0e4bf8ccc14988cfdfc0d314aad283f3d7ee45eb0e7842b2f8b572d229c3b55f9ce0d7c2bcb1e41c36b5ffa8fe759907baa5de97fd2280797d53d8493f675edcbe73e28cec283b7e3714418ec847172fb7916e05ddb78788bef43c8a1ff0bb2d79d01ad2537eadf774e1ca20ce6ecfef1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36e3f3c65493bed5fb0b5a0dd6d48205084bbcc1f3624c3a3c2af2bb66b8b5ab5b45ce0d2054a3dc9551bca00175d800a5973dd30436a4a863750038c387ba41ab76ddd8dbf5c5e3ee8f239ad94a3e88eeced2661798b5dc6795f9e8da85bc690090e832af547a5fb1faf5742e93aae4bf44fba28b7720f74a039f2e18667dd2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28068b4e8fef3e5ed4689f78a5b46cf0f11d99b01ebf6182a6c2f5c98bf6586377251d78e8e9b3597dcd39e0dcedaf364e3db5922384a3d1c2a4139c5808358f8699459c4e4071fbf20749ca118966564cc0b70e0487d7c2ade72915a958234ffd35724159137db84591bee35d5356e5136b482405f09f52dd01a6754e9427f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5d6772ca7ead332f3200e063b5d1a110b406d9af6cf1a7055feff904a91d8a09964d75880ba604afd4110b4b1539ac363af6dbafcce75bb367a4e64c195349b8d190bf8c07ff7cfb1cabb3339d1b808826d40d11f338928219ca83f070dfb9ed1dbf52479a137beca41f6f8c758d2b04660796eafe4b5fc338fcd46dcb191a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0d966129d7f2df13396b110f5f9a42c82fc02243fc3ffbce258f320e8f39e09b5efca7433863de34e137e8870f1bbf15d54550297b57d18894bb7afb7c5fd2c300e12ac7a72ce1f327f124a94c45745d9fad010c56a25422e91a7477327b0956d9f2b3f5ce279e7b306ddcad3e55412a94d416cf2091640a493132b702d77aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdd2ae76517dbc498ee94138a7d7ae7300d05b2bcae807476a9af9b1ace3d057ecdfec7902da4afa863ecf2a090048e1f4f164c17e75be8ba760eacda04890665dbeeaa1907fbcd2a92c677926bfde106fd25a8fb25449f75b40010377106c0d49d22ca3775fd7dda7d261d9cb89b93119fd338673880673af498b1f0b6d12ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacd9be1c2b364841311f827efec7908610a28ae97e5fd451acff87cdcc8b07a53f6c60de7fcb4a9013a2c109c502c03e858f2ebdfb3e331a29fba5a58ecf73f22b20ba24c54aedcc308526a2c482c572c68ee5932065d3bd9c8a625e04b2eb466aa49fc1a834c77622e0d897122a0d7e87cc52f0c86ba74b5985eb50e5905acf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4c09e95c4527141b2c266426a0458360a639bc64f71dbc9efba91fd59940d2f0c8c27dd9dd76c8ac40b48d07d826c6c8f644c806497665787a647fee9e4286d6ae0c4bf20f6c45b5faf06a353f675cfaae22a31ca1e8875e0708b9d541fffc04a1fdf1f49327aa4ff95539a96de549a83dc3e2e27f90bdc7e5a28860d713a6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b5e2a21a3b6519c7d804c9a6955ec7cb55f5ac24a660ce44b6b3f44beb9b741174940ba1306cff621e3435b34ec4efef55e5e754ae3427e4c82b272b208d1dbba2e53c702a416ee14623ff1b99e93765532bf623e5aba4e02548a4ade4626670176f5c7e6c5b68849fe530cb0e233360b0c236949f6b7439ee7db9365cb9026;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cafae02820cbe017a60f52e2f37241496dc8c04c6ecc91bbe4c066802bd0ad011acab962deeb599b6a9f54cf38c0a60891dd0c6fc72725270e4c0178265ce73c93d5db7b549276e023ba2bfe1036fe1504b097c58f52d9b1f4f40386a772cf8028281642ece14b5c74f035b205b6affe8ed9816fd1d30cac1955dad8a787971;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e35e3daba63d32d25a778419f1d84e6f8f85ba1ff8c141b8f82fb9d3844305ab6ca9180592797d48ef3ecfc7f422c0f28065e35612a4fa396aa61522445e62b9b87f90e78f150060d7e42622342a711a535571601ce970fc9354976cb66dbf71030d78f863191e805ad738ab79178780202fa49ef3f0dd715e7aad307e122a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4bb779c16bd102573039e623b1856b4eb777fcf2bae2e6d22ddc690f28a66c962808ba37a9850400c5f4f2e65c239b54372376167eda24e71bc9925ca585295724c7f9bbde12517a7425a039a6ac3f5cb630f8e3001c2be6d02e3411a05ad1332276cefdcc88dd1f9889cc9d87a0fa277f1027df8d761586bef553cbc9e7f319;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf79ef404430f1ca0d4164dd7bd2a5fd650a3da64f683ccfb154a6350cc1751577bc09b67273a065cfddd9bcad2f1bc05a9b4f1f8d41a9af39b0c9de04fcde12c62359864798b739ba5e47adba69c64555a361f1dafb3b5b49f59fa5f4dcbb9d43b02945bac6a9b0d971b2e2066231c4602e53008522202b5708f18ec33c47dde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba007fd145cbe29da11a99051cc2ef648378c9a7e6fe10f6bd24f50f74d952e37851231e1aa754496ed4070b2390ac2f07968c371f4991f0b310f7bec2c0f599c00dfd52156001ae1196dcf4dea4c017e2a0e7c0faf288e220d9a716f2887e9b8a6403bbfc29f1ebd8bd2bbe73b4e19d1737fc2b8650b62dc5b90978cea00ef6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6286014dccf19d15effc9e31bea0b197e60fb19d574054d9176b5158c7e10885ebe44065c1b65a51bc9fe964239a347e6c892e84a4be0d2069a1b677f20c9941e3083778eac7abff6f5ba824bebb37da2a4897e20d158598469fdf4a8227938741feecde39d4223510a39e4fdb68f52b441ccc6e3f37b4f5bf9d66e69e6aa2fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1509f96d257af0f98d86018e50e5eca82c2b0e0891462baf391e7d80295d97cbc46da2b2390142950d721ab34ff75fa214b56642ad0aae903bea5fd10b734f0b77942aea31dc87dadbd513dbab45c2c8ecb25b802a0a583280911fe0897d308dacba35d75cc05ef0607ac9eea5010aa0ef4aa9f1227bed2966dde9be1340d46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67818cd41dd6f596e56157dfa50164bd4d2fe3ce070a46035094aadf97450927e675a6be83b25e4b924aefc531f81afdeff98847092c348c8457eb37c28fef6266a2eead0c0378414cd8281d88652f32833d4d8e6f5f0c48fe7a75e11e558c5cc534cd905093e065d84ecc7b3a2e092a9228fcc0d459d28988c280f34456fb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4dfc3dc7f0fb991d5654ec609203d1f0d6324fac8ab419704df7b27aff4c11c05ad05fc29bcee13a61c73ab7f3f8f18ac4e927247b27ce78bca7baa2fafd77aac56d865c58abd4bbc39cf2c5344e9bd2167d4d6bec1c1c8492e648cefa8e2062e7a844b7a4f8140cb4f14231ceb691fa269c280ef61c091857789ac0393da01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h455deec1d8232e5745f7e8ad393cf48efc1c93d9b954e585462bdddb230a77ea298dc4743af6d8835498213a027ae05b35b647394e069a6adebbbc84a5adb02509b2a7f476b877bd6789270ab6da0847382f8292449f524937602ee662a4ef14c05321ec1502779b016fbec475bd9a2ecd172cd955185243916f7c73c7d61b43;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h490bbf4eb51f12518389154ed3c0ae8421dd667d960537a05699e998910889bfe189bf0574cfa3cb838c6be45cd333fa347622e975d359f83c352ffb51c27aad714070db5de4070723797605ee642409620e94e4559e7fd01bff191195f8830b07dfa4ce6327b532e69b1e29a639c71cf5e851798eeb8dbd637b625ef237a710;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b3a25c61a4a8d02fe586ae56f94d4055f16ded8de8554dac066eee35f063ff3c44cca249fc30aeb525450258981983245552a4317bf661b0da8ac2116cb630241720575ecde7502abe0a37052434972c56b5c738b1ffa93a7d2315e446d39cf357207692c69aefe597e81f6f8678f2a13bdc1dd31bafce24ab1b5667b34a204;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h630a211fb3e94a86361b6a365d9cde6019e6820479b1aa22cbafbddd3bce9300fbefcefd53a190cb92c7107b79c4d81a9d279bffd933b68e1a1f8d1c9d28b0d42bacdb0b858d12f9efdbd2afb44d12aab76425a1121b4c15c66ac5ad4883b71848e7a65fe7b04caa2645f8e3d543688ca491c19b0cf8ee26bab4794d4407a0c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6957888da5fc9521a205f43ead6705527b97af0152ed157eb474078d421e9579b27a6b9304d8cfb361b37572f9e0a873471b039de6e0cbb1a00700cda1e198b63e9056b3b82d0c5bf38aa527c2d882c5bb3f7457aa86aa7b6ce7eb309a0e1daeed38b4d114ba884c43c149fdf6b2f1735cb52be3dadff259968c2e6ade2fb16a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haedb7f90041f18ec87b3bc6361dd08cf1f1a0032a02964336d95b6194e53b61f73572e99d76da23e489775d79ee662bb93f75841d928746facd69eda6ddb7c8f1b5fcc78c8a4079862dbcf517d1d46b64e72f644cea113c9e9844b78deda4de24203922ed449067a46b423a41dba3a4c4bc80a6dbb88102fbf6d170a8106da69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d2b1f72bdbbfd81bf7acd9713fc5b49e469b304d6a316091541a24d0443dd387c04ca634ebfc194ee0717b43590a7100c70d223f635639762677f02f26cd357f9f321b458cb515128c28e06f9b91f449b0d28c05ac030c06cf62bf5340140ee09d0a36e728ac280aee78564883d2be9eeb6c809313357bc894225bc22b9633c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24657acf50e8f7b27785993ca0f41f222dc186120cff2913b6c74d36973942dbf20d6be41d07240542335c10f405522132482778689cb71761c01313c9a4cb04cd27d637024c2b5f157eeda5c021049600fa119a7ebf3f8f727251b16ae44df8d57c23a76490cc675399b4d340a94735616fd05af86850413ef9ea99dbbf4d70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h113ce4c8bbde0519bb251a8d2203a119e162ec35428fd1ced4f2520d3ed748c1e687f6b48aa3c04229defb9fde616c54b8c2633ceea0babc7326a8afbb1babb3a0af4f298841088450f4655b8476f436d1ddf35a64c47dfc0682c705032c586237a45a77201dc1b87c2e04e90754362b5f275c0e9192fb50ed5f72cf2a23604b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfad322b06f6295ee5c697ceb39377ee9102d27c36355a7fcabf667306b2404428db87f12fe7b80d8afe84fba07520ab685b7c631e23d5331734af55d00c2a9de64e654ca118f5d01b556859b1443dd5796f29dc7eea31b97be2dc53b7337f39a51ebe600ea481677361d7375187f427d7e9f7a43b2035749c6ddc1366abc3fdb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfde355d9a4ac6b702686fe24a54f390b8e0bcb590b41b82b0d89d43bdb10ddd36a812ccbc9cfaed16ff92bb696626e87e608a7a0a8f98cf4c2cfda971b472423dd1a3a98310a3e051b53afc214fa0a2e903f7817c3dd169c4634d1ddb71ad70fe1e1a5fc013e21da4b87293ea431a59ef761480ef59db4f26144302386137dc9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a594dad03c03f44fe2cce25f589e29ff337cf095f624e71b0745141cc31655336e5a79140c54c7fbc44bc41d3a8dc82a5b44fe4e97d9775d8ac38c2151be437a52702950e709b424f7a68376f972f50dbf1669459c50cf9e3f05c225a8bb73941589a22891817509894e0529a2b10e3907717a9eced9544890a3bb36971582f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18f9b65f110c02a672d20d7d2799e2b8ebd54a57e94984d7db1121c901f92569c441f33a6f37df9467e37e66b19c6020662e69067540452bf8374ca23cb65f24a70856f7106d425055416324dc453cb77e286cac9ccc5edb7913c7b0e81ae857df8404a02946573ac626342e887fbd0550f5a153724202d7f79171bd7bf00700;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb36f0bcc243383570843601bc6d1c1078dcd909683ad0aaec6f3ab8b100fed6379d2a2f5cf11de29a26cc0bdccd5610832e96f1d5b3be670a11f35383a993d3cc58a15e323f9537b5da7353b0e98b7c373924d1fedd55b11eb7d234969f0faa70f2005dc14c576d1f56b3f1c8d0a5ee83b22cfe451bb55d985bd01115fd920de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22ddfbc467fa0b8ba860002732462d9234c27dfc4e6e34102dbfbc52da91e66f131bcf3fafe87ec9053f3d850bbdf3ca68fb92f25d3689efaaa0d11db33911223e9a43b6830138355ded3eb59e965a7cbe535604673bd7f122abfcd382fd1f63253b0a74d9e1bec6e9d8331802d0fe8d6932eb62e6d065e7b8dbf502c0329fde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35fd332c78b3aa7725dc1906a6d3208fd7b5706552a426351bd42e2b329aadb24d3268491cc68c303fae028a488c86f3ea67242f0fd456ccaf13973dd6e16f1d82b48d74e435ff6989078806caa40e773e3662a03ca55d294d5e16bfa2176995a60d81bb1b26070f8a9f519a5b6edf245e7f004f390f7fa7aff3d06716695402;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cccfb7cfaba77dad151e706cccd2302ec63eb4fea561d5f1025cc02c5f067bdd02e24e1130033142f9ef34f758911138ae942db8cecc0224243712c7a90c7800f084528cf36400f358ecb4675e828f228cc194a4da8f06e263adc0e8af99f276eb1603716b48b5bbbfd0b2072f514654e426343049ba31741f84a60168c120;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h135693c676a8a687676e03b5f7189d0e6a6fed49803c00ce6329f4209bd271918dbbfda8e0a280625b3f6ea3452a3573031521f6580b5909f5fa9a285733c74298c43f52d5ce051931966adb7e2491039ade115cf007e77d8df5283db2d3f5f0ade45bed6535da6c0f30433659fd56fc43a54d59c2539d03356eb6ed6d169261;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7940d25c7b750127da95fb19d9a4d9ce1030ef70774f864ca9849f44eafeb443644f34c7d8598045bef6d1401901eca3050abaf9e01b154981d24b1cb65a55727528c6d13fcc309c1432b04beb600cb413ec8f45ff73d5f67a49a1748d6afdb9555e257e9f02dfb44e58909f3782b6dbada21a002672b5542c0d2156608c7e8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf80d44ed4ca4c5cc03edf61852236502ff6cda6677af8fc9834e9ad9fb7245702a65e70c2ef68ce18d486e2e98f216967a3394688758254650ef8fc71df7e0625904c20f3e3de33b53f199e6f1b7eeb10a56d22984e6ac53dd1686290d983a22322a058ed49c26a5ed10a05369a777b4633cb4d9be0c4a4923f38522ce76b2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48aeac85bfe669dd7191705411ab60ea728bb03bc69786db5a6f0831862732699d1a565aa707377d4a57e78821456e78b219aa1af60419d1da28ff1208250b2ffbcc90f481ff5572d27a6f86de56422829fdd18a0ec840ab91288b9536a43c6aa172e78fe88df8797f3b0fe9c9f24a1778d946a59f1aac3725e01e0e585cc61a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3a5acff66dfba7addf91309ef88f8d0dca69f45c321471d64cdfc247265614315fce38123f72ae1421b437875eefdb5d5469cd0e8c27aa9fe098ed7a816dd5d854770759faec99c6a773db3d8f5eb93e9e1013649863539a018e0df367a99ac0b0cc9ea96805275ab599575edb30678190db1c24588b0c43b59b1f2a1b96476;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83f0fc2a3cbb28fe75e7949298e6bedf4594fc84bc39c164ad16706953dd30ade7209f390eefd2358a39d74367840db922ceafa9644f0c66e5411e073978869858c28da6996e510d15aaf5671f5dea004932eaf92022a16734514f9db61a0d5038418ddd81f54ce9f30fdb0261a9fa36248df8c01426125f5d074a4ed08b932e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4dcbef5707f9084d2b311594c2268e19f71c57016fdcbd44ac7570eb67f756a6d0cb513fc1d92be02aa7291926bce8deb1e66c2acfea8bcc58070717b04dc93635a64a2ee290e81bad75247a36803f09b4a9dce84d3870964538461ba2aeee6b9e17b736bbd8e8fd879883ab8d46850b2548ba0c7721673921e8cd1339177;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9001594f2e971c750b36b15f4e93bf06ccc53d62709be0bb870d3e9560050d02df3f21ec55a224a547e3e27840d4b1aaa79058298034243571a9d488522c33f2d8ba0a4accb0ff423783239548a3400c7a98dede130a1c37b6dc06aa5bceae93fc0a03801ac3f097c7e8cc2af97abc220efc1e297c7265ba5d07cb9a19d0659;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1315e4a02831f1eb67642ec1f8ecd6c56a436cb024a8512231ad8f51af0c4ef198e2047806f661dbb1d1cf3cf99c102b958a332838651ca617041ee337ba7b165527fb40a6bef4469c4b3532640d67743f4d03810b7ed1fc5c82324bfe3ff4f6238b74d0bc1870e0374668c4864299376972c673aa7d4005f53b7b8f439cc7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae62a7efe4ff49c32aeadee13e8fe42ddae941ba8d19185000c4d3239c9a6beb1d64a96f1c8cecd1ec48981ff5b44ef67213170d5de3d138aa4a9ef59ad08e768359d84ebfa120b12a0ddc7f9e60051e0bc26a3e8becc8956c016fe739d195395f5e2aba836bd4d17b6d91fca55e35699a069bcf8075aa7fdcea6fa9c6f12ced;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2413fa9c730af9792d015d71d69e8e78cd62cbe648534707ad3a4f38d0fc43a30cf947624a90067e9c6802d318516aa658471e5caed83b835b4b8c267351c796097937ca892106e9874d83969505b53cb1a169bdb792e3e2231bf9e8c09d9373fa99c65a1a6b5cda2b8c5bf21502c1f275c1bf9e551ea4e9b099b93df42c66e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he07f5e677a65d098fca4553d7175cf77503af5f779ae98665455763a2371b7b1881d1a3dcc12bc3978b1d3d36b25a771616363e19eb2d2660f8122429999fa2c2ce8d9d2b7167d838933200d0b151c6bc31692121645ded122df8d0e585441b303cf378b43f39ea038c53e45cac6c9d7ce1b407f7887cfa194422196105af99f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46044da85458e747bb2464cc9984211cb140bee5cb8e17f016437e30ff3ff9584d86fc1e48bcc7931fc743a86a51497d41d7f0bc2d65a1ec9a3f84b49d8a151ef432220540a9272f49e4debdfe67b8f75afcdafca2916d06db60ef7a79ce6eeb8d7987b7cda39eaaca8ce3214c971bb8abf21a452c1e91a645830956c49f23da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf29cffe82d8ac990bd6320b1f84b10af5f48cf405d2dec626159b2e1a9b5e14b7b8fa9954095e6c6dde6bb00049a9aeda6149d2f6f082f458694d674f578faacb456ad27735e65059e5abe3b1bb0dbb96df209976b3e35dcb53e3a451e56599c7641f9d3c4e2736ea8a03b000e587d36c1247082c44b2f44a00e1e2734ea034;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39fb78f1eff3fbb11edb2ef09109444075c2c8978dbded293b953e4279c83b3e6478e4c2f83ada585503ed7ceb91d78020aed8618019733986f5fb8f73593f42a6ddacf641fd52a13b40d731740bdc34125ff781c944373521f2a4ca6ae6a0faf6bef579a2fb0e862c318e52d5fd789f920e15645de71cadda7a90d18f6cdc6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h741dfe32712f5af6e0d0ec2740cfea17711644897bdb10852243e01ddbfd6be76988da6c97db1b97c1b4da4a2f1070ff2dae128a6a798821c231ab3a6ceb4bfc514e8933c8ae41642e2cc6ce935b855ea085826c24741e0c8266eb18f736758f9c6ddf84855db184418a0e7acdd0a6625f61a58d05f6ecabe09874638d3537b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdad9d76b92d53c4c1a325f3c63f39cb29869471fecad06ffba4335dfc3bf463b321cd55be15158f4f1c243dcd57e181a024444d40343b0194688f06fb4304ca6b09499e337313654ab5b6ebeebba5066fd7cc0ec9b4328085dc8f148861ab12edf789156743bd9d8887098ffcb23825e1c4cfcf72ceebab60516c30155126142;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h298bfa582e474b113f57f30a61cd4661126e800431388c9e68cb95d7f71380e3474076127c9cbc2f72460ec8ee7e5871274623e2b10f903a0358f2861a12ea12ed026b05c0c319e767f974c1fa67bec68b7e9081aa64de38c2e177bf5255e7655a53e5ecad6eefb2fc4df87873de38c36c77e01ae58aa3a384a331159f59ea88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc767e56602c72d1762ed1c43d288cee67fb356a3e224d13ebc34dd5d88f4f3b44469b9614d8a8aa3bbcaf3191da071a349fb213f92f89526fa0e790178f48e20fc9e11b401629b1a097fa4b5b0d2c6fe821c658934d9173f5652edd6e39dba5805959eb272b27def2e4be915fffef44a2fd2db8895af34b9faa9f38f74de6d72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e695095ef58bf0d0e37303356c4f68a836a7d03a1c63bacc6f359f822aff3683372998c534b0325f4ed7e83946f3640d06a548c03f31b94e25a8b6d4169659d2181ed366641c018053055cae94d68b9378cb9cb6dabf1f357c6c3a3aba6bccfc6697ef1a477c597e07834a7473264672c6fbea30a9868816d3243992765015b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30405aa6faf2a77dcee709a240b1450584e52bec8361c0287463474eb1af256e2bb3e4ab827f6da9efba276dd15858d54e3a2c36ec2a75412c512139fa52ad8a29ac61c32e75ce0f7eae0dd82860ba0b7d14a1cdba6d91ea648933f4a5d7123fedf30cb3098b9cbc80f21da711406231bdd4a92b6f79f44a0ce57098a92e871a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h797bb0c0234176477ff743b4d58790bd24078e2842e988b8cb5f4f8eca64677440138af921d1f6998dd8f9680107b98918ee94d4403649b17392d7ba47d0afe6a5e66f3eecca810ccf2d445f6434833bd3fe3e7ff093ec31665df2a82f6c19259ff6b1684a9dd9d0dd4c853003473316f1256864794f6b321205b17108aaeb14;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a9abf778ee5037b8cf96a94d4aa792bc5f4d2c2a72bddfc7bbe2546c5e9322d0ebadd9282831e270cbf04ebad3dddcdb4b6689e0135e24ce4ad4c488b5192926a2daca153e4a53ac5a35696cc906752e9fb01326d4fa278833a20db3dd8900a482229638f40f4bcaaaabced4eb055ababc21a9088cde63d15209dc91125a909;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd1d7b20ae73c30af6fe23d008c14f6e71fe85d59a5608806c4c095773c50b97c1701d058b3859a53c67c2ef9aecb9d5d92b7ee70e634c4ee981ba290ff30e864650d038c9d8b2844ed3834ec7ea4d3edf78dfc936680f5f3ffd3f677be08d6616d3270490807736076a006e7f091ca45cf390442c62926d4ea2a9c8befd7fb1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1f2b90e1f11c8695df3e65265c9e4f4e7ab78a6c866929b868583a42212ef0c76996cdf5d3c4258e6509c8f979391e0597a8b0392ed0bb82d0831ea6ae3a44d4154b9765c0c177e99aaeb688d97c0e8b8ba542f546265f0e28f514b6f5eba4ec03e92a59ffa398c420bd2d4a7f63379bc2064963bf076ed38ec0309924da8c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6876845526a553ac91f098f6664201265ef99dbcd6feca1f7f3900b609d0374202ef78b45c9e23e2f3f27b93f30652ae9a96729f8a1df0c622aec848b06554019086671d058f62d9953a932721381735126c9a1dd24646c20b3ff7848e260378c6cd909aa17dc3c3579029094f753455e6f170c77dc9ed80a62e7067c8d985c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h779fc3dbeb66f7e4555c5c1bed5e430ab82e3432a5af602554b4426bd7e7805742b56fe69541c5f9317cebfd1e27bd55eff2192fa49a285febe2f27ae216e2a15b8cb915f3d2e7a939fde9e5e2491015c0b38d8ee33c822a733d702f6ff1a118f7a3214431de58f1dd4625f2ba595a5e48246bdfd1799835a4a004fc03c751a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2a80bffea33f1e2bb0d8c42b2e18c2263714f256ef1ef0197f81350cb5f181a5d26e05ff4a59f809b9a043435bdb77a7bf0c41d86251a8b2e36636f3fb9b0229be57d1edc192f25f8e7eacc459648f208784e762581759b8dbfc1e79d6eaf707dff00a8e36d87641f90f53d6c9e33eebc97444d3444949e2573139928c1c060;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e5ca35a9e0841db8029d3486b089f42b404d0efe24e07e6edf02f6308f4848e74969d2bf35e8836421f2fb17c2b147c9b5026d91301cae3a9326e7c9631b896ba0b1df23bc388e184b8879a57d7f3fb5b559d1c7ec96d7a5f9f64c91c0ddc8cd363955d86ac9b63232dc64d3d67c8875aea08a4403daec80bb2a183fe355064;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf99a083e6b7a3eb9741bdd4ac978b87eef8f1d96673e491a08ac7e4635fd11cbd33b7154c54d7e967de70ed225c5270a22dd0cc3b0e8da21f7f45d492cb843d7538cc22c2e59a9c33afb9bcc5764f5da95772c70eb5ecbb25c3c497cc311631b1f273e86230925407c1890492742b534c8cd9a2adddaf2718d7d1e017abd6b06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4deda60a67fb64cbf8f8ab22feb79426ece2c98214ba14327f4fa1c3dfaf5ef674fc28912e6848ff08385e2a6ae1677ea776363ca9771722729b38c6fa5aea71f4a880011c60d5a6b8d0ef629bdffc23b4e6fddab74a68d0bda3682daf42fdc95a3d6ca24a58dc5ab5df1c47d172084a4d341a77fdafdaf966f55077cd6b7a76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5886734607981a49480e23310e5087437962e7e267b16e5a1fb2058d8b97281f720a782651b191a36c0253e3b0733f4dc2ac4a97d1b232f3f1efb356ad3e3d7717dba2dba326686e964b08769c98a68bc4b68c389d50ac960fd9efefa8a3977d156948f1314faeb591eb058c34328317474a963d2af7c640a4985a74a28c4101;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h367b8e4567d9dbababaf097704924abb9d9585005802d0b80ca0e97652df9777903c30b7ed26f3a7511280869255564dd9eb0123536bebf1416608c45d6a12a4e0f75629b02ce62192bb77a63f678e29857dc1ba4be64980bd1392c66fcaca475b2b51a54d0b009664089a2f3acec78253a8d01ad2aa699dc01e512b30e11c6c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf72baa278c387fe8589fc37240381c76d9ae59fc4db64d617e70d967415263c8688ee08ed4f7f3f94b96fba7b039cf309068afe41d444ccd0755ae6876a0d9605194f3e30c607acd205f7eed359d3156a7cf2aaa84ccb6406179488c01ae2ca3bdd867cc8b03b5404412f078667e9c0dd67189f917ab8d57a1bd27916c069d55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc866f03ced4e8c951811896416d677328a6433faf6d662213f1771a3b5004875e23d3bda604acff69562fb35eada008b3e0fa6b00b08c610626f6d22b3d96c24ec6ede635ec584183d83ad3e05ad565a0fe0fe06f990e7ea4f8d0874270cd45b6a44360f2ae3bcaa558219f3390ce356f02508f5e32b3ab129175c95092c0a21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf605c0d673d0b5864edd06f70ead5e60af16700997e138bd548d197575b13ba40d452859cdcceeb0fc5761f284c3924652b51cd5728af85ac31d14bcca3c86b61c408e1cc6ee10225b4b3e5d8b68115b02f09d732293a78e79713a52c5fe881f762f2ca60c7332f88043b041bdac0c3ba03a8872407b25a97148ce9030492417;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d732746f65798878139f9358a061f4762f95a1570d5a5b75230534ef1aa3dff51d947b5f5e98b03b84ce14650c1517da4e32c354a6240741946a4de93358d17f176e5a3dad8eb9549d83fbf6b9cdd2340b09720aea809b75703b580153d343940aaed8fb47f7612edf64a0bca7622ed1d73ecafdf3037a1d9f041fa1511357e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he572009b08783724e10aed437d6c9bde9cbaefe7c961e2fc24aa77f30a79fa7461b8b27866d48520d775f5d3c168c1945aada4882f19c6201daeb45e9a79cb574fffbe9c7ffd584a1fdad0fa278c75276d4290481edc7676d3edf43c89576d1994359ddeec23a1926e91145a13112434268ef9cd982df40c416e23582df47d2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5ac5b7fd49a44924d6579c7b714ad07d3db720242a5d0a58853e65498898f241b057ff881131f56d0080a8393b58603de23228bad9e2fb01ff1a9bb54225e34b65750dd2545e5e1d6e41d3361f302a369c9674dafb0aea402320a7073cb93318ade814c4cb2cbf20bb122efe02c38f7e237d38bd48296db4a9fefdae2d6ca88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1aa28d5fe3dd9717f9d6fb29a8369c7106d2cc4d51e12b1f1be8462b55aee78798b234bca53f85533625fdcc2489e7cd772c768a464edb80016b0f618b3e385ee05e4e4077acc348e34c9c9af2a5c65b7c4b50963ae58439701201f3893f6ec8a38b4ea49b1ad92df3abfd2ca58409850d084aa3b7ca962d8ff2485bfc968f26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde4211ee03da6dcc74b3144f69bb4b31eec9d00eb9e472e299b1dc05a49cfa55be11f0be1117ba6477bf6b8a905ac1566eac50a2c06d36ea894628b29fc3c07494a1526a3813ebd1afc5f0a6768d00db7e2855082de10a150136f1e5685338676ba6b56f7e66b45e890bece21e8d900bc51d0e40df29072fcb2f9fcdfdcbf18e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he57798f6485191a6234a6879f548673692c4ef2299145dcbae23cf53361f0ebd35befdad86f384ce3558f861575156d8fe07de049c6fd6f0bee37055bd8f4ce02c4d8fbe3b8e86ec607f1e2a4a7e77711eb2c3f1845f4768df897a2f848a6728117377a3ca0f3cb65149b7e4b4d891624d487a2a3db5d925de010bd920d2f541;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bf74eac2c9fec000e8004a063539db297530b54c25d6661c97a2897e8b39687888d8e5798e4539778769cb4e29c14bf2d77939a7f0d4909eacb8b6ef695f63c3bcba303aa66ffc5326d4c0ce52d859f2b0b82b66a7d7e147b5226fca318de317f9a495326d307847806ec519a2b97eb75127f437528402cf6e7a3be8b23c9d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50f8360705c8c0f43fb9ccff5f028edab9d8405a90ac63722d0648db47bead7a52a38f6508b7c1356c76928e788e47c25c85e9b8dfb39b3f0b32f796c73f31985b5de5873732889dfe5216a25a4365fd7abd921849eea373b2e933427bc01119750881f6b76221f2ee08d76818d32e8b6b6c53db4964b35e4ebb0ace7e2c9be9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20baef57eb71a485aeb6b432dd639d20606cd59fa8c8976968dd2efe634adcc4a3877e4d0b1f8b24594c6e3983f6bc5c3f5a0f5b20d419eb11f570d907fa47332dbc3c5106936be8b308c518fa8dec4bfe48bb0820ba8b2be88a5b03cfe6924749bc9f113d250972bc2a9736762360d3c2c77d0b4263fbdb695319d7dd5b60eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e8e4d7e47345b427b9bdec1514311110a95f0ca3601cd721fb0f73ac6b804a9cc57845a75b30fea55c477827a6758299fbdfb452d334942fbc60c651630956659ef143820f7e9a00016da264343d33e91ae64f08f1778d2a6b9693f2e2ea9ce5bc3d02b24818e58f4a0b0c56f5198e52422982c4b2c0571bef83c7a70f06119;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h144d1c5864d356d44c60a9ef9004a34a8ec2a01170e1b09adfcf166a12e279b172456379da37b359ad335147efa9be21503833098c7a19252fda69c62e2b9a708043d84affe2d8a75e95a74a7ebd2e0d105eddb72a079f5af9723b3c2937ae35c7c95935a4a8733712c451459c920ed9080712a13bb5b3a8f3dfe7b629f8dcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0899832bd4772917645884fc313d17d6bbaeb480bbbd75b390c067b0252a3e533dcaa8ffa9d044ff49b710682bdca217c3568f11518fe7990ff1abb6b128a0688c57c537b3609d7d3f9bcb2659a60496b94fb9fd31633a74b826fd54764e4d7bccde183f53dbc78685850e0197c966c1fdadb8c17e102b7ed28064adf7f558;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70638c89ee04c68e67bb3b364f9e6ba54c9ae2fe25f59690483fa3fdd7166a2339833a8d2f39d7671cd04a692a2bea61190e9aacc3fd32af47d8dd792434e16f83d478f55c95a12700515432cbdeede2780fe7f11440ab44ee2c36de8fb3e5359ebb695c53e5c1a150a779cbf901792f462a251197f3b9a9df5acaec1a7af14b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71cfbe11e82dc66f50d057bfbb93bde093747d4258ef279da1c657ee371de33316ae54b9bc07b07c461a9bfd0d3059b7214ddfebb9c464d2df4f79ba6db8db93365e774e98b6829975bd877b2b4210ec24c2ac2ec6c90fa7afbe59b373b62f69985c78fbd1beb4a86e7a73250a9187e7ecfa81f85492725c08b8b0ca3605d975;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cb5061ac89aac0f9f81a374bc2380b8b3eb7cb9c8adfc9bd21a9977d869e523d546ee1eb4f465c27b53736267268672942654476c9682f98cc9eed7a55503b5bb073ce1f825887750a7566e0b336afaffb8d85f3a774790d9cbec29a6e61385721d3dc1769a206e31619d8c2794526ed19af70bc995dbc79dd731d0480eef3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6127181bd0851b9ec46d7b9efe49ca913c60a805df794b4102030d5c0dc1dc2fc64c949f8a763d63b96052df73ea948e3a709914494658732bb48226004167410e087eb813d198a76962e39de26c5d355c8122273c0181d0fbd1e36beef154d883375408dbf1a747fb6523bf47b415091057a7a4f220e60ef5cbd728011150d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda15bc8e39eaeaf363e7d11f5c7ef10b98cb60278cefa3cac0a3c1466d3bc79299e3a1914e83288defd2d5225b03b4d15bc69b2d93d6e72c73412cf50d4dbc395b9ed4431b1d172c350dd44949b74e9419ea6ac549a10eb5517f14fe59530220c4c2d17743cd574e0d37a179a73aaf82569c28c23af142f9a5b7451ebcaa694d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he98efd7fc01c8b75b32b74955733e04c8722558bc3b4e47c04d240d1d5e467814476ddfd0fa28fcb4ecd86582c226334272543d4874ca3bba97a3453448ed2d32f6c03a1dd1aa10ff0b4d7c247a27835cd3691778dff5fd20613c6294b43628b7d5bd1f3a4952910f7872ce178a0973ca90b60728c022a96bff5aaa1d8b05a83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60ab7c0571b6db1a574ed528c22b59e4afb59a6f9e99c05522fec9ae2c22f76e4ac07542ae0adcd5afc675e24dd85a9de7abfb4f0a6e21659db807d95cfcba9c59fbcbc772143b3b9d04c0a1c8c5860508fbd8931dca99fc278b58d0a580d9437a18b1ce91447dc1a6a3debe1193d47b488af8311bc8de793c1ad86c39352bdb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bdc6cc4a973c4d8cca7b637f932f8df884a8cb56534e3fa623abf6117dac2fb9486dac0e50b75517d19006472144a5824419ddff823f4f85a382f8c6b03e2799f839a044aa8a9a960d073bc8e1ca3130a7f11c9aec643a11badd06e0c49b51050cf5386d61fbba0a40355141e48e43bd2e7044e1f2311d89267233c462a5eb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfd392b0e37f8298e120eacbffc010b16738a3b29a4e0346ab01fc38d0e0b13c74063506ad1745b9ead7d898763434e7f78327f39c3d357b04acb568e3204ee98301bea2aaa221d975ea45cafed73fc377494adb37455160e32de52fc3473f0c9f25153856af0ff4f5be66a28de62a8a627a7bc73bd8c00a6a8cd0348c812e75;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef8d0e782a2bd38654d720a786e3a20373b7519ad0cde4fb4c95985794bffbed778ed539d1731e58fea98e4b5ab1b763243076b5bb65344823d0761ffa992f5430955bb40fe1e5085024bcae535e9d01562f1cd194d8bfe9b6adc794be3a6d25fe00f135f2ee646a6c154ac9d7d7af7938a4895e65231a7cf60fc53863496ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6abdbe59fb9e0bf792766139a8a937abc9ea64b88b3e9c62410d691608e61155d8dc5e8d58eb29d6fd3969a60017eb40bded4b5bea2aa165409834b00556b645b528004f6353b5089ddb880e8930f54d32adc1070d958f0b6edb077f8ffdc2e1a7115f1e8029127f60282993caa155839706763cc9212da32b77aa6f937aba83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h418b925dd0971f1fb7b378be556298613637ec7af16a30f39335697a85653e08ab9158a0195997433498508b3e4d7c7312e86e1e38cd091859b1cdeaac4fdd3f5e532b0c1ff1cf58aa58128733a8bc90317f2249c966505cf98a2d8a3588a44e808920942daf735db3ab13a114bb93e3a243cafbe8f9a5c4bbc98cc5342be8c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51beb3af36512b88e1083f1a70909a5d408c39ce48c5a720112572c8a88c9f2342359c3f2b8594bbd4bf103940f0da1e139eea2f3d44c69bad1cf6e99066544989ab13bd7e4c207672ab2905010cb18a46cc288540a334f976c868a0738847c3cdc74a72f253934d2e927d4f572cf4a49d07be92668c52a8344f81ed8b92c52c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cd99a1417c73ed1ff2f777b441c3135072131de50a334293ebf5eb36becf16ec93299f5c4c88e96233191adb6f4fa163a8cff4f139700717c1bd6cdd8b747a12c464324d6228d7d964efb7ce1fe79d153e48ae7855f8c0dd4549edc506fefd51a9ad5351486ebd8c74e72fa5e497d53ba12756def20ca66f0c9b057b529f5cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8786fbbbd867cd39fecafb0f8ac458eec6d69e9a932ef502202671f122a16607590536dcb680a890b665d93bd9b39eff50211bc8f51463cbda65a4f055b3fe1bf925c186187ff597ef797376596c963f10012aa67b80338a3e7b1496ca672df2fdd4d208f560acef19e11ba8a18590f8445581c437fdf1f48634d06b4917b96;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e6b7a386997cd25f7fe2de6e2bc1672eac7b8c94561f0381124d802d72f67c3a22ca1e1abf0fa59c74ae47c7c30191c1efae43d9cc0760d4e800234f40e3a11b970ca32cb3b255c3e29d013320a732339d03bccfef13c4dbc4d7915f2c15f56dcd2a705d0d90f4e4e4ba5cdab9047170c2f9bc3ade9611c7c63e601eb418938;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d5b9fb835a8427df08168f247e5a105c44d4b74df4de192e9f536ead2a4312e8a8337237c9dd1e95e79a21335126763d3944c55bfd16e85b6bf82153f5f6949e597b7998703babd02d737ee791fc9beac2af6d8392fe5e12a8c3a5d072396bdbc6276cdf800febd46b55d71f9243691428581f953f5dc23839d653abf10d2b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h769e808c953c9a1f2851f0912d0f10abf2706614a2e3759f36a58c9441dff880b0c6310ed0c0e2e57391cebf30e4d95274bbf6a3e58e9d79339f0b8ef8604a7965d95bb0238324eb9bee9161aad828d2ce2cfaf883de89659905d0085c96e990df1282302d9f8ca1a8a71ecc58f858c388c951fe3b651b3f011e7431ffb69798;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd49df076f3ed7020c61671871122f0e4f395f3f7c259ef3453c567e1738978402d155f740bc26498e2b9cad79403f2d7e2daa9fadbc13e1096390597c2f76e2b2547f2ff329263a7d6327da34d5b82767d5a4f0ebffd963d9e084379658396273ff53b0f4e38b0e1f6a3ca380c8946a5cd924f948108d2a4c69e23601be06c1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc50b7ca6b17a2dbf4a99197c19e05aeba217f1c38f332a32b7005168182b2cdc6dbed3dd8bd10e625720fd9b0a713ed5ecac02d868cc6f2241050a09597c6a3cb0b585111a3db8b1e72362cb2c34870ebfc4657442d616cbf9e353421656a76cf889ef460bd37cd3e079bee61da5539490c9cf5fb5580eec391ba38389a77d72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb455ebc7ccdf02311b53e5b3501e69ae4932ee8bc8ff72b0251bb76db5ba26574d53717dfa46ef2740bf5d6d33b246ef2ac4f6a2b55be6f4245949b07c0d092408125a5333f7ef481daaab30e0f641f4784f8ab8d4fe4227e6979c8b91e3f1e5fd2afd9996cf8c33e3eaf8bc69f35de4135b48b6beafe8160ba41a1cdf55a874;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13409070e48d8cba5e37c96c33051d124d0b9866a49e84b59e3806660d9d8b41dddb7d89af127be60694c33dafbfad1b56afe87d354f703432ad05de56e3fcea5ab1ed61a5abb29d0d4509fe69cf7c7e12d583d482dea302718d61485387dd4e542ca2868509c900804281d8e4fd4bbc55c2e20468c23875f169de1b59ad7b1d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd5ee0bac25dbbb6e3b756833f03b375ae5b37a5458d6960a1790b76cc1a384a38f0b224d22561303886741f242956c51f2a476dac5742d5fcbfc13de114a986350010e32b133d67d5b0e5d1fe231e5ec7d013203e609090d24d13281cd7d79c45b84466d14d0abea012c5c061cb936ddeb9639d6565c21ef15b38b116719a32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5764f74da14cb6c4b125204db62ef93ed467052ab8b86419c51901bfca227cefc82059c85a788b287bc799a0ba624158d7ffe99bffdccf614c9b7a09dbba3f67278e2ee283ecb9c5940a8141283a3a6c2880ce778df83b1f432f9b8bb3bf7654c65c0c55dbd95fa793c07ecc22a04436e7597de3933a46e6eac396155e94a1a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h281db063b7f90d96cf0d41d72b2f503e79cbb2d3b293fec096cdfcfe1b2d321c9b7b8093a0a1992229b8645265dbca78def66563284a86772c086514e8b047053d4371ee164f556bfbea44b00187a6d7a1e24840823526ca332117dd0376cf6fcd5e06137a80ef9c6a65c1f3f826d45c92057fe0995c3e84dabdde49d7e0a997;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed09b7749f45936158d21ef34df458f2595919ab065f11554e19f794ea5b1b7b858a5e11b26cd9e2129a1ee593b301337405ff13d649b23546116fb77578358b74bb26c5635e929c9f5344ca24e2d2b28e23c810f70ddf563c0d3a64fb9863b0ebd818410724ac2a25fd631f20eb70b038d341b38078618d5cf20db0ca15a8a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e3f19748edc114168418d5d73f0288ccffd810af2aa57d2950c07a0da30d2ab188655082ebbb4261fc85e8d3fa56e74ccf8cfd721f0f33d1ca7cd151bad926abcf6b3240b6c29317d6d3893ead3d196f63456a378b8331cee660e7bde359cfbcba5adf1517072e915b8666809cc6c8ff7a778d79288abca41b83294d6b67d10;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf822ea21a2542aba2a1149198575474a33c73ba6dcf1d602fa16d186fb2b6f315ceb25936cdcf50db4f045ce5bb6389ec36a9f81b47e317a6bb3bed63110e024bc6ce5fd0af43e794319c53c9eb64e06493d432dac4c994158aee5ba09024b0f2b7438bfac89b488c930fe55a392be7bb5da6054226661b702c8900df02d6c09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0b493e446daa43c6058e356115ca11284fceea8fbcd38ee2e0123c63273c10ca87a53a3eea679737478d1cd6160762dfe9b13c48e8228a4487d1869316797ad425e3e6ace04dd1f3e8e1095ba7359cbe14c42a687d5fcff6289766b0e708dcf8185229cb63eb632747506c724a2e21db35ea899fbd66e2808b722cc00d69bbc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2d9a07cdf38ec23a34b439082b1fc457a2596ca530fc330f9c333c42ab593eae842007569c1dd65be5aa089fe8934debe680d17c854581759e6b6283ca4b11c26a5800f3c1642845f72cdb018dae743ab0e282bb846157fd29526d845eff5a51728bca9dbd50bde10a9fe64fb0e60a7f9cd15e55460014cfad4f43d200fd7a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a315122fef99b7495e762e855c5cd3628c41ef7a63b5fab4fea6c14040cfae4ea710e7cb32a16aef91dfc26658030b0a8b109dc4ab7b37721e28fcbcbdc4625a473ee0aa42a8b2e5b1fe35375821194776b53339b2a839e6efad0106d9d25d95b258c7536e164d76343a6edbb1ade029df1ab06e23ea1e5a7ff9211b460fc80;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ec37a1ae53ab189e14194d59e41d6f7d99ec5d717d3c86f670dc61fc352433c7bd273a6811fdb4b0681ecdc28d53cae33d0437fce21b7c8c649c21a76df2f80c563af0a8060bfa426dc5e4e3ce21e70bcfd3b0fcad21e774300bccd91a7c884cf3f33bfe04d97ef46b3cffa26044a19167fc2aa78e1237bba5d22edfdba4c60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha09c580b8bd6f6d9f179814cb4e8b4cd0cf05298c318320ccd511168502c88bf2dca24337a85433d17e538dcf7ca2007db19af5b881daaae6fc13d4294e497652dd04bb4c5c3f3e9071f942fbd28476d70f73bbf6ff51570d492a60a6b7cbd4d60f6dbfe4db7eea486619871ea06b2ae53ffdfd475b797eafdc96e8d15c32cfe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h861cdfc4edd5dfe70f761fc408acf4166833e585a5ff0c178a6d1a2bd7c162c91c258cb4b0ed565ebdaa0c17c8f5b56c81788c0631b8bf2c37c348c84acd6c121f33224be9778a01833715e659406ae696d761ce610cfc509804cc9f19f5db3dfef75f2b68eaf85139c309ad9e99bb5d6f041cdb02513e2c1e6dda9cdaa5d8b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h362e50f5b00fa87135fba1c08f3fd588039f76bf24bab692841eaf5ff96cecf807ea64bcdb505ca5c0c43b7468ecdbff78cfc8463fd6e064a760f114aa9d2e86500fee8eb7b160c2bb294cdfedbb51ec744bd4e56b8473863d8f6bcbe2fd2b7133f72b580fb7fd504060a1297673e7f9d7ba96af1a44c0620bce5185e882ccc7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf63b9df0dd1553b9ee844532d108a1b201e5a605f0bb9f5a3bdc1e4b7820c4b24241ef43298341526ae01bd1d8ac2e836c147b6c62ef393203516a1d3a792e8c750c165dd44a4eb9c3d0be657366bacd73d80608917fbacff6b782df2ba1dbbfced31536d55401bf6f4003f9258bd8e1c4e4e2def458860be12bc5e641833b02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb739bfbaa30f8a6d1933c62290b05b756be07406cf6011ac90fb8c8f2769f42a4e7b9884cdcf8958b629f93f7e3f9fc45ec97b8a43974b855372141889f6f8a7ba67428db9eff9881387b18a6b7fa9a95ff04740150167751dfcb3d1e30c88e85960a0161966fcde1752a0c017780c2ee1e8326bc6f8170fd48d21fadc0ef6a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80b41ab36d8e6a3d0d5dc0a6a917d7c556401e1af21c9c0e3aea18e21e5c22a1dffb50d595e626309ff8a017b48a711b05b6f0b6309fd99259f8990d5d03230acca18369f2930b9c0213e51ff64bf3b3a1556dddade2de6a63af991af320eb5b8a95420c0601e7b7af442d08571f5b7bcd9c4a0785a53487b0e5ed0bdb2d1399;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc86908269ec188ccf22f8c64ccd9fae9d89b1013eda84987695d79535d657c54541c1cff4641d5c1fb547aa7af7f39ab568836ea4e2c35d1f78147a8d21fff9a0b047607c58ecc5c4db54b0712744dd38c4df703cefd0f312889eee2e872e26304c4d70c06b31737c0125d7cc992c47bae5e8811e7af5cb93800848c2059ff17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d31e99a077e9d367fe7d3de25538a0a6846b6cb6ce79b1e068f28704458312b2a4f9429e8cb87de5c3310c2ed9f5b4eb7bb44136b3b5cfa0a5e4854b4acfa910e027a908414a0370ae0de0eb073dcb0b8acf4f5c4fee56fc1d2670a60bbd591a47c00ea2c3e982f9c3860da67217675e16211c51810ea388d3925c59e495be0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65cfcde1fe5e8f9bb019059836ef4be1c61c14253de14545ca86dd305512b908dcd30ad220c094e63025b7c3a6bae94f05093f26e68d4e4ff5e2fcee9411f7c056ef5b3e26dbdad35840db3b0054abd74381014e1b5b0576b94f755840e7691f5c5e1e2d7d09d74423cecb5c51a6c79c9c614d2bdef64a8997428dfe0cf7f486;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ff24395ca6c4e2beb2633f5fff17f7780e0c25149083dd4cf8c540ea398604ae347de75109fd4c7b1dcd59d496438a0ca2b595bc1e29de6f2bc062a8dee7bcb7f125b896514ed3f29a5e9e570a563ef3053a37b5d3e1de7dc78cd814d1ad7e5b9a0a9296a7e20b0c53aa2c8dda5d5696cdf5132af1d42eb00234292822b4610;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3205cdb16001caaa0544abb233d02388cdacc4f9e4d9683b3dbe4829b7eb2e8e13857068a14ec9112b7a6700ffac441cbcc37172709a60fcb1caff20b774c48a4d5fd4ae3664c1df25a09469449e43ccfc92f4dc4d716030fc1eafeab776a84a7f6e27fa07ed3621ee5f69470f2bfaa714f92b6c2e3c2d9876d6815037021148;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8080d1ceace16d27a661b703e1b9076a993f3f626a6ef0a071b2db325ce8b2d1285c34c26719df419755ef1a6b4cf7428cadb5e43f40af56fe4dfcad99d6c2c0db9cd5be07cd73d264707daeeff6a8f973b9c72df2049af17ea6918a98d50eb4c88dc63babed175ade653ae2d7cd04f7b3cf960897d3cf073eeb3d08e3b34318;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedf4d2a9d20f6e216298d60cc449512542ed71fd7a43fb6c62154612e6be4685c03fb034f084e8fade0538dc3d8a85eff0ac2cc471e0f915841b78408cd315bb6b5df2455f7fbe563c472b0c2f8416cc44fb02b596abdb7328549e0d5a61ee3d3e523998b1152b7bb2b2fae3a09abf56b14fd5433172659296ca9c777f451261;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7c0573a42fa4fb64e63337c0380476ee1086535bea133529390bf7ac5a2924004fa66eafe5954241246b9c938cbae9d9d3f7e2e36128e8531d7ae2ad143a5cac88145ffd00bf639a633c2644993813dbfc8a4682f8b915cf24c12c080cafeead2a3d08d4a2afb9391bd7a11b23b312b7cc564f33f6f6ca0912ef0f266dea862;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cf14e213565079142a885c1c1e5070ce903a9be3cb4adafa495ffd728925bc9ec9a49f73ee847c9087473b7b4c0f00581f84698ad8c2e7bdc0630de1abb2b4931383220cfd15015a4bf5e1c9d6e46c05683442e8fe20fca6b0aa854cbbf3a23868cf9180ca04f55011e30afc0f0bb26e76463109f9fb7297a3a74bec8a9f127;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55d819acb2f87a4a5fbff7db42ce95f13957a629094e5084b64eaaa1b85db29e3ee760092c97fbce2b0b1aabad15ad95fd817ce688fbb671b996f2ae2968ad4af993916a569e7ca6c729ffd95ada6421d033c11fb13ad8254d2b88bebc506d7977d73920d067594673f70c40db3425e993c272c455f76001c5212c3f93d14eb7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd481a0363169e9a2b3df41d543dc9af4c7430e7a2927ace7cac509fbe58c8768e4f8c7d283ef714c4e63e8b4f5d5db0c51d9cdb9e81fcd4376891d7a089b7d0c16fc1913eb7728a4a1269b692531298ec6ff791798cbb69152e0089b242d5dc7b22a7916a866e476988c03d068eaa825410ee33545d3e86e9b4eb7fbbf6b92d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a73c5c8ab781d794a91b3fdca364eded78b4e04ab145f66cdcf4d5ae7083fd8eb0974c35c251d09a3014db73e7ac17c9cee7f42a497e342d1b3a9f0ec284e0492a1b7a0401d73b0fd6bba6ea38d86c643555525385af7046c0a02a02b70e13af0adf8fc2868cc2ac65d7603ac77e578297c057978b0c00fb54ad5c5b980aeb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae0f81bbb83ad21e2ac60c79c12cbcd24dd288a02c748d9ae2db5c92acd17ea50dea3f9c5cdce8a295df1544782fdd899d97678edd40d181633cc400ab0d8fc63ae03b258674333ad4323798242529c548fc8a53321dff949462893703899151f8ad5bbba2f7ed5f28f8a0a4c717cc1a5f65877f1bc87a455abfdb1983be9f4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had52b1a74907f04ba618d180f958f7401a9cec893bdc7c5b9e7241ab3b8b4dcb49cec9cf905373de2a3c3925bea50135ebdef533df4f853805c45f6251e7e98f631ccd2c8d2387d70c73bb76d7f498c51f4f14e867d9a6ff284086522ce33977d7a2c1ba4068ce2d215d5566dc392e4774e6bcfb698a22614bdce2b4a26dd819;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d4964da49297e164e91e7ffa40e2c547d565bb7cd84871fbf42b3e73e3cc9353beb267e4e5dad7dca40070a6e6598e4ef5a93bae2dbf78281a113c1445abc4ec350421c3aa4f840c6ded9c3372f7438dc7e265bbceceeadeb4cc40f1b47acc9f7ad7b2663c854d8150c7882adc2a7c2064307bbb6e500d9feae5bab2f7e56e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3fda764d85b09ad1a76ed2c06c97c0498ee6c4fd2f502ffe9bb4cb72250c2141a27882856e06ac272d557590b84802c2887e3042fe34d8e150c1c10ca175752fad60bdf675df441f53f1777796aef419d42c27b07f3be11701d1a3e6ecb356b91b34c661ef51b5d70f60caa211e67940cf4e5fc15747b1afd672a9ee8724d72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h279206963618a8dd6afa360f4437cd92739243ae5b184e4634e681758bab21e1269306c3d8ab4a75da6d9805540b3bd7a0ff71c0b27a291540cd57ff57c3ebdf8fef2eb5b8a87ec3e4a4f0c6710770fd92ebf0dafc5bdad2567dda0d7c1e126b6f0ae8936f1c5923cf4da988d4a93bd025acf0de16993f5325fe1d91093a3cc6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ff94710d3e7b2055c86a2803c27404d2194602d47bb40c23fe0e87530c59f4f49d441ffb9182f0c146a27e091d77d5960ee6624c352318ba291a2f4e065ec58ccf8752e2679173d562455c5284447f74b9e6bb2a9870634d32dcc412be9bb065df8bcf44590ecb52eb6a5a2c8802dbdd5c59d935054d863eacb67f9eaa3c81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f473cd736b5675a89f61a4c7466f0234e7cd859f07e2b7de41fc1d17d03f9182591eeae28dc4ab13778a21f65b4f2b966a07d5b60e9c6ce23fc64497dbddb0b46a7e1604b84229902335eb91e2c02d6ba7c45997ef49eb31a8c79579dbd38ee4dcf159626ce7c643ba76fec2728896578d5366714345caa7ed469d82bf2f58;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8699ae9aa9faaa1a6b5f4909bf57d25d4daee0c4ad6dc38445b2660f7eb587c7d1f753cabcddeeb1746fe3819b57ce5253a48b3d5150da01032326c986af353da35d154fb062a0b9fb72525ec7a6fb5b0c900a1d51d76d7bf50ab1b2a693280f6b03bdc1182abd8b6a8b00811e54f40ad720404452bff37b979f6a1c63f46695;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha26bcc3a31e969dc3a0698aaa77a28eb4f718b31e0099b2d6ddf6f5b2789f141fe5408d5e2addcc7ca042bedda51e44d37242ece400781eb251e213da74ee4165610f963b83d1dc9ca11decd89923dc0cc728e625a240985bf8228ed52974188ac18391221a096a9a4174648d8667b9211e79fdbdeb1655d57447baa78dfc19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee7c7062de9a394cb6f30498eb1896497c02741a1c9cd7f2d499a71528005b270b342351d611acf861495fb8b57cf9bd8c2da12770fdf92848fbf7d7d83f635afe8e4f288f4ca0d930b187bd438ff398171401e6c96b863a0dca29a4e08eac1e5769c90514ddb60139b63182dc794cd0fcfbc755b6e0863dbd11ace424ec16a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5d04375e87dde223dfa375930e1a28c2e036c38f8a041cd1c331daedf9b0198a1537e5961463a7f6c041bdf2e37e6b8f7a3a3a70354d423cb7e767b97497c7ed1993918249da6be561eff09ebf2cfe872eaa8eb21b646892d95ac0ada97016da76d2c6691f8e975415bd3cb92ec643fad64cddda876cf7e75f92b2de8b891e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88251733f3ac5abdec6daab13a0c8210a1ca56178a5fc779354c75b48841eb86c50e1c5c76eb4f065d22b29e4b131360f9c8f2b4f6fcfb3d804c1a36d313127112599e6cf02d3f85a4657d3cd3fbaa33bea0f663f87ca8c25618f566e956aa2fd4f2bebacf1217d45ffd769e8c5b6af78b39e921ccd75619e10ffad73eb1c9c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fc726957758602dee1bd3fc66224a515b5ed143c81fbeeba3f9d9a84b158b89b358f7a28ba05cabe256a40ef508924374ea73174677a208245b71224a4d23ee5c24a30bfefa77e31dff2eed1abf072eedeedfa50ce51f44857c7aa30add97aedd09353046e3861f6edafeda5a23077325fed74340be6ac45c0f7fe085995aeb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb90cd4559450bacd20365cc49e43d895b315723d63e6eefaa3ec6081fe1a602c28ede36589ca8d12f77bfc2f9d7025a2f92e39f76636eab738338edbd458616fb4aaffc80382642f3ad3f921d42c233151dd208be928d5df1ea202100658fe54e1b1bdbefee443fcad34389ab496fd82dae4239e6d9c8e737ea0be62b3f460f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8de066fab94223c8fa50ba6514eb815217839eeabe6413fc71d55f1ec881ed65b125c275e542629da4b946b910ead0a88b9e67dcba428f2b34b240d20a0d6c8b9bfc8bc9dbd55fe7e1efc39da006506c65cf2126aa23ddc20d24727089e4d481ef4c5666458c917d0fb8f89286c00d751a2d270f522430aecf5d88c2a27a62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b855a2118b01995c537ffdf3c7afc98aaecef365e75ea534c202034b643bfd9418ed115b43af19b1341c1c5b49a480d77aec204288b18b17bb77e81b041af91e1a54b7a70bf6e7452bc23a001a256a3c2ba97029820953653277726f2ab448f2a4e29c905cf36f1a82556dfc99d2ca5ecd73f4bd4ed4b367ff90cb52c53cb27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefe9563916b0cc6a9ef6fec8854c01b4b1625bc04ce4d7d00ce522723324ba5a9b162f8d06e32f515fdf12cefbdf2c3dfd47257ea1465c1946df8ab22c185b6baf93905b53a379607d4aba5d59a9953a6e6782a09d7069510f580f52b02bbc9ee30becde5eb0388bb235421d9e37bdd686f41b07fc5d075e24783ff007054c12;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha23d4b86c854cf6da974e51c5f2f6d7bbe5b3bc44135d1857973bf89fd06c8462b47ed2987d19c254e9597b78385a2f55dd6f786281ed00b89c944d78960ad517de543f8374e459dd1ddc5b796c3bf729ce75238ea03019a918781515162feab5e9cdfbec110137b1ff786c33cd327dc5364c40cc3fa1ca1cf83d4c04fb3e9a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he31ba2178ff27d8accde2233357d66b20dfcb7eef1fe8f51cd1dcd9dc327f8e6a41a21d5280b48f7571b827c522f77f994ad666366d9ee6ee9fad05ca8952e59ab4ad5da814d33f731ed56fb7e5f71b52496c7f97a3df9dea245cfaf8bfe335e31ef688f1f4106e65b3398554a5f250795537bb92d49e377156c4e85f24e7ed4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2b4adcb2e77d8f747a4646ca0e055a212348387edeb144d538f7382bb837d513c402a8ac906948849391064b9d5bb7505699ab4209b2efbb9234dc279a59b5caa5c7f92e09ee7137d5b951f65389862c174e417115221d88a264adbb5de85fb989edb7ef75b082fcc6c3d784fbb629b2449d8c39ada4e8cc95f248ca5df5a4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbadf55c3ed554597ee8dc9f3d53a36ac59d944f0b3b5f90b799913c7ca2683adca01a1adbdd42f7592dc7d9d18cd62d555f2baa8c9b3a6d8bd14375cdfccd0acb721aa81e38f3d8dc8f7d39c110175431834545041397d4640972ac3039db67a17b5317f02d4d8bf491d0bc8d6727aa29f00ba268f858119cbc8831383ebd39;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4210b2667235101763336afeef2add1a7e03c85a107de723e0c0b64d014962c8f22f01489bf9bacdc4a26c969fa38f71e2eae44fd5b55489613fbc87e215fb33f70dde5f055df16e9adde9305155b8bdc24b4331cfabefae883cbeeb41df663982240a911fa5d0ab2ddd591ba4e0c1052e83b09532c7abee592c48afaffbdca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b2cc031def16d61362fb5fa55e960640748a2d2f2471eb716c52a6ab4d77896fa61205fe6c94b81a6902da097065479f86f53a5132474c65c7573a9ec3922c02cf41529b6f1a04bb9d743820a709d0ac5f963896691172f7511b84331187c47332617a0747b38761fa3dde67006c85f5598c7a8d111c477b450dded2684200b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ace07c927360d46283245a02994833f676b77ea3f927d31150e537b5362385f63a60848630e3d349baec965701747f520ca168a23782ef00ede9034c0e4bc5cae4bf942317707b90f9a0d6c66dcb6e9b30038f00cd4690c5ec56fbfd8853fb9d552e39fffb8f6bb6aef59a3997dcb886f1d4c1638aa96e67d6e309479e377d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed2e7aa0b29ce7259068e798a67fe0e0fe8f47da63e076092ff83958b6327e92c5811a7e7d2664837f1ab08bba649aa4e310c930697fbb4bd51c38ec5ceef36d0c7b01042fd55ced4b16c594087097bc62ec1740a831c275ce51e53e8639d8b0e4182e30e4eb0d5aa810156f499628db4be1732336a1c824a0b313c50b5ba3bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6aed52fe6b11a997f5f10285c7accc430e796a9920af68c75f55a140a6554fd63beac85dfad84cfa9155cfb85f2b4c10de81ae9351457b54f6ad6057efa12903156b0db5d0607acced54b28f0d10b6dd23ca6a96942c134b3c7e098d5712286caf7504c9dd80507a5c32191f12e270fe2e12ffbdeba2dfef8fc75d23a16f736c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he639eb35e670f1e342c5fef12e13bf151342ef5912fdb26656df3a2e488d2e076b39f8889f433c92f7a61eee3e764c648b6c0489d9512673d3d71698ca4684e5a45e3654eec2b3dccec8d832ecaf098049a2675d9865215ccf1a1cb54f6bb8b951b59c3a52fcfdb995f505ddd2fcc00df12ddf947efdaa3666611624985897e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e42745563911e62e3953d761da4cfc3b5d61351e9848daf036a8920773f44023cd51377fb08f469945d55120511008a640e525ccc5b60bece490116f81d7e33a7360fd868dae37057cb85e01a2554ea7296e5b9c32a7502c4c6c9583d811cc56d4b185a474644ee5b14ffe39b332bb26feaed3720ebce36d31bd09ec65c86e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h448970f198cd8c081301ec7f3010e274a246dc6c65abec5818535f8a43b1b04dd352c6f6d2c5a0bc65fa13b399561c76386406a18f82cc930861945d068bae87fabe5db1b4bc8744a779827773e54cfc7ebe1c595e0ca7f1eaad06826bfc6e6a1a7a4fa17d56ac2c5b9a809daae8b20fb894263072d32b6c710f4c61f72f8af7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b012c1fc48fa5ebc78aad8c2ea99450a6b00936dca978efefb556149ed62688dc5cd229f85755f842315ea49ba109b2ea4681e272bfbe0e26e40c60f3275ed1fbceafb8aca448f8889f947afc9f5dba6317b5872e6c0fc1048816c19009a5e802951d8738b662a2be12cfe422e34247e2fa83ba5aa66f29581fc95f851c3ec9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3861aae4a6be45586ea3551f4bab6311e439ce8e064189ef261a3565ef60d79be9dfdf324bb6f3d5d2d3b976b7ea5bc24439995b2b3c0cec6721db9f1cb68b803f9366975b74eb2e5ae7212873ae52861b8401f0cdec7e3233083c2993f88deb8d9dfb7c40f78497dd151135b3ceab270ecb69ae42a4c0bfbc71cbab8c82d6b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc448deb0f6a7cfafc905bc8d98c2fc2854e38643c548dee29ff4cc812e5a575e9ee14235943947f3eb40c8c1a554f2a818da53333b0dafc91f8b11234820d6fc187e4e93d1511d5332f441fb5145f303eff1c0534c13e149e35110cfc7976c75ebba91f3e2461be6fd0b803615426ece9e007c47f614d63105cb40fce24fb906;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7298d7240162785c6dbcba6213ecea8367b980a5b49642cf4f490957c07686502375757337b0ce082278d2b08352711d031fb50ba1111d4eed55198141bb1f3a02298c89bdf55f8bb22ba3f77326e9ec95c287759bdfa1a68a5b54518a704ed636cf1797738a780042d033986d934aca33a3e3dd039906381d264d17ee6fac23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb0bea98930dbe16271ff4438ab0d97ad3ee5edc95d380b72d3aeed83b4b7922debc435812f19b80dc31f72e1ec23ccfbe811592b3959eef5be95d020e1be543a9a0992ad2fc6d45c036490073f8a0515c4d085c2b0743e8a416b0d8eac18905e43f2eec816b043bafd0cfa66035f1a47ff6e9d04fccf7eea44c6fd4c65e03b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2cbeda74e62ac05d7a5debf0738d02a633c102457199af9d4fe1bb274826f1cd27ab824cde1ba1e2893a4ae9e172bf886ef0b6788c8333c82b2748eae0035e381ba1b150debf0b5e6d0bb168274f2fd38ef279f332323ca1e65689b0cbbd43f1254fd18d962082bdae9ca0920ba0d81541cf1bcd82eaf194a3b5ba5f6be35fcf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5032b5c91e39e6f0665e118b7a559ecf4c283f81296d47e0b7313d20552bf845ac0ecdd7662218e91bf9f8f473626f6864c8d738a0f7011d91ec699967839b2e0d204dd2adc795a448c69c5a528ea4eb39bd7f77c1e0b3910a7ba29e3070e980b5b0b90713fa213728d886370774b1a7437aefd5a3a282ec872b73a15ea47c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h368dd375d8aac6a88b568a1da2b9dc6050b907f4a64b9438e1fe91f58bc20c5b6cf67a40b14506eb2059ff391973b2ec79f1e6c1877411ffb84afec3346ca7e888f0b693971e52a567c907359146310a470913acb785de1fbae025d0b49029640d4ec2a42c81da961f5cf9a9062d5010976ff70e57ddc7a822c4c6e506fd0c8a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h872c27f4d55e232e543ca50bd9a36bc9f086a97f96c2fd10fa08f3e9a8b8d9d4cf3ac21206d3200a84731f5f47d55eeb8873c2dee55af12f5245015022ee3ef2891327b00e4243a1b6f84a9cf38e6dd676148b958d2276164012de856aa6c00b72a7cd97b0e60f1dc43cc97ed94146e7052287def5caa5b4de3d436ac95c9d33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4944a51a985166541c2306916a0052b6b43162fef759de0c3cfc170e7575d5a7fe3ed3d71d9f78f638178df2fc44431b6f94495af614744f90590a3fc64749555ac1f9b18d9dbb5027f99a95982142f6e96d0aa809408ae36c605d8d8c36f9007a619eae25685e8a4da6abe22c398c30fd5ed52479c10d185adde13db02e777;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5631e177fe57005454945b010311460bec1bfd0d33e43b88c1b247edefdcacb05a45ba1eb9de7a03a5a81a97365b48d28e3b94374166fdc45cd3463225f8d5ec3bcbf80b2fe84cb91e9bffd3823aa73e5b997e9e10319c68162054165331eb7ebea7a33ed9ae81b7a3b85fa0998533fa25fe63df0c36d86af0a65e2d12f6ce40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9332755a6d52a67bce4bc7e162043962b7115faf3a40e7e6fc16e2708143596746ab0a8fc5259480ffe485da7a9951da7a9541ba96bf8690a57a565a459ca18472d82c8aca218626649101a164baec2ba5fa8f893a11f980b2f3570073661abec889c570b62057be9efbfbdb298062a52ec30ed2b440c8ed0f2042eacf2b76ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fa819ca323eac1474ef38eeddd43d4c615607ed8d63e0709b139ebfadeae373dab71d21e86f579eebbb643e030b24eaa784297363bcf4c8403929f250418acc7a650f4d6e2208f59560038828af478f195812a039f2484817d4b790bfaff0e7e57363893367edc9dc5501446c87828541defc647365a74e9555ee609f6d7ee7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa99d29198e19a664beed4d974163abfec6bd5b6539a8893fc5ea91c273df2b6bc078864041cd247992172486f7f2387d4b46fef808a5f8342a1b543ea0733f9c754a8119a3b2b7de931a1ce4765572431c1d4da324a86ab47ffd745e8372807fe52c17d5074578649310faea177883c01ae054bdaa60c918e3a9d74a27447ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28be606bc4c2b9e1f9ce3017affe9819abbc545d1984c09483dcc06863346307bc045dc042bd3e8ae969c8545e5c9d0574b90bd42284853e822627b480ed7d9f9ac54b5ae5a285e9420d7f3e8cdcafb9d8a8c757185d0e978a8ad838da39a4e5a71bc58598f47b5a31472d28e2c4c6091f3843df002fa5adbddfea0ce84a3aa0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52a4fbfe425ca862e2a6f1b99513e0d75f50cd8181673530c01e81cb6440efc865cbb331ad537eca793dd64515f0bcc7c049513762dc8d440276a30852fa5913e7c42d1afa6cf46962982a38479e45fd5cbe1f755f22e709a3dbb36c183357208a81b757ccf1b19a2c5a574a595223aaea93e0a3d2ce8ccc159728f053ece741;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d4b1b1828cee6068a68976cd403858234818c54521bc882f2a331e2159a11e9679bdb51a89d6edf02646ff5416b56cd3525e8efee2f871d468716120ae625f0ade845941479ca747a631541932eef42409f2a4f79a5afe53bac0f71e1ab7e21721971b7bec746f78fafbc53e4f7c2bf4e1b47fa5f3614cefc459f52c3a271ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h258206736dfedf814adcb09bbd3912efe35eb26e03d315ce6ecdb540b61ff7650a3e42281be2ed115fb894e76805abdc8cb53f5358ecdd3af2951b077cdb1677902d839ca1aeecdb4c2e46ec4b03ad3cc1fbd8c7447a6a56dd3d5b8534d75342688c3e8d535a5a19dcf7eced1e9dfdf021a1d5e90831246f6ad922dab3c773ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f5826d936bcdbae23ef98ae3e0c11c5449edc0cb8338b3a3757d4a4bc66dfabee9e75efeffa2d4e4059cdd36aa3cafcda5200741e43729a298815ad17c8eae35fba6c6029aef479682528445c18ca489213d8ca006e0bac32003e7f3cb2244934cc987d8832cc765e672e06deb54c6620020a0ad9ee598d217ee3727a1ce37e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4127181976cd0755ac00ef2e2ffa09e4737705b0d86fddf4b318e05d90a410d83beb9dbb2bb0754b88942f6e91b009c1000b9ce3d09646c23e668c6e41074aecb870b0085b8baba57a2b331e5ea56b9bd2d1ce43533f656b2fe0c642d8cc12ed8ff162446fdd2b587b3b906c0f005786ed7eefbc36e1da5edd3329a50cdab6f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d93fbf09b1976bbe48b8d2deea2ac60c0a28291440c396a014ffd3ba29175127c789456a3da09efb37fc008e00e7e637ddc13729297d411415a9c5f8f9b54fac0199529f6d11d47b02e75e86a68f09ea63abf5c88c2c6ed39ba8cc3ee5e0fea45366028b0c3557d3e4e66360afffa480f1fd8381811e9d3fc1f165ffe1eadc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a569842f3d01411d0bd3536857812bb36619a89593b30aead1d4f923b537b449701fbc57b8c22e2ae61969123eed60b8af086c989784b1342a7333815c99b5800b8d61f03d9a2e109b35b4c095d4ba70adb6576a378caf053d219587b686fadeb5c499ce34bf918c074594056bd712bfeb4b42aad8a807f62bec14475f11740;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45a4bacab6b5a57df3f75724ac9b7f4007a4ac287879fba78b56dc2573a21e17dd8b2f237e09d906c572c72d2cc2725652474e89d7a85337db16b3c14157ac38ad325e12522da5da381bb604ba09002265ba3b6a720571b954ff3db04f4c27ef3d82775b8c866649c4375cf059bcac7e528c40eec12d13e0fa168fe548a5e265;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a474cf99b5ed6a4d342b169971370e78d7bd58a2aa31706797730d0826494cb10b7c219dc49e15e5988a4d61ad677fba9b31b9f94c40a21ded940730a9a5adebe6204998f2bf4193f909a1ef1dade92e894a90021caf9102fef94f75d08a17b2026e5dbf16a8bf8c73bccec8e618178df7fc5a568e34406878dee0d19b695d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31b0b590ad38abdabe0bb699947a7e4b6a97fb8be265807016450cd4ad27ec985fe27bff38157dbe703b00ef882b69ebf5164669c3d06c0334a086448ff302ab681e3e8ae9c807aef82a5992decc4cdf4fc46eb09424a7d6afbf0f6182f910880fed52598ed1cce20d0d9e12e7c1ebe11bfeeb26fd343793494191a3e11be3a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h446e57f8bbd4480b7aa6f252a0dcbd3e42a6ce56ba303fcb19f947b0c2f7017c1cb238b67c27c594af4e2a1405b513b727f8b21e409efe71660cc49884b87753b5f9f8a934223ecc1173499692553c1f010c6290ab36868e6488a9479f7be357fb3c6df9e1c3b48df416c3acd7d6e01eba3bc8d050ea85a4e6fc6b34c1abafe2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd76982865c49f5b325ce35ca52b2aec83c20c221747db0c43bb9d9514609b1915f8de54dda313b6f7b2b74bf3a4dea3cad6c29aa8aaed70f605a70b0507f54c3d2cc577ad408f3584522e7d454a05f341d39c63ef616ae76384c6fb8d6b95f7855852477c811d276b09521aa2215428c4f20acca7db274de9f3f6d28e05b830a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habb5567e949ace7f7461dc328591092d3536611a9665d8f3833f3eea96131ed36819c02617bfdfa59f20bd89b2422e8a48170b7706c8d5bb0cc57c47aa2f9c9d1f51a7a93ac99d82407a1c9ec10c01b3584b9e34a1cc8d1e5818be494f094068b40af3aa4faed9ec35bf04b6c73403e1c14b2c0f16f230b721eb095791d9996d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46bfe0d42a3afba09244d8c632d4cdfdc0012552aca85782ef8cfa307f686e542f85c89dc08102e0b42bbf0483fed43509cf12b0697830e5661ccc5097a93c6f00f521bcd4c8efdab662ce508c22a55511f23bf264b671b70dbe88dcb8408e62fc54c48bd4ceeedb7229799eaf7b2dfac915cd3d6661471e3649d91214aa774f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f58e14c8cc594cd90a82e8b8bd199ae4b53e3c9ae225a487d50dfe45f8838fc8b0a13f9a2e5faee9566305f06237f1b1e5bd518eabebe10fb6b655e9524104340b739fb910e9989b7c838828fa6503a2fe03e1bb53256f408dc492134e251743c5d1f1351c4780cb526b60b09533792031a0f42da8eef90d495f4fc5153df62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1bfd432b2b008f890eed7b9da7f2648b3fd84ed379ce02c2529d6c4fb9c37e0440586e1d86c3846bfcf829d418fb4b196f3f5e7701fccb7f7dc3c5b4420c05bcb46bc796c70334d04e7e10a25b59a5804a18c97a596838cd1e0c0ff9f608812f83df4455c045c405fd75f54919adc8e8192315e23e1ffef6f6ef8d8fe418ae7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0cfc82a98cc6cc4aabd5dd715b6ee6eff3a0316d9f8456e0c99ae63b22718509666b616f2132435b9f7867ed751aede8ceea3ce4edffc9772446528e0ae202c248f7d5aacba3fbbced1a7c75b0f195a087ff47640a5d01fb34ba9ff20bf20019e3c742ddfee9924913d2231eefae5145e936703213ef82c95a6ecfce1f110d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9af993ddfb1e13bb4f918ec6db4df0c0019b97606279ad49e4fe1ebd330ada925039cf368d0ab8bd5a9c417295a9cf04f26b11fc1d0b1aedfe6d0c86d2db7c12ebfaee04d9144f7603d6eac930e5f0c998c9a73a79897ba328690ae6e046f63e7a16d490683487ef6fe21ecda1672a3eca81cb57c2a3d81114d103782e53e4c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5429c57a8946c727104612ce3d9c64e40724e0c5c5c09df0a7094106a82aec2e3ddf43cebae949daa5c5eecab90805414dadd1154909e05f92c9d036af095287b6270bd16335813385371ecbc31b72a3cfdf47fa22d7bd6fcec9c899b2cebad6fbf684cba88fb55f6eeda3dde9796921d746a4a44b73851f4eb1f832594f59fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc073cffbcbbaba6946d36de7e3538761d4bb22b714ed42feee022c3c04d6a15e008e8c35c30103724496aa23a8b2eddd338b334ceb8decfda819e9125276ead9c7076197710a86b2bf77afe4158817fcf5fa51d826953871ae38c2fa8557e6d3a0acbde9f900e0be1f23e3f99a0c467b33ceef3d938f055de36387eda012bc61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4de8379169d8f5eb0cb01cbc5c9629e1e6d21eaa86f5083eab6daf2b39ec3aeb4e83d15b7522a9082df1e740f8bd8efb8446c177462f141a2fb1445800db0ab227e37a235e1141cd228472d7e1be59b404b9109a8a643984a89ddf5a6b818baed49d098ee3b97af46ea087999b154d323d64e6870c9d0069c4a6516051792ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h388b45a020e805a9582f7e20f858be7c3b987543e1b078bcbafd3758c12a2a85fc7b137e8e455df99a85ffbea7b1219db1da4b93089090751dd31633a6f849731f61457a05e3e3c6085d11730b24811ae8f11e6df00683c516c7f6f63657eab30013d07a55196840f295a11b15b03773fba18af6878bde6cc6169f7519269c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha296378b388a8b4dac81e953e4211c481a9038ce282890dccf56b5fef2de57acda6e40cb1371fa11dcce7ff0f5b410d85582be4a555469934b558cd85e642e163058caa738dd0959bfbe876bee50435178ebeb9c66a84d05fad1f22cb97e26a1ab8733bb151bc9f5d85cf2cc3e633497076282df0caa867c922e48f1ff785f01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f5026c0d666a4e1093de5f9bdf1121ec9d38368d5c043b8eb525be0e181834ae23bb1b292005454f63662cb18c886235fb513bdc7ea7c315affc361100cd2add41b7c5e9270a325ce4ec7c0db431a4b1c0f08ca3d91b3f972a2706ed706c1e50580af4f68d7d6199f8ad345556cdb0ff8575cf2427b602b03bb2ab5ce71b598;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67feca2665652566466a266045d9b003746717e2a71a9834bcdcd1e86e0bd749f1a66aad0684b21f203b0b9012da4819ed2f49584afd3f3ca327dbd6e41a588fe6dd5739ad6549f19a79b397b0d085692d48e81ac548d97a2818bd102ac7f5d2aceffe81fdf0ad6e60c485da88ac7fa4d94a6f36789eafe0a96c9cb87d65db1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36bcf1ddc745a17eb7d18563f3c83903cbd393b312ef93feca9b216b7570d5854ba08d2afea825801ad27572d5b681f780807e4c200d0edbaed59a5642856d7f67f24800c2389c03d59d4b6dd732d237429367f34e39c6a8992d5f972532656ec75bf91d70eb20c70bd5581ef8f41c175053d3636e82672aa1d0928608cb74b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f7a893da596c7a4a8483847089df269aaaccf27a8ea9bf4e25874b640487df94ff57a6ea26d36c2553dc0f88acffa5870380676240b1acd825c91813b4c6cb1ec85e4b74e530f2ccd8e295cfa07ac46a23b356d2ea79dbf4e34db5f4381f7fab612bccf26b5469c5fe2a09cd5becaed09f3fe7dca2b4de7ce209dd90cf07346;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a4259d42b5bac4ba6e9fecce269ee91a5d0e17d561ddafcfb177ce178dfc61ab9c76ced6435211721d312443bb993dfdc21cf8d279831847da10ba59e3a18a5495e249ee5b9a0c27cd7e26940829f9e045f36573a9dcb80cb0e71e910f2ab0a8aac8032e3526fb37e75581df6f5f18f5899b48a38a61a022ecfac1a89934d41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7212ad6501f97589c46e9b1409f678622410da17b0c0133ba909a3a41875da5565f16435d9a3a923163df4c1f07a1f70222d60581a5a27cfeb0c7e23b37802eebf94f97b4c75a9608e5a31f2b4630048a150cc1a0f6b62746618ac9200c2a6a9077669878801b1ac54e9a16ed1111358a3e7a57cf89c3c73d28877cd5ea35b02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc50b1ecef5339aeef4385e3397f1fe1769431209e0dfaabc668e4c499f9fec4a62b9f357117eabe9b0ef8694e1eb59226d0fab53b75a2544c736e3ca6b723282a935a8df4849fc535b22522aa2a82a11809c35cada405fa49b91dd037b41674e11b8d456c1210cfcc0b87614daf0c9a895e4eedc6a481dbbd500858b7b038ab7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7f9c98e9c18622553973b86e9a0bdc3686ab166309a50c9dcb02bbc284a7c519e7bde1103706caeabb8eda8bc739d23b09ec4a7e7c63f127dfa7f1a086fea6b24820d1a62ae29cea8c4e5bef8b5cce4d4c984d7af7c030c84b722320711c3416f31b7ca8f224882f89f3d11522cc9cf69b8e86ce02d289b5b6094eb2b04128c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf539170c26192d7a7c8cf5b2ec5069cd85b9659290d008115720bffe58de31b0fcd3da3a9409f94875ba3181ad58f394e326ed1ed645caaa2ebc4a10846ca5df1017a08811f5f1cf0663ca85684aeb1f3586db7b58e0efcc510b5fc2e47c645457e6ccf4aee5f8ab6a62dc5503f87811e0a3174e0b0c0673021a198097915175;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h151be97527234c48738ffc093fedc2c2a3f83f2c4970f761d85ec3b857d0fd7139e112e73b18162613223eb988ee96861bc6ed7abcc0906ba00a100688b73efb05139fc0f9e1f1ae4b3df2a5d8f8762c05c26a45ed6ef05e815dde6fd74de105f8d110e0938b7defb8ac67ccb7a0093254ef9249fecefee03943b115a0a4d600;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cd8e738e7d6bcb9c6817f8d0f42af904c8f7a089be48d2ecaf39b3d4e3c18923169ab7b95d9fbf83ba7cba535fac137ab94e0cbc8c91a6f35622856568df83d4eeb5660315293e316ad551187fb3cbd3b022bc5efba001d584722e0470acb37514da5f3d832f2e943ba796242103490efc9bbe67b86dc058a2f38901d5d4cdc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1367e74319a82d9e1f445dd717d6831de6685797338ed1e32c1f187fb05ae79bf75f7dbfd90bf229e37d3d867cd3d8ca4f317dd8d3b4605b25e52e04113de8ce2a13562190d42d31fc57144c36a67a142dbb60f81e001c2d80b1ad98aef9c05675372b1f510c90154e1149eace1480a9ab8b087cee4ba1b67a8d4c4951e61e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb740e5a0142a2cb769f0c2bfd9d397eef39e4f2fcd19d64fadc08af347e28510666a15a12d102c0530830ec5fae35963d5fe8ca663b31c858ae5a53cb10890c8c3f073030f428ace7d0ec19330b41f7738138f6cc35e1fb0a2a8ad5ecb0d5143feb4eb5ae4b8ce9d69b1560f964e0bca1b5da10d59352a492f76be836179129b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h862dfdaa6706b76a7b1e3a079e1c31d7a2e72c6fb0510f02b14eabc4ab3c4a0c142d8b64d0b62020d167ab591098cf4f700ccfb7f890c7d28c5d2860d178af74480ab109f7dc54adb7e35cfa110268121381d9eab17b7adc373147628c3897bbcec9ac6ac3f087edfb34defe9853a0fada629e114788d02f258c56b16c128590;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha021e00ad775620d9fa9f1c8c53c6223cd6f6ca57ea28e3a9626ba2fa21d0f369d97ef2daf2a3aff561f64a06a9a61972feb93ba96502bc6c427bc26b96a49974d583a07fe6c75e339d77e03d2a8125bc6bf218b74d200cc1bae3c9d09be301194111b233ed79755b7fed0e0b4de1c1a6c3a5e0b64e85ee19f2afbf39eb5cf65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8e745225bfecac22149ce6c1142b5bc299023427f6239fc3922c6341ea0ae55617cf54a78a06d40069fb0a370ce6db4c3451f37d4a51a855f9589df02e1efacd6fee8369222d0a9c71c1de636fc79c861cbfef33d359f0ff5282ff4d6b15423a8e578c5ca9e44c94a32a5693f275318634c9c57bd68694df3228c25a85d25af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3893b173a84095f778aa73c7e2c0d1834c541209f92fa8cbaf126009ba46222d55340596fa1d77912470c1a1fff59a538e00ebca9087b5ef2749c2c7d80bed8a45670a05a446ea85a5dfbb075b6492bfdd84ea0e13b594f622863bfb23bdaab56b30783375baad4409d30acb45e9a0240450cd2379bd83fd2b41823b32fcdd94;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7c2fc229878ec2d2bddfb21c1d81fcf486a9f135b18fcb42f023e0bc5ead12d7e1204be809ab561312d284116475e53d9820ac10920372900fcbbe78add1bcfc1ab6742e9735f19b1953a4ca9b3febe34aa95665d42b6ca6cf2cf57d01ce2337ecb297bc48109d5df5f5adb956a8d6e3aab710cbb04044bfe1b32bbdfe799f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c307471c2db6543056c7d488e4b155c67feb362436e99a926237dfdce7b8116abf7244fa5a332bb3c36674a6e4d2454c7da3c3597f366a9bd900e21dfb497b43e0f726f584fd381bdb1f5652a000892fb7ea8f111be63de81cf5986743e1793eb72bacaf95535c85fbaf9c31db7da62c0198bb21de1f439a03f4e3e2b9d82a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h404358b1f72145e85f9c42df6dc0129378620bfea111865fe9de47be38b2473ced7c44545c01314eefe8371e4e418820dcf22e6e85672e04920826ddbda2c22507d631c81cd497986f8270c6ca304e724d58f82d2aa497596cf4097124157f5154e02fa26464b2cf18daac03beaf6f8d097fdc7b0311644cab2ff9b014cf5afd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3d137d802b356f83879ca5e06f080b7d4ca27b84c28ea0f0b99d1ae6c43e285ad1ca7b20175100bac1a3090c43ced2d45f9124b126647770ed0afd363bb72148d75695ab905b389d98a36c3667d1462b77bb4760612e574c388a0fd2e81004b45f2f582021fe5b4ed9c6497dd41eaf54659614516f18a7fa64ec0f360475d06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50769bb620e1eb2c5108a8aa86d737eac6fe3e3dceae73447b7d1820c5d201e512ec3e5903e2ebc86cfffdb61704c5377977fb9094c74e792b3ca14526214fbeba16c3b792271093421a866c900b186fb0c19f1473c319983e2b34eb4c7b302cf587de6111172e1e310954fe8e05a2af8d2e7b27d94d316ec536d5d1529a4665;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62b95444a957872ed6bb231c552d21110938e6ce361ffdeec89e931d4a82958b9bec8afe7de9bb7aad0acdee95de69bad915f5cb8cd6d42870dcddf964bb3c9709e573643777fc3f2e7231d2ac7af2eb1ab47a1ccb23b7809d710f926c64d1501692370ad25960d1c62aafe352d48607f27d5fb847113fba3f7f83c0c6fffbdd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a84c984cefddbb878fdb0efbcb8c058ae47e1dfc07466a02335de85291379bb67e55734d2575d25a7558e7d8b9aad626b5aebf0988fdcab7514317b795329adee348e67b24577e39713410760a3a2c5080263cde9481ca2f305c1a33d537628f4d14590f052e22c9e49f06c6a55007252d39ecc28420d565f15281f09b1f7c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5ca008574e4ed6f7323c7764031a7743a744c9de737b6990e0a7f411840a092f0f8fa78ea8380fef0dee09ddad658c5e39fd5fbe6cdae7c33943018bc6280ff0329d487bcb3c0c85da7b7ced8a700b84a5f182d736dd32a547b55d7414f571ea4bc1e3033c16d76b33df58b31a49412eaf28524da6f6aa29868fa0507b9d3d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf25415f8efe2138347b32ee21e19523c02c859c4b978b97495149b58dfaa211b7511e85c34f84be055a46ec22685a6ea862ebf48d9655ee4b89cfe6716cf42ca1850598f38e84874da22bc1f7d64d33cb0bc55c956bdfd9a5fd53b93e962d53e05fd89e1061f90655663007a553fd54e1881be3162099ec66114c93b479fcf48;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e2e9156db8cbe8e6f077a9d38edb304ebf3a6d125b6ae21e4b75f1c0e2325446406146a42d0467a31e26d2e08a12f52036a405df2e189bd11a0567dd62735b95c95d9810e0d1ea54cb53ad208016a517befb72cda17843070385329a69b5fb26d16f1bb00c6465ebe2dc4c8ce9cfb1572e3bbdf7d34de9a7257adf611ddb87c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56b307fd8587145e24315e627387354464beda60cbea57c2684082e26d61051720e017523d3ae6a15c257ec4ba6c8826a4347d808f878832f7216aa5670f41ce740a75ce42e5a6ef880da8d2aa7a9a5f40ddb2f309ac40fc524b8185a9465e31703a4fa245301cfc1833553e4a410b0fe934f855e3394600972e32fc858e3ab7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e18a535e2979295a8447bb38ac2d0d7d21067f57990af9b857e7ec5c855696910b72b2ee35525730e4dfa8b158077668b02cbb3ead78cb36296fe0512803cf87669ade7a9f8cd28747e46169cabe190a01e2dc28a50e46df3fd3db8737474a27f371c0b54f302fa2d88c0ac110f1f46102666c6cfd991273eeb0ffa32a54ae2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac56e77accf63c372d71fb19a64f17ba7f955965da1f1c35cade242cdf02dcf4162fe5a49e935e0ed93f20a4d9651c42232bc12a413594d46f7422d5f2bd9194c94c974ea71655d4f67a165b8669d56e28352057f8596e2b005dab9ed5593282818b6d5ad26a8c9f9eee3f99d6b8b08e08704831f7648f114b97024b19207693;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94e4aae94d6e11bbc5383d486518f67abbe89de4dced3886682484c668dab237970aa5c4345daac1d219da44e08e9fefabd6f7de41c4d539b43e9390461c134435fe2b1535ddd6baf5ac96242ef4da40fab19765cdbb6e4f0f7f538e860326392270dc9e1ed8692cf6a609d909fe4b149212e953f8bce9ff4c874822857e526f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2682d28ba58085a50503f98028be1eb5337ca1b5983eafe4d93b149a8c70310cb4ce0743e937d4a81e014a09e784e8b879b89336f058882d7d927b88e2a53a254cc3927eaed49111574bf2e3b112a3f2334e85ea89fc5760b889ac70ad8f32b8a24d410bb83714382f964fdbcf2bcef100cd80a4e2538f7907308537f267c7e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee34d6b3fb4818fa32a581c3944056843b6340aeb71c4897101174d08a9cd47a006842c56a8f4fd21cc41a129a21032de7f778c8cf1d39fb3c1b1fadc2085b59611d3cba5359a5068cc4585bd6cdfd707709dcd73d05b1baaa214c6cc694f9884aba60ac147d26e4476522931c4b3273614d2b063d455500b341bfb2591fbe07;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91a1f97aac2f6065029fd97a6ff607abd56067c2533464f32c4f89c60a9db2230b9ec36e692f25c4407d1a99e72c2ce37b7d5cfbc0d04ed7b8acb7df0c311e31157f99b1abfbb0a9e953123bfb444d7665b361bf8965de3933882b80a9cbef3cd5c6f87a3468cf837401c62754de92cea9ac82cd73073f27734973847c8effda;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d7e6290cdc782b56ce4d39fc54270f71c4ee1dca901c32dc62a2c2934a72a1bbb36c82759299ac0cbf6fe2b5330c95bce4ab47ae85f65c35519b7e430f8c9bb833be306e9acea043e67cacdd6d33d107a9fa1d254b60a7ee942e4c5c90592f77751e4639aa4ee1849e18546b5fa3addd8df44c0c49514673e2bab4927c7bf59;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6237800217f3ffc7fab77d4ad98ba6e1922c471f38385f7ff286cf2ffc41389e5f4fcb82c97d6de8da8e6e393f010ae8777a8922ea2ec281e73ed41ad1b4425118f2018c45dd1c5238ec12f74746cca1f495d76647664c93170a77317f141a488d7bef14b885826401280dab7ec528599b7b7bc03a7f5192ac5f9d588883ca12;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81de610e6e509c94cd119b06d207d5fc54b129f9f5ee2712d88f8dfb63e8b51e18615a8375f8f1552bffbbdb7f6248d62c933dde6ad88666f20349b4176dde6101d5e3f2aed4d1b97f23080203f3b4dc0eb38f9aa2a4f2433f09da7e3be7f5ff482c576a5a613fd03cfb7a10980528c1e754b37834dc34063a05439b23e94349;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ca4c1d112d9079436af76badb8e5301a2c754bee8c35c8244980932aeefbc5cf118ce9ba57facbbe61e9195300acb2bc906818da7b7f3288e59b3a570b2eb8f14d52f5c197158fec9a77f96a6f831e1f5504bbee7fc5c4b0da351cc9e46bf1e296a28ac188895a9249ee48c3a49db38d4b20887d121047d9e6b9e3bac5ebc19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h369b35500fff1dc0c8b8597aafd4f8acfc33cf60d49dc370ccc52a8ecac3a74c6cbf60e5f8652da2465abb65f1eca5997808e7fe7f90d5f8723cbde37ffc9ea185d2225583a135d685eaf41c791ac9b1dd8a0c29ccf9e666606059d21eb4a5331e894ce16a540297131ff66833865beeceaa0ae7b5da679e64a080a6efb80cc9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h638dacb576ec8e564774a6a6d82920b2e4702e909f9d150acede414cb1163f72a73d8dece30a9726174395fc520d982f16eae9a608e85be8b48498b89b807b57619d82feeb71746cedb8bc2c1d5141c6208f5e01605dce182f92da217e1d52f053f847f4373d909c13b292db5959ae749c7ce646ed220c82308b9d306743bf81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6fcc6e98979f03221e8f4b4779381966da05dff6546236bc845c5a1d2b4ffcd99e8cf9df43271de4c696ec979fffeadf8b4917d7b81184f3cad6ed195c9276da2e980b9dc6eef246229dd97b6f6d0aea1b14d4b7cd885eba7e930529697d4732a546e76502243b624540d2cdf6482102315daa3dfc7a08c8688a22b2f035298;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79495ab2c5509044c2770a8e4605359ef0fdc6eaf85baa8b7a49a9863b2868a8a1b50bca789862cc62f58bc024c4f3579f9e59bede085e773b3873301730ed0e36b4cf342e7bca1cda67d65ab4ea87ff5c25377f89fc19e48a6c00e0fae31ef61de9308894f18a85d8b906f8df0b6977bfd398c0a0c21522388cad6e1327fbb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9262ffde7b2503e6f946d6f7b1396f4faecb843e310c66ca28a41c4a34b9b461ce10c272c2604df956e8f60680f68391ed96a1889c9b7a032bfc56216f2ee656c261ad649c94a30fa028e9557bcc5a9ee8697cda838f1559a1b4c0a5373550cd56d79cbf2afa89c7a85ebfaf53e1d3b3cd78bb04dcc28bcf9692768308d7ec2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdb7f2abfababd7fbe72328cdc0c1c303998792becc3af9545cf33c2c38e85e6ca81b24a4fb566b7781c6e48e90028c986abdf675f40a7ae352ee52507704ff1273b973c156097519aff0e945891ffc1c1015cb19f4af62d3fe3ed5a0caf024c098602f5edb1d9a880b737dec23c182be6d8394f709e5fba6e8c8e22fc4e2f3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbaf6ebf7c1a9e50b97394461ad23cf95d16f41b5a3133245b4381a85bef9af4a4d8334b9c8f240b071f6076f153c12427d1f8548b950ed1f9c767d1ed63bc7b56bf341bd294c71b904bd98e183bd5400a7152cdb64053a73f3face687b05d1418b9da2b73b46e0012e0c101076885cfd6e951b89077945c1b8b9cb67b1aa1f7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc2f0b55a55e0184c2125aa357b7446239c7dfd581c56e8fec759535f23c7cf8c482bdb3ffc033fdca3e1131df7da49277dd99bdeb0d8bb20a9673dd9957c726218b5930901f09b703d9d29c57ab85b4aaa2f55ef06363dac0930fc464a5382bf02915f9e53e5483a769d366c43a3ad95d5fb87b872916eae8907444467b70db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc6622ff93a8f96ddfa421ebe10da22586abd7b1ea48df9ada8bff1ce81b2a24ccf9c60e95782c00f4801244c9e869f54254f66ffee465a76d211a9b432b65ab4fe0e96d2d9bdeb93f001a0198ab635328acd2cf0cc2eb40c997f20abc7b566d7c2bcbcb93e53b1684141baf11d80fbe6118ef6dff4cfe8ce3a8f4f2e68a44f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2017d0a71eb7f720cd19cd852e7b061d7c0998b8c2bafb48643be04092003f362b2bfb256afe900bf77d82501ac9454652564fee8e69d5674229b7ed2609156056bcfdf65c76e5192868a15e6b41b359814dd8e584cdd91fded6d8c6180a453650484c005b9776aae5a28337c435d00e755e1be4b7c06a2de76d8a3d83d950dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6035d633a2712999b0e34dd2d2c01a8c99d9bd5c34a88598aee373593999edbcbe2897953264272cd0e31dc6c282132ca55b23931ec5c832ec6a1c69d2190c46fc058719d5b8bb7a3b0261ea0b3664063043e57b61f9383992de48ee4929fb00926dbbdce09c33a21283e518650098af420b9af0b3c87efbd87a50065261aff8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he696c8861321b6aa52594958465d6720b68efb66adb18af0ff9b1f9a80d318ea76e3e325f6de6c4ff0712a73fcb17daca53d181813b8c3319db4c370add1e632171dd8371e071f4c7d515f5c8bc46123387a70f50d3cf40cb393d63e30f0665b7098a59d80f01931dff51c781941abc2c00077e985ea6df1ddb0f35dd3717418;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd25fc8616bd0777e41ff0399dc4456c884b6985db73c08da7d25dbb1ecb48faf5929f1a3c57f95cb709156f21d3eff506989909f6a0139bf763c2f1c7702415479fdf13a496381a9cb09e176b89394bb6fa7ee1d205a303a46f95c2b138cad9fc5a9d19ca54f66f4fc2b1d28be57afdefd52d489299ff77238f6de3fe2ca7dc9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf4623f11f6d64fd788c2fd7b656fe9f5909b42e4edbab1281e3827eabb7ac0e08dde0809711a87f90451b7931a2fb615dc171ed540fd73e73203b572bef463ba9f01a676ac193881451883a7b94996c9259a1a5fd9bd3307f891cd63e17141fd7e23b269e7f8c34f5fe98773bc3efb99da105ec45142766ca787030f485a611;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf80d3cd32810e17c48c99ccffa1853236d2fe5d07eb683d17a4abf70bd862be275f52e8fc1f6b89c9772a14f28c02c4d8a8d6c4eaa2fce16de4bfd0f13acf1b00d9df74ea23deb2817c7987a8ccb6692155c3e3936ef1f182d9a509aa3648594303add929728f87c1a204253e54bb1b26270f4486fdc70b488d5c165e591c3e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4b4c1fa38ffc5c72dc26639fd7d918d0e47cd7deb69209aff7d77751e832f5ff45ab76fe3644a8784394cbfc59264869a2d7bf59ed962170982c849d45e8e11fa016e30ee9a6b331a00ad27a393af20585f3bdf06e53868c39b4d853f3f8d99ee494a976054ebb80eb734e9449fb01897183c0ad9a95c03a105942c2baa87a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9e1e69a09b3e83d9dfed3279b1690ea9e97ad5673dcc19eda2bf628d1601989364f11b53b1868bb387f42f1a1a781b8c8e79d8ddfda5905fa5ae639e9ec7779a3dc21f2808157714f43dd5df3a6c42ebd9a004875bb069c3e66fb7f04f8e6666057e2b97656bb8134ef4ce3ba5f9c993c8756d3bf471478d5ff9ece518f893;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44769f41d81e95853443a962aa2a1fbd09d9eea25e34203a5c01b973f2a40e144990939f9a764f7eeb6268cb1b2c918943f16e59db4bc19d0518da18d7a5c3feaeab6881bfe7719d70057744c47318e774e3e47e1362774b437abc071ae6c64d8d99a6476cf34be616ea13c97150debf3af726118f3f46b54a65cda97e011203;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae37ee4d192e2d42661076f836b2bee860a62af0bacc81b1774f9d1a2e6376261921ef8c6ec16a095e1fc8b4969690c01aed76872fcbb753fd99e202f6685e8f16735e7720e3fa19305911a2430dcf9ed4d6b781d898cfd6c3974233811a0dad4e84157cbd9dd13c45ce096096eb50153edc7d7e0b37b731aa25e744566405e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2864a4f272ed9f80a591cf3252ae80b123f735fb093908f4e7507f5c4b7f656417a17e6637bcf94a708909f03a995a01609e521af4ebed41256bb1ff4eaf9059d383ee2f911767d9daaa934eeb9a63dd8426d865335958320a0b35550da0656d51087610d04287505bec9a220b1ddee67be0a44eefda778b807a2d502c829af7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h934f61175232e4b71517bc45de5e5ada87af5444425c8b49cfa3f6cc046e73b4e4926bbfdce4559b98093973c7824cdbbcead0e6ee8072fa34c3a4e40f44d21070163a0639459e428978793e8525fa05389ff1c9f9b9b00418b488f87d2d1ab4f6c851f40de185ecc46fd63f6e7b923952b9f4a1d80b8ad58bf2ed3b5c7339e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ffb52c1c93473e7d0896495be7394a232adb32613d20f4b55f5a46a8b5f33f3e19689ef99bb2c1b4d1dcd87dbf9d6fb39a73cf64897a2556c20860faf857334a45cec10821a9258c3869fadca7a41687751b5db1c7eac9ff8827d825ebd90fc9525b50884e9e6e0dc706693b0d701ec48379e9133950a4d995b561f5c1d0405;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a6d760dc44c51abb3f60789f80c2e57bba2f67e696bcd4eb20ffde87d7d0befbb3f04423067b94811ea0d4e331752bef08a13ee547ad38592e64e809efd0d2bc7d2532d3d74ab9db1cd17fee1056fb2b9bd580706375697d1d379d165b41788e11e85008a326d1b9ee9b11991eb4fb59c9085da9799c308509730ba22cc9893;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac2527d3226b3829f1349722fc903ca2e0b9d0971ae82db3563f9b056042549eac4d70d72e97568699cfb37240c6705f6bdf040a71d198cfbc01ed3ac782da7297a2d6c07cfe17f5069cf03e181317cf935411a365aea59950aa6257055d0127062a00d1d24b91fbcb325946e799e4676d43aa49be854c032f35372858762a9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha39a04d226a2ab205fe2ffb8869f3c8bac64476414552fa7cdfaf80de4cb5552f85d25ad468644d69eeb3ed3f25ab27e7f0225031721eada6eef13970ea4ef9ab1aa98baf2ee8bcb710236b8f6763f04356489020134bcb65a5d846f1a5f9610dbf5c7a224af54049883e42ad4f80c5ce461d5426a9a65dffd0b35ab685b134a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc09d5c181b3e83f4cf6984553b1bd4bff991df24dbafb81ad903d6a6a1c3a5cbae004474543e5218d227d49c108da85e4876f9979d2744fd2dd759cac38fe566890343803d5ccc4d4337f5cb256c2c3daea5d7f1201e394bd10a2789463cd87361399e10f48ac4ce9465377b2a25799d3476ddb1e4aaedf12f73612a81ed7a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fc895b3876dbe9d97dd048d128118f418e49564b7c45b42a586aca842fe931c27e88e8029bd7c3bf09749f029ccac749acf2003aaaacff3c86b4d10aad4ca9b9a2a21e78c1e0a79b2c662892f865b7776c34233f1e97443b8db6c0c41ee5c5b5f519a6bbfbd14a2057a66dda9d107777dd67d75d530c1a8bde6d25706acb149;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4afcb26d4ee6058356a7c5d75a779f6cdde688731cf9a092ab3d69e1410f0f13d6704a164c400c2926c6df62b431ff250cf38e73f026a46da466aff48c81620f808bdcf311917c8f543bda0d9ceed5efd290cdc52d44945ae28c03b5b76ab47540e4bbd0f76c4e809d2fecdf20099d6786ee1448ffa16e405681da4b096a1927;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd52e29cd7314f202f0ceafcb170e5ef7565e512749d811a55fd312611d4bc855c34b13211003f9798e550a6bf67c7bec25729d1dee99fa6486265ff0986649b24ed4254ad081eb0e82d3ee4c815f161e79a09654c0183b5e33dc23e4bc6d69f852a4700a1e45db2a9508ae0ed962ac438cfd42f1920eab03f2293c0428de577;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa0b0b5f8b469fa33a73488431efe44f8c05826b22b6b53a717e28d0ee499a975f6638e12ebef44162200bebbd550998177baac33388d94616cbd8ea156519251f733133a5b5954629bd29bfff01be525f5bccffdb042ba057bf692c68f76e85b11c2bd81f4be03ee7a9ed745a9b65458b74a096c2e854c9a7e0bd5e7cb14243;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbaf461f76ea3e260593372871f18ab8488b8ffda0c6731029768e20bbd3a7d9737dc41a9a52ef6258306a64c652ab8bd46534aa9f9723b1ac8386cfbb6f9282afd0731af593327e8d15d9e4f08c88a2c87af0f685caf2fd2159db5e46e8d0b68fffc9083326cd7d08b3baedfa5a8a2412381a0f69ba3c14c25823ccfbe75c4ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5a359ff4c56838284885e0c374cc76fbb1fa02f3e28091b851822e2f0aec4adfa8e969e957dee7986441d3563ac1c943ee8e41a8345e7fb333cc56321717e64eabd919d99e5891d01c815f7c320c3d3b375e229db9ca98bf3026e28a9fbe4aa78061ffe665eb0fd0bb590e894451dea10136aefecab06916f91374c484e55bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc0060ff09bb4290c928c53681a84d547790e043cded8b6382da680a6bbe03a74c65e3b8059e93f16bad3affe36fb88c274e4c2646a70896fe5113d9f90f634a3a13c787be413102874492b9bef63b608f661ca31621d580780f8897bb297ef1c3d78c043eae55ab52da770289b87bd46baa14b2eaf94b01c240e9c449e1e29a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91304e74a7801edb589c22a8bd65f3da1d9011eabb634a801ec5f94e95a3e63f73de5d3b5e941a766053403d1b251ff3e1e7a2df4c42321bae2d2fdf8626d571ba2bb0e22abbc1d16849f674fee9797d3725aab88c833abc77d4d0c7c095ee8f451f51887ea107c292dac586200ea3ee386d8693367c2895268ab01ff2a19fe3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73f20e7dd22d274a16510eab9fc71322d2d590d225a7e8b6ab2388044a1f81f3f73e2d90ca1f20ea8f9a9ee241e86e2c223c4a47db82c4ad989cf2bbdbc4fd1e43b40adacb91b4e7e082c3397ed401cd02b547493806de0c0ea99dcd6dc1c76d48ab4494c2c2e1c259c6843922d08fc798a138c1c2b74757d93ecfd1be6bb591;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h666f2258a1e46a603135a60c5d258256713c931a1784b0e15384e0876f44cbdd01525d76db14b7d614c07d26a5c437560d7b5fead594a9671b7a075971eb91d7e949d6f0ac1f2b05665fa37217c7738bb6588ec71744c65fab6d955f31e03215dd9f6d0acc89b3f64226e4b7495e07ac4b19a003d5ca3067c8194812f729f01e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4461635bbbf78fa8c2c8a8cbdd6038bd5445f8a08f83df9f4eb2cc4cbc9b2ea12510ddc2fa8eba0f0458d1d66ad96cfb790db7d575f8a74173b8255b649209ed0ab4ae89c5e7d0e7a49123e2cfaf4f06404cd82773a8b034e8a37061602cb8af1c5b6177a25d4523114563c183dc9bd28d765215857add9e87ce8d93faedcb3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30a972be8464eda354994949deaca8f32967a1572f8d3e6dcb179531f9080060472cb3e275ae7a3bff8c45ede36ddc0b60f75356aa6542e6dcbbd3af2a367b660aff4569419dd56162b5b6606639de417aee54c1b62b54e740c1ebbf7aaff35671f86c9d81de9aa1c36d4485947dd01d378fd77cd334654afcbd18f5b45485f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a9d137a3504e3e9d7d57817685a0715e091d58af931f4f8007a9058fedd86acc993ee1060a6d359247c686ec5be319ec60ab802eaa9837d2cebede3d686b244b5873f0f10d1d61f9c4ae5ffe566d4666a01c5bb6d7339363fa1118d14eb838b9d6c1f397a2a6002bc71f90a5f561df549b91cd352a4b4a5f52134999a6bcfb1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61aa69bbf4aa235a80e4482ef279870ae174b95c8da78ae1a65f2d349e284385f61e2e7cc0849a060b7ce704c3d443f75482e1e789ccf543fddbaa008264899e3336986133b886e3b6776c9f3c26981e48477319d5118e2169d1b91440b278b2b7f4453211c6a17f903ef8612deaa52e43c13105e843c96c4a62000b36c4c0df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1118d276d1d527128f28061e08b330273ff3366e3c38089eb5d4e0411ddcb1e0fbb9258554efc5c37397622dabb3bccdf78682629bcb3e53335b3dd66c49e6b9ff08f2a5c0db4230785152ee5e564bae31f9905851d863cf98e63fdae468ede046edebf10d4782c469448cf0e427133833f812460786b72dab9d07fc7905e984;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7233883a4be66d29e457679176c8295ea2d0df834ccf9075486d7e7a702286a2daaac894a9a8f2bf37ff51ec1f6f3c2dded3e09c735a39f5e932dcd47298965a72d1af7cd56340d7dda6cd44de8dec97322c95774e39edf137c7ba6b9aac0b11a52f9b3c5854323e9a8b48d4c0819b27770743976bbd39c6a70cfc6e219aaca9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1260edb1e0fe7305c56840103018a31e7277a06da65c32ab9844ab660209c110b1dd9f9ca94599591ae461a9552ccd0bd3654133f4e5661e8c4bff423bf28e64790fbc979bfb6a06a8182b3a1a1a2017644f8627e27f321343d395c40f8ee600a75f6d37aef2909e2aebc251b6c6b61082b0dc151508806fafd08005db361bed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa26076c7cd07c1ffd3a53c821b945e1318853e97b2ecadba2e0393b8da8b179ab9b3849bb543dd47b582332eb5a408b37ec966a8fdb671e7b54265eff81b71a5c98500d29747b3ca9af14064fe782bd4a655fa3eaa62e9881ef968e706d2daa907aff9e489d97f0304d22c5367e3a8943cd03c03855d1751c458faf013e074d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he63182d917c125497763c15c9bf7affe57c5d6361559cc384bdf42201224906fa954049279df3e2b25054996cf6df2600ca47dac8104ee1c2ad0abb3b9d0eee975e9133456020f57fb321932e9eda8387ccbcd97f3645e169dbbde7b850957bc4ad3b487ca4c7bc5ac3cc4f9a7646a63532cf58aaeed5cc895e6197ec0b44435;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2156427f93b1c36507741da857cb664965dc758e0450413fec6eabae245b54bc2f342e51b3ecce4d9fc18319861bc5abf47a4d7c224e4fa0552a0568e07de269ff9dc71761a1a176e6fe78721f6479d12471b81fbaba3a0bf5a370bcc2bcc4da1379cbb3d50941fee8677317d2e78e06e79b453c0064739aeca739d052518ae9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2333453245d2ef8acbdb15e2531fd720614816ae260de9c79058ed65c827c8008f8840d259efbb33a2e43f6b3973562ecf9b61c5a6eb96c7abfd9f223fd5f26bbffdf0eb9db05ef9cdf727e54773fb154a437733c6dce73b8360c99a02c869a1008da062e7af0262adfc20e27ef34cf1353c4ac0a0fbb1b787f7356d9958e219;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha967282d73edc6c2a64088da78c5ce5b235e256bf248cb66d4baac60a756a3abf956a448fee1042b03acd85bdf1c6379fa144dfaceefc7147c7417445b6b810261b8b83d8578518a6476449242b17b550750277c531fa75e24a1bdcea8eaae2d28d268acf4b2828d15bd3696aafd11eee8cc9027fcb52e93f6fbf59d85b9e294;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha54c52f54ae320b4c2980d902e67ff366ec43f40359c81d33eace8218973c6f77cc81c5b13def2fc29653f4be83a9900a0a2bab29618cbc6803752ee8dc0a46c86fbec254238741aa6e52ae68409ed88f940f58879eaeb7f873202ca1c195b987a185f2e80be1fa9d53d385cddd1e5faec136e2641894e56351b479d7426fd79;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac2737e8ce049faea83d3698899b7fd33497c5cc71aa7fe108a37a94f8e6d4dd8c412830327ba30b5476c77f2fcca3a8c131881c4dab1d872012bf2dd48b3516c25029e19d150c784296582d8559a5ec5b553be914739670e06df57f069dd03cb35b96cfb1e9654076376bfab3563c8a193ec5cf77faf113882b4424a532e2e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26756c734dfa56b770fc3c79485f6f2830707f7516829189ecb0a73bff3c98c6801754444481b040c2ae097a6c2741056d305ada83dc03c16eaa67d418a582815385c698f06363c7b6836fe33d437227f6d39151e853dd91a3568d68b8f0c3e81245e36e7efdd3778f4e2d19b11257f77d573c38c8ce055451b2dd399a383e60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9be41bda036ceb6e46bd91f27356e211b786bc90ed3d98124925814c219b3ef217eb3582ff501bbd0cdc84b88895fed6f38183573b3829bec2d6467c993a013c4c623545b28506eb7123a93a18cd8f54f5c65debe81b8645785206995fd364b2f24fb67059b662b748611d49d741364493dfbd4fac01a6089a7c38332ce1864c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb191c5e044f167715371b7add35ccc6925497dc9e43ff1c0eab1ece0f379fe3fb20d3d307cdc7e51f9140880e0a07710e467215c6b04a2e358c77b9d86aa13e7310dbe97397b81215d2fbaeeac53073d8f6f093910c7fee6deb42863f60a10f6ce88ffd77655b1c20d502c00f802913bd85238aa1b92a3a24053fd8cd3e3d4d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c82be6a29ca4035d74e2fa46ab8ac040c3e05a8ac62a60af906307f0bf9fc264148bd31697a28f42ade16fc3e5464a0bf654ceac90bba1a6051ec54fe8c3150dd5631ce1ca0d9fca34b6f68328be137c4ca71668d86fb31c916b8740bda1ac3895f3b961951a8760a91c8b9c5fa0e4fdc7ef1a6ae0304c82dafb51850c4ddd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a37d7f56e80566a1b39e03ea1cba63fe008b8bf65fd8ed3e98093a0a052e3cdcbb9aad937dfa634c260357963a69d098802ba3e486c6d3cd8154a904b1d02333cf5fe8120658024d03952aa1e99809e6efb6699164c286b06ddfa5e8df476ccd362b2a8727474bd51f61e9ffe3bdd54ec65671f890063506667d9554804822;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6dd43a3534838eb06569b319d59481ce2b6979a998501c3fc83f1da5412f4007da0e48de6c6a992cb2d773a858dfc6bc937818aded0c7ce5907eac2929486cac94bb3eb208afcd22184b541a7a6d51f650100697cb6e812d0fd3e64f756eaa752f9252a57f2991ce2b509867306985c7b3fa5327b215afdd6b8058706435f9e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc87d0672be319ab79ad8e3f91af9dcbeab7a48a034ab9d415f9996185d5c1895e7f2f251821d47dc9f52bcc61bafca7051d424bdc34164434615d541b0db0ff2a750f4e87acbac93780ca1878330d9c09f83a0e11c1b1a569e7c387bdf3e0e297d18f3ba3ce65106ab406bd9be87393c47984cea513f1f8c6662798d36319524;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94454db59a81824b090b11a5905cf15201dc4143a8c554ba682e760c5735c2dd4e2d3998f02ee6bf2ffa20c985fff763c37ccc494abd28afa59b91269fec01bcf496549ce414818680562b975e67a5b28af0b8baa3e9f371e8e4d4767ba6401d36bdbe4fb25e664217961d507639179338fc21ad7b1690576791afb9e333b600;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4ad8265ef8060e8b33284152d6640bd57c8598c270aa2b4f7c50700a84f0a3976922b3c74761eda1d3e470b58d7dc6d044dede487ba8687134589b54a30a79f452b889bd159cdc5c4c1d58718ccd11d6a27ec4935fa65d3cf6a2bfbf853c9e9e7d83fc2d0710fd0b774b3cb5bb99c7218f5c7c71965507527147c732386fb1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc489b75f3f0dec6d4ba7eda1e394b1e49e7d4fac76c48a3479b661421b119793abeef71f5579298f7416fac18f632b2b4985d13bfa7465a2770702844da3117562a0b5ed6a357bf54bc57fe2ab61f3ca1a8cac9f9c36e56e99831b6f419c63ff5c803ee7986d0861f345efd0f5e6ed9ce45f751ac66d7d4615a25267699eaf1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc4763153fe08499adfb639de01da35beb2a181c6335e1842f0823de7da512d526d597bd205f6fea8826d0e9227ce767169cf2f531e01db7863ed3c772bdeb2f50f0d73cf6877eb05f0bbfb52dc77b053a85b6890718aaa53523e30919284a4d543781e9b28065ba3bf3bcca91e3069b0d788eb51c76eca9c66b7d458014ee06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haca0c7c970e7bb8ef05c872ce4a9073c388249ed2b32b385713422e9a926f3fa8975ca8bd822295939f8de87a7728cc00912372591192b23335289cfb7fe7170d713b63f6ad7f89abcea05911ef84cc44cc41b1218e462d47fb734c727fdc630b76713f4479c59a09318c9e55fdac877c6bb95abf20b85a1a6cad220b4653ef7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83b3a6c2d9346787ce9785d0546670f84f9a03b0d421569a26ce814dbcd9fff9dd289a850b36d81c8af965c4dca87c03d27453705cc63e82c786a6eb2854e7bd385da5b2f822d6d95a09658b2469f330b087939eb7c6848e9eb445235246ab858a28c0874405974db5e8385dcffcf968923dff0a02d1e0dcd2cd8c0416246bdf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8a9aefa99f3cb480cfb0483e3965f53ba5db79cffd368376a2f0d652a1ae186cf85af68e6e4fd393fac68ede2609541c624285e968ce5bdb7e0c38e1f6c6574925e29e8542d2c8561a208b5916ff780e17dff4b15271ece4a912f99fe3af8cf0403e2276883538e3139b4a483f9d4f36bfa385bd191ae6477f356a13a79b1de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc355b1beae62ef0cd3e09c5ed7426872af03d247babdca9c0487af985735ceedf0242b236cf0f25d0d2dc2af357b885437153a6fc1f4cc9536eea3f0e66db4b390abd4a1b5a975a776352567b48f7e5d10124f70db54e33bc8f231ff88c2dc21220f18a0b5da28de4a8697384436c50b657a167463ad3d49db8f0ec50e9f6b34;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37b4e7a395e9a82f6ab6fdbee47cf19aecadab2301c4f659d3806c0d43184d6b84e64793d3b6d777454e290b9f2d4dbe066c0b3542ec40ff997a3e15fe2c33da414c92d91936cb539c4cd85e5d21b6e491fca025bd7c1bc94fac2110959b3783c58b5567e0b05efb3dea2b0423576b929e512e4097e68af2462ea5c31e7d1e66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf3ac522e7ef58a02eaf001e4f775d43f801ffb6b1b031d1e4bf2443f19820bc42f6727102e080a3d617badf05938e2f241f58a68ff50254f65e6fdd71a59cf896d9bff5000d7374bf88343e77ec1e40fccc10de16263d3e30fe25c2da5c57243571b550f66c06c5e1d92362e676f86d95750174248e290f67c8ec218345b292;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8f87455d7ed36fa67958710e687726d3f5ae3424cb9ad0d71563d636c8ab97d561080dad821654d11695cef83cbd76af39dca20d2dc12db7c4742e13e01cdd3f8a3db98877de38de5a36991f7434791acdc166c9cbaf1e452a6387291d259769670393ee8f234e08ae63dadf0788fbd76a67af4df03fba904424e6cc9fe1400;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3534f00887af2528ce6c924f9afd1f1a452e86d18b1c66742488d6c7584f124d34ae94a6730302f16980b1cdc7a02915105b0507e2c76392453e6e79172d69018dab9b5e606fcd3886ac4b325ff742991278121dc3816ac697fe212adef22de290a034f92109caaadbee6d325e69319e437cd623fc0e29ae7689464faa2f994;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heca5d6961c0a417e5725c04be3863b116c9fc6b625b58aea93c903728ef5bd1f0ef75629cc90dc3e5ed147a0f951ff0d0b88df58fded8995dcdec2df41c54cd62687019b364fe0f8c91280e29ac7a2ab22326c199a7bd2bdc30297675a8f9966faad16db948588277f4f19b0b2465821bf7c03d9e9ec89d4dd7d02a3f6c46ed7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3aee30ac6ef6d428714d7b44a857fba32dd5d9fcc477629c525df525030d4e8ea2bd9a3f929d2315f7121924505e1b3a7a8f629da60fc4ea1ec3475548200d69135b3ab34bf44cd61a4e3b7005f1d5aae6523438f714b8373c40a3526117e42673cd5f7c6e37aefc201b8f797fd57a2ecf740ed17f2f60fa083fc76a0f86a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15dca47585c97b6e63d6e03d26e9d8a9d413d2382bd81cb511439b7d64c9c5f5833ec67271ab847ef5283ed0c5a36a66ed05f7c76a759647adaf21df04a4f417bc1a5d8b55bfb1d1cd9656f5336eac84e952ebc37b5982d9aada9066007bb041841542e9cdc33553209226c4b7bc2ed86a360cf758da274247ccc88b3a41df7f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha40db154f384e76723cbc00567f7745626d5c493c2e0c6a7815772cf1de0f4454f3cf74117923704fab86f0bf6715d3ba47de8d8cd7ed314ab90ba69bfba279fd3ac20158a2db39f018e0f9f28f8a0dda0b165ee83fe084f918c7fbdfe1558ef07f8b867b6696c65fc6f306b5de71e3a7355b4cf8d4cf1e80ad213746110eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9a42188ee805c17b666843dc0bd2ccc40f1720bb86c6cdda4fa2c79f557f94acb690cb74897c6c3801483b9ba2052173e17d809d915ed2a1fc620c7183280163bfb8654a8cf1ca5cc89445bf8bc2561115a356df2b29e9ac4823ddba02d0cf98652081264d41f767004a44503eb326722d5136f509febdfe72604c8a9caebbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d8b1a647aacbf1dfed2546282ce0e9d81dbf0229e9c420d95709d20c1b0616b582f3aeb560b061d7f1e4759a5a3e7082ef6e2ad667ec7ab8187fa784fe70d7d8c0bc4e35a6a8ff321e486920d6a71ee3925620352b1a6594eb54afd98250101d9404b43bafa13ddb99f68d2233ae59e3ae69bff6401330d36246b899acd78ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb583385a4d419411be7a12eb4876016bce095cf5d2fac973484f29abc092af728ae6b1486f6c02faab23dd3ede65618055bf8c41d2592f668abb8aa7fcadb30559233412d8d58c613bd09ea7b5feb4916583c8a61e29c2674fbcc92f5d2c502f2f5520ec2532237aef046886348d68c70c08c448d9ac262156661331b57c1ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2905db8c8052f303a12ec718635e253476debb6b86515cfb433936587ffc7cd78cda239bb2c73c58801381d8e0b223a97584e525b1c4d61b0e0ba0b6388b8c8b37ab12d32fcbd64990b8635b871412152a1032650b4c5860e2846238650f999c8e7cc9181a97773607b55bb90b3cc1340dfa5ca76713584a37df891e6e09fcc5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd17d6b54fc2ef0c2632d2dce300588baeea8eea11993cdbc01252cea91acabc5bb74501653c3539ad316d7b49bb6a590eeddda5f72f25122dd2ebf2ac76bc30b233efc420c65802f38318203070acfbe1e5c903c643019b32fbbd2ca089cf2423b69b5551a4909bc0b0916169279cdfeb44c61539f20a155855492cf89b245c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f9a167cff871dd6bbed04de755fc55ac8114d54ef34a445489726fb702e9a942b95a5707d07fae8b2a467153c0f6c9c2af9e99434aaf8f1aafc0a62b22f76074f74f8901ad93a75dd68efb73f7eb6c82419b3331e38c5dba72302b928726b6c668942e2d164547d55f5563e317668be98870643224c77ba5be8ebbee1bdc367;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e65df8bfce4fff8e8a21b969c5b82a9c411ee18847b4b2fc78d25f7896cbb450e9d30fa82f1a8e1b4d09e960be6b2326e8419968e2d1263f8164b8de0bb9688b99d89d810ed9f3cc4bbf898c550bd02e3062868768cae81de067bcf81c8179022c711541c432e678eb37100137b04c306183cddbacc9fb2e8d1125a3a30f317;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h766608b1bc6d2d2c89faacc0554549af9da0b1bdee2818d1ed5bd54b23dafe9af2f95dbbd644d60299854b4ddb588d26ffae6faa780ad2c18f94c024885db7d1cd53cda42bfda0b9046fe18b0eaeb419323b54e3e9446c8405c2dcc795c3e00336c80381285b15e8fa9c734a8f0df46ba833b344233420c6e1b6ab41af263e91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed83fd16bcc9d96caea97e1cf4c2b574ba014ddf89a62b8a2d570b380fdf4ab08b5bc8e7cd66b8ea33227d47ac1063a7c10baff39eb2bf177d981177bc5b8b2def4e2c118fa91365950cca779d95a6e5170c8cfebd750735c5e47a9b8046702dc52f637abf81435c8978123018dd304bc7ac69f18e0f5d9075e89dee582c59ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8033cfd6d130f9b43b5391a2e48167cd9303031003c1096e309164e21d83a11ee016d1013e3ece23298f60221c395d4c23828a473f3499d38b938f4cfc5ced72f75b334f1ecf19868ecc84fd8eaab09c714a77ec87d1324942cfc58fae9b6047b209ce587c58dbe2786102d6d042c2dcc407f212e826ba34b2b4ce52f41988d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19c399310172787ae96e1df94e23cb47a08bf0f03b7c84e62313bbccc44f65571badc725a6808dc94e1a54c75f116ef8209fd9acbcead6d043dbeb4e929a7e77183022e5b059fe69ae94a3228a084f1158c0c57b544403446e9840cab23cf0779afa64c94d70eb870f4794817fba9371383548f2a55de2a2520678b2f36ae12b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79e74986dff951265c5af91c034a070152c3308225a4770b4bf231d78109532095e35a93554be30df3f649d44bff4cf15393f81dbea43e4e38d007c72a1ea5740760557ae0ff3f4bbcbb8b197e0f98b601685f82c70afc88863dbdf7817fed87c8a4f30b1fcf0eb5899de0a4682fa038230ba0734cba8bcd451effaca071bbaa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8af356d13570e8ba83517b9b20051fe66ccdb0ef46b08ff4cd847f0210d8f8e9918178b50df96ca4f6d8a37d3425f3cb3b3febd43ad4795ee811014ee0f87aff06087494880f7d2e87ebeb749d859fcfd34bf5936a2bc31fd6d5c44626843c28f59464774c87893f2e816495ef3013240ec0714bc91607a11716f085a74a604d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3414c75073eaaf6e9c59d6d6ae351fa9b434a369cea682c4ebc178ffe529da2ecc4b35ec006192f7cb318aa8e6b72899ad479038a69d2b06b44cbacd40b6abeab4303a3dc6bdedfd48b42f0abf4aa6e4c7a21cb41f7d5f8fe560467ce46714ebd00164d6d52d3c758672a87cdf0a06f31e580b787bc32d3023193f923b2c31e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9929dc3de4f2aaf3d020738e3ff97ac61bf95ea4e35cd54c32d4284baa9af927efe63a58f60cb242b5380c51dc85da04c117217b3392902e5f86d00e4f140538bb52981e41b15f2e260aab894659088ae650fcf203d9f1ca2ea0549ad76bb51b47caa015c6e8118185589ddcd2578865f33be89c764024d53bdeb240ce97b1b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd529832755afa2fc05c36e1efdf898030c3bea263e8aa7f77dcf6bb3e4af2abf79b4860426742b4a28985f7aa066a3e7cfa07a309e3797adce09d7f5f1ffdefa676b8551843d5ffa5789ca5337bf05df42f7db4f05a6338441517f118962d08429e380bd41c784c2276cd361cb228f8bfbf6c713d62e9988f128d0808669dfaa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h244d85fe2ce6eaafdb8bf27e809f9361060164d909248d2ca15f739bdf4070f2c17db784863df4e1aa4c017a500b28153cbff526c5cf020eeac7bd0d67a7deca5ae5ad55295e83aea48e77df729ceaa226312d8e567697ff6f36623177d69de09450b8a8da10408ba4180d78d18387ad05b28592907de35ced17da9eabfe3b3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f0256d9decd8665f11a95169cad617981666965affff05da8126bdfacfcd5282e1801b0528933127cc46b3bda5956b360a1afce2f2c635f2d2c9cde8ef90c19887d17cc2a473df98db0623d3bcd9abbcc13bb65f3a140cf3c69c927772d9d3d99176bb0f8e2f8be5632a7f132b38d00d6e165b55a5f4e9db40a4515715e8f3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4311480f1a65ef4e8a9e7a19c10eb78558e25e944374813e555c3db5139bc32fdcce4ac9744cc62fc7a312fafc846133a8ae1559223add2ec2525d04573594c3c6325a6339ed5bca5e135ab17271240ac9bc809bb865d355972b600204ba40c18b6ac0255643bd65e54336fc85cd20dce6ebb5f22c425bc4cac9f428a419798c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37a5b55a1640a82b11ab4a927d83d1864dd5cd011e5bacbc975c1ebc5841333dc4cc4aae36f7e2193539c97627d0395cdc37ddf01780fecfba89dfc87380142da3a9d79fb4db0b2d92770ddc7ff66028777eab00cb2872b1c220a6b7987db64c70c6194629fb678e83249423b74d85dcffc862a3dcc3aeccdee6ef6a891be98c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2157b46ebc73da6cce12f1269df8b1af5fd27cd8d49f31b41c09110390edf08fe2fc40ed5cde00c10bbbddbf6b0ca9a86d0e6ef9ee32b539b18b10f9abb4de66eb0b9e385224f9de2e414688e947f7722a5d28beb946933fdd100fa955bd5cb307c06603d60b7fe8af9a387228436b5ed5506587f9f906c2782b0d925c3aade3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b4adbfe170379a65274e04c5d686e06b703a5a9ae316b6f070bc7644c43a121d4bacf3f3d6b346ec79816abc60d3810c58d57a78f4b27a09c9ecb344127ba89d5d27011d12119158a80352f7c042ecc6e33ccb6eeeabae5421baae9090528e774c984a09c6f7aa936664b6c9a4f06f81416fa2445458ae3fda80b331d69c69f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d2d10f469b54ae61fb4b40a91e7eadc7b88655f64b57796ea4115ab92d0211253d8178a7f637cc34b75436a214f2eabe2c5a27edd04229212d07572d8a8c6bfbf662fde00098491f35c097e4e6b4ce491e24d460c885d6070247baed4547610c9b10e3ddb8d28c327844b5cc71c378d9c40edfea367550feed5c5b83d24ff3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc862f38e7d7fcdfa053e834ded88d48ba804b5ab2226541f396f5c90fef19839ce095ccecdf6a31444361d552e8591b93c790192a004f748e292c2bbec1a080123c2ebd3d0df313bf5b16975765aeff2f2e3e0b4b0e01312942e767633af79563584d9252509019b156832e90f9db820654773fbe7826bbc137fe1f9a9a52a15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a6f3bcc8fc6a8b92df504bd52226cb2f898538995097c92bf0075a01ce91ab0ca6bbba4dff01f72274d9ab33f2450c1a9ba3db7080252ccfbdfa62c613d5af994894f83527f89a53db45df13f2e2176ef93f0d097c751daf5e9cea6f36e23a25305c0f6144cd9605c4ce7fa6d067f4c9404ebe76086258a8acfc14a923feedd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha213205729ff9a0b5fa05ac6c8620454f26db79f2d6960212e20271d94399d215be214090e6d6662334690b06f98f6d1d71c39e1f616fb9120eaa8c5a87f7442a4f00c6aec816585ba7d08b6724dcd531c746d62ae9ab182de040c480a8992d08d7f4d46af3c9697262c22cd008105921ab2b57d4bb34b5693f5a3fdaa2065a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf77cd0450b5e0c0913de0cee6f18bdff0baa5544af781f290fac9399bee45cc088a4faeaaadedabef0b20ac8c0bc43de387febc56615050e6dfc2bbd757476220e55275b2be2f61472534c90bd6d443a864c3e38c3cf00a6f8ebb55fdb550c9534703d72974702416b0a0946ec3b4f06a556330960e895a096105639dcb2550;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h118fccc5dc6157d0d77604e6a1e272252b6d81817144639f228a5f413e8257e0c928c47eb98422efc29a1640187f2e1820d5baab6419a3fe4a93f1300fa000a282ef590dfbb5f0eec309c457060dec977e0fe7c0cbeb210b37fad8468903df491f5027a81073ace58d3fbe6ce9fb67712f27f17ecdb17976075b87525fc2d0a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcbd4a14bd226681647fce8467862d5a9b77e4ce0129a35f99f086b33a9abfb0c72204f931f04a9c2fa6bebb776641612befcba7ad574703a7e5356fc7b130d3359128c12bb143f4800f22742e78ce6b9df85abc9bfdc4283e4fbd4cdfc9d82651728de86d59b00e4c0a60c4d612df10ea180ff8f459a65040ca913f35c990eca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h465f9c7d93958108ec92572def9a731267c3c10dbdc82726276e3e6b491e1c4855bb092d5f0817ca59470530c66c311f2350440661b1baf6b50bdae0a037ba72b1ba8ec729ab4573e344e0a5bec577129f46c54a562360dae783537821bad1e16281af529f1198080738fefebfef57afc1048e87f1091a9533db275c6473325b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18e05a61568fc690f91acd554c70d812f62ff5812458ac888b86f4b6a6b5be3668de464873a5088915c6f482cd79c886ca79e6acd49d0eda22c1b8e80ac7196e76028b88490fd6d3182c695f8510fc1c6f182b0de0470453e2625bb87aebdef9eaa40584385aea1fc134c238a89a2710d72fc43c553675648cfa4d64b1446f15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha77aa548ed145c0eb31c94f63e92faae2f38569676203c5dc44052db385adc04264d3a114749fe33f969843a09ce3a4e4be4be50eb261888b8087384598da7df52dcf9d6efcc88e7436f113bc9c8411a0da0d9d40d33e5d1e66432513bb2e58ad85cb8cf75ed68529e889bcda184dd33860a4f7f5dda94f21fe3ad6b17660498;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22fdd1d347c01fe4bdc7146495a004e94f6df7279066f52363d21d76af950c19068c950320753d457b69652c7bd011a6735f4af3c38383df7ed87d76041b9afcbb8bae6e7ed069a0d1d9f051fb8281a42a41af5c0db1eac35da80b28ec87190784c8390935dd03eeb594fb2829ad164c550ce7b429139a037e50a3624c21a3af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1eb7580e1a4aa90da68db85a169bee80ea1fbeb68c6a69d5db3df9884b658dff6f23fb8ca966020862c36c6c323c8001fbdec6f2bb6035fc8a08c9d3abd429ed900f8f64e1f9a88c038a9cc36b7ea32c2098f57498ae7f065fb1b9be1c38720c8b40f25a404b83a4ac7c7c423eefa9458cfc8df97806a91a35226d1736d9d1e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1094bf556970f6e9d136ab5e9f86250ef510291e032c26d3c40889f169a1816240fe0f6386c8d79757d84d46aa011d9aec528a59b8db565068894b40128692b62a09ecb3f79f3ec9d9e4b93346cc9cadd4279e3c777caf1a77f2a208d4a55d39d5ca7bdfe707798dd70b39030c61f84769e06c5b92398780e36116289db14a51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46cb0a900b22e6409f12104f682628925f576fd3c0fc1dca63f2db73c5d7d3e3435d8582705f01af31ab354c8c91058c1a15c2fe745d7eb60b5a70f35321aa15c6992b7fd56e55d537724130cda3fc8ce9f3219626a484bf130ff0e133373ff1bb6f0d4d19b65195a3c9e1eb1e509cbf239cde25d0f0ff3ddb7b16d06e2f935f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57e0c0e6e9ef78d53e2bdb51bfb040e4eb11b5227a5ea914bd7a870403e3e0ba69e9dbbcbc6d92adadd47bae8b289a7b504246d660345b988e86b4a92f460e29fefca26a08389a40b09c50516e0d4e8019cd40dea22636905f46cadc3f25bb9cff47ecdaea2f8069d5c9f7a50ccca457a62787e85c0be38a5d70e91c1ced1c71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68374075b990213fa739c5731b58d2bf4976c22c31d26f01ae47f0cd2f48ccdd8b4c36aed8f5d5b2f749810326f1a36ba4c1cd583ae8ae3815889342617eeab26326fdb037c466f7cebf247ea72862d5faab96e8b8d86f9bb0d9049df92a517eaf15fa20f8b8e05287f829fed4a88b533eadeb1ba4d14565888c87a1d548a1ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67c9772e46ec5a4d6089a20b184d5b4c34666ad21b9c421aec5d1d5e94f9c0e4a6bad386468b4ad96cf5472d0684f17c4aafbc0ea4553a9da86201ce3e9a59befeafb072cb2f8c6707da08697f0f313d3f68f65f3e1e8777680b7cd8ed8bbeae2a85587bac19d4a4a75439bff35cfa980f19e0b09cfe3b1179da2820cf753072;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc107edb792c32a1a6227b9e051edad24a49ca175490d4948313c744ee2706a79748f1d778432b81807c3416bbf9b0a7cf4f73879a4e601b4931dcb1738f61e6e5e68df0e01ac81c7a9ac9e40ce4049232503d54d8eeb1846791ccd6340363248944d098a45f34d96ac43724ca25cc71e65024787ecad98b3a13918ad0b84ba97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf7b4ebbb1004dba014398bd5b951b04cd15d4fdc6ddeee335d86566cc1cb64611a60d4cf594c5fb454ad1b2df77f536a23ce5e7276896acbe3af6de0292a0188a563f638454b2274c093b2bcd037717005c48471be3cdc1c719c07718f5d544568d7d0bb6c485354d1435aa467c9aeb5b5815c980325fb1bd7046e1dd88781e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee513bb6fe80e98c2f61b68317df2307e57ebe8f356e1200f3a10f50bdf1eadfc61a60f88ed604e4c64ef72206799cf628ac1185ca79fa7aadc87237313dc430a41b3fe0e30a0a95155b5e84ed37fae55386a1c734114b8bfdefc9e43da617c6a56f84a9b8cf6f3db0655f3349264643a8c195b45ee4554c2e9ce6d161a81b7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf08494d099571b85cb3d3e7bd07cd17e1b2e15f8dc321eeb221a09a01e9208e6fe9da399f771bedaaf8d7326a397869bccb516a2326b4407e858a5a74e94f80b5ae67b8af3897a00a0356d309aa0c12742e161f31c5463d0c3b8d32e9ab9596a7c9c5a29d26bb524d906918048336f4527edff0f9564d488e9dd4ca23d892136;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1749c92edf5bfa4fbaf9f5ae545877ea8d4fcbccdd2169b8d23aaeb7a0882dea1af4bba5aa397ce7090f619015d48b06ae27da2e38926946d40aeecf4fdb0d446c40b0e0ea481b3e5c123888cf2809d8b592f3e2f854b329074ea2bbf8a8585ca76d4a2bab087264399673f8a20f403df5436b2254049ddd6ed08571dba4a7bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7df22ec9b406a38d1541b42251719e899f8b55f4f8ecdcb546adf6c1fe00467ce4eedaf5480d80937ebf47744b2ba7bf28f5c9a631c4b98421b904814dc5d2289ad4b5f51acde6d173b1787ba8500e1899c5988597612466728f0dd3b5e130f7341469c9fd6c4a5f2dcaa9ac3a270b2385660e0cb4fd45fe30d77d11a225b90b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbd5202af53f22627da37260f12b7fbaa56ad272462de24089691c64bb5938265d570767858a9e83b9e2a4383a6b393d67851d4a17d25b82148c176a39ac9ad33790b08d85b6d5ba296eb76809ae6344eb53b5e939c2c476c4eb334ea90b2fdf19979da0c465702f2f6e40fc65a016951133c26c26ac4c587c6c31112613e988;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28796b70e183b526237b462ceca05f265483793c56a11941f4664fb78dca292e4b07c2df5a025486e0a0491aab6d5b118ff3043a59a270a4878dff4c7341bcca3f30354e75cb9cf5612c7d7165ab063ea439dc7777266fc01d6ab09d0ee246dc11d417e658b91769c29666a7a672d56329c71aa923efb09c0d1eae8dcca89905;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2e2a11705f08a7c4a9738cb0f8c3dc37369f40633a356899fbdb55de3ea179015556c90a4b42d275248952633fa02c2d99a36edbd691f162e497c5093946f06bdfd48086086e41b7e48d788179e5fc3027a2855a16f8d67348ce58d379351c127e876b0cc121535187671602da92895cf6969c6930bd13c4dbe80d8909d7a9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e143af571d88329d670aa0e0d039dad9506dc45114cff77d2f49df7d46a9c7d85f08fc67bce995bb48c383e878cc85db0acf952ff3053e74336b121dc20a60d0bfdc5b38892a1a99bd8e63c048e91121063775ed268d9fe96a36e60c4e0a591e374e4a64d3299c7ec8fe7c0bfab9eb5360a3c5034ac28b3e6fd6f24927f21bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd65b7524c587d067a88cf95e1651cf6ac9a2063c856b72c4279eba1429800995afcd74db4e3f3def912b808eb9773f9065c151c619a5434797515c5b74a14de8d718ed4d942a95ed85fa67553509960b7582b1cc2c4dd128f3f213bab177798e18e339f7c28f0a058754a14f8c3a02de3d6030c4b5bdebf1975cacdd446cd7e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35cc9c53ad9b21214771d73d012f4b7cf3f46089fa5f6336678d621bbf884a997a993b407b1885383b01a25df64bbe858c95465ec1c35899cca71a5b51b44583b49a06ca9cc45ce8ca0c6d179e846c47200d5dec93e98bd9223d313563c9414e2231eada0b9df7aaf2ee715d5ec2e4048d2e38e28490a27337f6d1260b7c64db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6be9f7a8d9890dc5896085d62dbfb01407456e887ab03166d939d13415a96d1a0ff39e6ff31fa35699cd3581dc219af93b5bc444ea813e9b05db956dc366efa375398b9b733311317b8c29a32bc5dc7bd691f39729def226b79e3e1b77e6ce6d393bb5f43a23771f94f24e0620e363e7b146f23a0a5e06038d7ddb9a3c926a04;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19a238c78025e9f59ef3beb913d23bb85a58e8faa98312db0849f312a46bf0462de0d92075344edf0406ffb4128b46fbf3335a044edfab5c803e7a4328e3549fddb5a1510916ece404aa4f1ff1c693cf601a057f75775b7e441107e9bc73ad3916b9e13beabf9d87016026ede9b5a9c2d7dc355e5f0554a425cde17716f2f4f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90ea9b9c8ae6409339158231854223708ac3b305515b1eb00c43fe182f21dc56419633588e397198856695483698673b921bdfe50b97dc13e1d04268a5f88c1d458aa41254f1178d60bc3c198315ae182e1b0864062862a4a7d6b0024b2e6457463dc476fbb4d1c11dfff64bd7dc621c6f9010dcb96b2926ef748c48f6691720;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc531cb02b11d783fc55520d73f33bdf94af5b10e5a5d99436116175d76f120d71fb8a33cd45da659eda5b7d01d4fdba9e639beebeff5a3378f6a7a01a656ddcb03cbbe6bdde5189b59330b5356204b36d1d77a02fe579193fb0aa5bd5c760f83a04cf0ec9df1a0c9cfd698685f8ac4030103cbe11833a162f230b5a29eea3c83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e1128c890c1be50c96e7647e77ec78cf8f848a9aa27cff2d3a1e4dd92c39b33eea997336f05585a07150be4da1c57562b444997895feb60893e98ddd5c2e565bf29f43d917e5782bab18a702cb9b259128a03f7c5315f1d1a06104b6496fa7f71852d401788bf70f730e090c3ae03150ade146f66452af74e28dcda53b476ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hddc29bfab5efddd2754bb1962da71d585694be832b73227ea27f8525d8715f6a4e672405686c401f0439d3d7fee7b2b285da9f1dc4b142a455c92723ad47c1e5832461892cd086c87c0714612d954ae0094a4020dc106c84931dc6aceca39d563403e20048e789f241f610c842f6f3b8ceced410ecfacf3379e4dca78ec639be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h894c602f0eab7fac30f279cfc0f59ab8d950852e5beffbbef27b7cce3e8908eaa00971f8a3a8a6c1da8c4772c2a12bd2ce6b2f75195f03e04865e6a7d0069f9138ef1cb294006524b985272c22b54d1a5109ec210965f6bb2270e25f06ca02ac4aa71009076739059be019d448574cdc4bf604392a97773f4c0409580d8efed8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fe4a4e3d8699d25bc724d7084c662ec1ae75c2c8721eb9b4ea10e0ded9ec5098a555f365fd80ad9ea0e06fed25e625858e738e5c013f8a9a6a8ee9d843ef09ba410c8ba12fa9d01c5cbc00ad68c155af47b842aae55cbe1b424ad7ea39ba8a4db2aacda2fbf10ac5d79b70c6161604c579d8a90d97ce9fb96dc7a4ca76afcab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d911d835d00c3abdc97e0ffdf4f612350fc7fab579cc01e2d370693cd216454efa9f3e5c3eb3e758765800c62e7976c745703009e8c32984d02af06dcadd509634bc8f3f72170538f8bc51dfaaae755802b11f903ab58be4e4caac66b8a5d735a20720a22e621b787cc6a0fa7a890ca064388c8c314e032617594b06327a724;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37307ba1682ccb91025b91b970c76a37f767528d5cf27e6b7716c98a16c55d26fd83f2705bc37b8634fccd4ca0f3f8e4af34b434c90df0473632780610b1c9028774c99ba4149e38b2d2f78a28cd4614abdbada8985601b0a9d52b4f063eaf1c11d934f8e563e909ac345b50a0236624f74225dad5183519f3fcf7198665428b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h328c593033388b6b6616786124baf669947d8479bb97be3f9ac05d30aa435c4c802bc3a3c42eb5f49ee0d96c36cb51fc52c8e4dfb2e90e1ac58b3efb2f45f5ecf484a4bf565bc2daf092f09476829c413e861b9040c30845c696277346af537bc06be4413728813f9f5cdc2f936fecc201a5b4757b11cdc7423d4f70a756d160;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7822b54feed619f04242abbbeaff7749d63ad29160ec5363fdce0b4a0ac38b8fb92f08e74158a8955e48727f80513ed294add87070cd40eb5689fd4d0e26b43c59b8564d61dde7ac66a15c7bc83fe647b701c7a42b24630e9a4184fd3b38adad26512c57da0ca7a2bd27109093101a1d306f7c17efab039d67e3c96ecd305655;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd40fdd3a6dbe2b5044929c82e6becf7dadbb3692f2e3a91abccf11b449ac0cfb83fbcfdd09e6727830becdc7c87c93cd96315f99bdbf2d0bc7e4734a7edd4e23ae280ba59b75d11949f0ff76116943dd7f7fa110208fd3bf131e32b244c67d1595f53b6606378dab6c56bbc5892349eb0be1c76822d122ace41227e70f0c8e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1111abe93de76c005f9a729c19667ee40e0ac46ab7dea2e16bf9891286836ed94fddf4c9bebf1936faeb1fee6778008b9f573cbb1897d4bc975465920ae5ae9e0cf082cdc0ab2a85a0a6c3a6db6886ff69e42fbad1d24a15ac84bfbe2ff934fa092047c41dacd8d64671211542a6b0b040914b2cb10bc747864357b89e1939a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2294e55cfe6f80af36ec7f5d898e1eaced6c18af46c2b079d053afbe821213eb3b805b4bdaed554a20fab2b730de0e7a8055629a85381d9b4d71b3ea490ec02ab0b5983b8e06edf582099f767570d18d1caad565c5a65307614ec7659539462da819211b97fa1ab63153b692287bf59ad1230db05cf80bdb433600562303955e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f437dd034bdab282c0fe50c816962f06f8c4b541f16ed4aee73f8f0d8ae9598acb7bb76ff1f78152120f309e611a9c4c578946a699a3a11603746c8f0e3108b319326ff116457550a741d34d7684ef58222901a7e7a44870c1d4246f0fbbd868efb8d4dee67679539265c13c7cc169357b71311314e8f6d84c7dffea6375d6f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b8aa47cee53540318a19b5bd849bf5ba788e4bbd278101664e63b992046c354aa5ecdbaba7d649a0e0156224a103a0500528cf3d153258f3d98d576db8d27fa3765f04c58cf23e279003ae111750a19d0035fe0d44eb9dfd3b9f70375af1b089c66861c84c052ce26ed27704d69748e244a636da42d1deb1bb8b3262556b1f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19effa3ec4249eabbd03dfad0e55a38abe9af22e8d168dac3aaef19e5220a643d6bbb0a7b6ca98a609bea3ec989c69f6960ed93651037a534d7ea582e4a4f286520bab16698fb1157cad972fa768703d84c243ccfbee7782042ceb19c52992d6b879354c1f887c8b1173f48e8271325dcd45dca6aee57a1e314b8c7ef1a3eb93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcf0034a331da5786bc047de37edf5a8b728cab4e06289620bf4743f4cb26d00f56f0f77a2c1811e9d4d775dd7a0a19d518855f05930a0b4d6dfda2ce5347149170891fdad9847750359743e6793cbb14e04e29e3e104a087ac970f1f3a2dcd52957fc2cbaee27d264d6d42d7cd3fd111df40dd830c4e5109d392b37f951ee09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd56b95095ab39c735911a6cda3e71c7016326e3384d979e8cee6123f48ebbe331d78f0f175ee1a5a2feb57c66502159c2581927756d21463de0745fc99d7177988d9b1d6adb958ec57c0c292ce6b9923b911365ccda43d1bf2e6a6904ee0956acdd662ee7eab9e3c24aa74d8cf01bf5d0d00952f04cf0da1378294cf3ba4c071;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa67fb68da344d31b0334642df19dce9528cbeca1b8b1c2483fdb7fa7c1045c333cefd77bc2afe8d309ca31ddd79140a2fa656d9f7c6d0db878092582b6dfdfbcfa804561081e97e3d065d59cce09ebf8078d3f615cd93f6d967b2fd050d935542fec4bd7fde01a48a80c33aaf58e7b443d6e4c5b9c8f4c50bbeddf89718d88d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58e7e665d27f7978d6a861d4082624d8bb2721e898727f771cafa7a9e5fdf7dbe58a52adf14a2ec97e0a9709902145e8f272ecb0b36e61e1a5325359cb705a30b59b8d1dee28ab47f6f9d7e21ffecd5c4aeaf31df7095ba033987168d22205c17fc72c6e5f5e9d4a8ec013f93bd4b2c61c6b86a823a8a70a05270784f3be0b16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9af1bb3e79db762e641f7c7b69aee613c48b2233a1f60d5e4d753ae9291af3e78a70b2b73754b4ce9f654d8d81b100c702718e411a7f86891b5913715c444373a881fe47389097f64befe061ace9c96ca9d19a2604c4814cfa3c7985b0cf3b1b1b0b82de7723f95e48f6e71ffdf5d1e178c981c6952e36cac4320906c22d6722;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc0bd2e39c76cebd9b7394a742ddd0fd0fe303b27789081dda4dcfa8724aabc92910442abc0cfdf031f5f54fca0017a2bc44bc0fa6d2ea3eee8fa4705e71f2cd667b916a7084a7049e8138a6be4fe99ae1050260147d3d5e1180a57364734d61f57e5f98c9bb8c32ca50e34595bce4200fe07cd4a1fcc71126d0c996870dc3fe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c0da9b858cbd68a9642ff546541a590257d9c5d869f9e69678954f8886a59be1017129e4dd69ebe04a2a12f449d64f621f17da4118544286bbac364af1549bb1a6a38bb5bf302456fdf156808ce0cd2bbdd91dec4f541d51be96997efb7978ab905d32539cbdc10638e29417530600dadc8e67aa5c627b508b24d051722fb69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34857bd62aa0dca9f7ab25f095e265e9768c4bc490a03f837c5d1f15ea5c9b7060090aa4518533da238ec888b0555ae51096509d59ae9593a80ac42888b5c64633aec0469908ecac59ea35e82f34d71981de130985d081b038210b1eeef66b966aa6ed780b5e98b951450df4a9eb10bf82f473b878bee40c9a4c70e7872d266e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5dc86e36b388469c4dfeae920603eeddcaadfa6b28a1ce14bced23d8f646807226082d3854eb4a6ae0c44abccfb529dbef9af5c747760a6056d9e0204d228720ba23750f1507af0bf9171210adc186713d497d41f30cf4cce10c157bde6d46f3278c277aa251a76ef589ce20e79ec1cb97ddf74ff1d8bcf98334fa9dfe86cd24;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had84ec8a81d1908534b82bddc9d32a82e64473c351c2d12ee1c23ab00485f2ac3c0c3757e003cb68ed0b071b4c3a4ba79f65d61c46b9f7b513c807ebe8a37c97d246e9022a96ca8e2ca3839567e07749741e92d6dbd02e4596d8cd51257ddea259c4f41dd0f68a2589bffd1f8293fb2a918d604348dcb057503d67d43a28658c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1878d3cd4476d54f4e56538cc5d323c2a07ddbb9e6b656fc95b7162462e66501708ee338b56e88999f84939d0b949bd8c529d4ea753570a8e7fc985016cda35962dcc430b7fd0791916c9ef24922e4be696a0aec310b16ec3ef9c2aec57a571db7bd1ceb3c94a9f3a82fc6cbb6fe53a516b588a58eeb5aedc23bf29998ee2a7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4aefdbb4917837c2f9a02f799cd748a8ab003068630e5a62beb887ea67fdd09e720ea3da7dc11298e3364053eec2dd969511833ae9af7395e00e1b8c09a1703e7b8aab37e07a43d8f4b2597f619860c957ae3c4b234a995cc2a9fef0d865c0ee1ec7efc472ae74691278ae238f4c5dd5b0f9360be8e7253b5dc199e3259ca1ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb30f1d72c413f58992e0a40e95237c7897d20130ffbc9ac8d64710ad9fd6e57b0e3dc794782af8d8cf7034df7ce61c9f64079ff48a8a07eed69e9fdd005b6a264a50526253b0231478bf22e54cf66a3089d5f1a30199e25862cd013c157acb6c75a5a256953af25ee4275ad4e1d74326bacf37c6992971c429d04bd3cfcf014;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71f319ee37af0e9db06f893ce77a4693ebbda9b6755ab88d145e8f56a566c53901d70907aed3c308f30135d60650c5afe1bb15dfc22ad55bc2ba45e307b5cf13a48903e1210c8401902d2eef21654482b8879c9ce62f0366f11f314ada8db25f189fdb862ffdd47d0f1050a646a425b2195d51612822dc4a01e898eee75a54e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf17c15e8dec75f883df047c0802e9b58dfd8a1f1f85fb349e83152d6bed23d617bb9a21c8cf6c61b55de01816994e09d360b2fc5bcd398de2f4730da290967e2eadd45f2afcbbb064cb662a2d38920f3d2a9692a2924b02231e2465f8bce4fc0ab8efe9bc2a86a448be7b9a390d41d11b79724511e9faf2cd8fb7120c760e64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8828de232b12cb831d000d93bc45eaf5b6ecc491c0bc009b05ba48b4a759b21ae687f33394001769fb1674d6dd14a1414168e49b6dca25bd56a475c60c4a9603966a3798b706e3419238bbcc35cb981e33870d0495439056c068159517b8355f73f04a23c0668762d5f60bfd64ef3ca36cb9bfe8488c940628664c6fbf20c2e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec8466ef637495edc0cb6d6555ec3e9e6530de976a99c5669795bddf93fa704af24179701592e9a203bd9fefe6fc71452ee93b6e72e807775301c8d42bb8026074c575a347fa1d2db119038c4e7ecd7653ba4322b4b005bf86b2c770695d7dc8cbed79c6551804bc91c9f197ad4d325788e9b8b45e2c5bb1a6d8261302d63053;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa39501dede2fef2636c207c486f5768ab8a55d09facc7d84de230ec433cbfc9db76538ccdda3b03a95b901c36c5c1b0cc63f3b76fff385e4c7ef9988dd092af20c6f166b24f5fc323e7db2260179456586eacb94941a3ba33eca5cf1551f9fc2394af3a79f1752e1fe1b7f18da77ccc9254041320a9dc49c3a4edc377d24815;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfd2d6d83f0f1d37d5b3d5027a2abf1640e967c0b7295432a3c247266c4a2669b3c99a55dd08ffa8d7b359925295a768d8f06ea322b2bf635da664f73f0c382e137853064c994ca4586793fe57a9149ad628a1fc1232fe3b55ab2f6ad64cdd90cc501e422b9c29bbebcdf591e485a5576c977eb0ea467106736c9dd854d6aab0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95f5f53eecbad9a69e06b62d66933dce07d7907e9e161b34987c2b7acdeb747059b82b2481d9ffdcd7aee28038b093d15060351e95e3ecb9efda9caa4616d253e3078350e9d644248785dec56373dff992170fcdc6f0efd02c2c37236486efc4276f95f7bbaede2aa177820720010d4cc387a07b4787c8ae9f4ab073360c8844;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4d3e44da88f556d56a8a1785422e5fa141663fe9b07ba800cfb51d0c46d7e4c984cd061131239626bccb3a93ba1e2da94d7bcb6d02b797833ae3987bccc9694acd5670af64f24daaff99226de149194a93868d5fac6affe095031c960b0fdddafa4bac41e7e2f149885ad4ebd692b32dfa1c1aa24cd43c55737a6d90ec796f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d77e9a3164ecda4ecd447bf052d5038decc7db65c41a684d185d223af44aa0626758fd20a66b155dce584b66a58d3256405f240cc0b2ef97863f60aee4915f49304b3502ce81a5945a346729e01999254d280aa167fa1f039a669aa34afa202e0b65130428ee74433186633f94384d479585dd4473f40643f517eb2716a777a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5772fe7bc40363c398f49b8bcac21bd71bd5e8ae0dcbeeee9a916c463c59661d1396bf66f7b96786d2e740bf2be4c8a37e98359099a5328e5d75db86431da0e40534e2625fecf2fa4d17797be74931cc7dd6e893b5ec79eaf0231153dd868ec11acafbb6ef913f145642261a992431a4a1cbfd65c521eeba8f2f06ebf7431f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a2c3bdc6e4b14852c33115f21ae9834f80be50c97059824d94b913b31dc6a1423f7dc199415e81dd78a256ee607da9f8769d4f0e2ab8176bacea0a982899fc2e40103f17792980fb1a8beec3d5c0510d60e21d5d59cb349f95e94dcb6b03741e35ed0412213e2707fa9ea4708ef226f7734e8d8fdb36955284e7f5eec3ac0d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffe8954ec45f7ee7cef8d583ed3ad15ceede04875895b550f76e325abd8b443f356b03047ef1509926f9fb799064057e6069365126633829cf9c8eff3dedad9425339f1e15aa6eb0d9e59dba36596ece536c080c9634bf2c7bdc1b5d51d800caabf6bc78a0ede80b924cf0c8697cd5997fe6fd0d835d5254235df28968f0f5d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97436db8d539fcbe1bca32c0dd48891f323c623765f96eb8061f352d2e96863cf5f31da9de8887441da91d96b9be0395456b94342401459756c640b54229c9f2cdd12c1a6238ab2fe0ee5ee2acd96c3812565c147bd8d5edce7e99afd93ed0a7be2df164221171d6ea6c6a192a0f5fd2a0c3e903035e67c7142db3a59216cb27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde8dc1881ab5926d3be631266e1922cd1b788ebfd54f1d807ae1b9ddeab04fcc8d57c411624d3c34d6a582972ccf17d688bf421dc356e509ab6ecf1fa86867b6b9e863e60e278d4f73e95e7fac88d65971416caacfee9442764a103e48bbf391b80749d8e13284368f13435d19154d4e858d957659f4a71a27b780738821406c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he201034e10398313df3bf54ec999f8f7bc5e66cabdd43cc148b25bd536794fbae8714fd4f89a271fdf9a0e9c7e9d966dd231b1c4a479e35bb2451918a439949f62a03b615cc51ad9e7ff63712796ef20dac02d028fe5f7004e27aa4f06d9ca037d3ecf9ec0f73cb451419da2cb947639edca8d35839e899ccd0666824f37b731;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7f658c6c96a3b58113e4c5a5ad9cd0e2d497d4da1b594056899d05da2abb33e5eb598bb1780572b4c1a717b907567807d4c62019ac31a751998664652c43b54d79beabb7679fc2db364ad3a1845ae278846c0919bf061221f71ef3f26891f5ed721504ba52e222eb0006754ca17031180263ced7ed10ea7e13ef2a1de107f9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44e0426098f3b96e70acdd7cd14316f5b5db9d46ff0b2aa4cfbb9d7b6cb45ab4d70b0b8d62ebdeb1e8efea8179f09bfae92a27a985a341f97cc794234f891e3674dfd8264a9aa640d4559ec3d6d96d618c1d17dfde340d8e532d926ecc1a81c4d812f17ecdac611f3d48caa3772c42946d9236d1f36cb8b70be3e350ff20180;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81d40c75340d52442c6e7a5cc3c259d3115ef15fc1ab08107f9a7d1b96c175afeee77292d2e5180b9adde08ff7195fb4a98a314ebca9376570ef1da5f25c9834eb109dd26a433ce45b5c3eee3f0ad2140ddc12c1fb87bb8491d7045d9f21dfe0a65123b2d28c146a731fb13f091425b069debd238d87f40c6af4f0f952815384;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe2cfe8783e2389de4acb8a655cb44ccd01678003d79035bdb2c9eedd0c64f2c08619b75b3dfd69d216d3fdd00c5311e7f7af7c8c9ad56bfe29819cee7c883fc6a9a8aae6aecff3139a7562464c5b8651af6001d0534d999049c905347ac0190e02e5c037cd332ce3db36466264cfabe49f8d59c2aa91d2c0621afeb3a823181;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d12820ebc1284b642eb4c246c96f7f9d699016e326e52744987e4173a31b624e2e725c6015bf0294c97032a24b9fd2733196741951a2745858617640a9382aab974e30b5d68b3385571dab797dc992ad39029f9ee8f76bae07d1e89582f6340249c6c188e409b5c337eac597b4930b744c2fcb191523cb3b829cf49b44813b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5e5603d6c5c941471434124318a8a40858cb2c5981873e22b509fd2bb09b8123782e8387e85ffa1c39897f27f0ae7227c778d4c7f3bb1fce05e1bab4cad4d71bc30f33f37a7147f011821ecacb1e3b9a34f9b78bc63b77b86bad24c1dba23e5e9a2074e4fb2be9f14290c594264f2ce778dd60681b97997fac7e5c558b3fc3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb41bc82f373af31d838773cd7c900e91306d5d5b4c2b0fe38e9005c625f3d4cd6897bcdd68618fd38f2be7bdae35ceba27d0dc1c047dfd2001e256091fc97bb7bb0bf8e9f8d6660b08e2611fe1669f68a84f57391eea40c7369c320607c18f93ac7db86462f553b8e794d49168bd71a91aba82d720d71d6746e74ee5ae3ea82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he66b4d5ea4a9f4004a53c28aafaf05cc3ddc539cf755c39e2c6bac6e3ee45b46697e4ddb5ce1550e27fe694b4336a8c2ccb63572bdd6b732f0b8cdff98fcd11c6d0d0037edb6e438358c3fec68fe92d47de8af73f034474421a383c1a45b44322eb0155aae7231ecc1ea44a1027cb649f4a8d9bff42324fdc5044c26540cc6ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f464429022dd55b5a6e58ba59ca6885ff1742fdc270b0018b126099d1cbdee3c22e67d27fecd99dbc44e0abca9c9e7f8aaaeba4745553c5b786aa192fec50a95eb9b1c6664d0b8550f58b9e847dfee470315a33a5f8dd64e3f392d4ab67bcc305672bf9222104583905c62d912caa0d8af4654b2212181e9ded44b07250e418;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb8e76c59462eda2cce2673014c3e30986d156a77a85a6173efdcfd7d6bfede8e9a73a21e102e919606dd346201f24eddee6abcd520ad5f9b741ff6647e8fef4bee4cee053fe7db1575e4d9e16824a36488872d2adce1282f6cda139bbe2294c6a7f8a83442fc00ec0533a349774c2abce967e95c0a70febc79627e3d377605a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h270561db984d711f1e0ca6370efdd9ac04f889f05fa6ab2da02c2316409fc959791766681a831bc7b3a0887c67175eaecf0c0a47d45e5691b9c508294227ede87df686bad969c67726202f0d0b742b86adfc1c9ac04d877361d4670c58344203e5486a7de6027322d66050fd2ff4b604007032878ac7f1f58644fb4a6f4b0c2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b1feb7bfc501e842d4bd9735e9dce0f29cc605b2b5e9382a64cad5cb8bfccdad203cef363f966f52a2d21146c592da523a18f365b85cc22e6a971f4dfbee594626500ca1d9c50e4adda506abcd5c69d774488c8fa7a744b74a93355e66e5e1bfc668f8628eead5b498e30a81a492dde366e923a12c4c67d1a0786fa29d96734;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha79f09e4f66a60b9c29dcdce88101b22135c264e73de85dc5643c4c4885258a6243dcb2bd83adb3802497e1b9c26db3c5edc177198595d85ece182bb03a6892154467967b7143aa0e464f0d817b5bc7c786f9f81d24982977de9e08dfcbb6e5ee44bd85b46a93c8cbd49484ad4bd3b3c2d58e7a1d076529f9862f72064558740;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha492d18427511bdc74d59a97a958dbd3376657fff22f2a52bf1432aee077573c58518eca6009f540c285dcf7dc9a62ae438909b63e91b16dd1a8c56289c7a32252371926c40d4d9fafc31c09891142922101ff1288cd100e5b79a38226c85d4faf1b2e6d052356029a31f75b92d7025c6a1c0608bf41fef14e42b34ca2db817a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8cd28b077851351debb423517ccc6e4d8913c1a23fb4b16686e64e8f964fb6ffe81108ba363d873b6eb9307a21500cd1b587d2d87687eb59fe9a5481c0f28fe3d3900de418f9131f813e05d7445dcb0f5719fee516209cbdf3377d1d037fa91555c575ca1c5fbebda5a8cc008c025aa3922c8ac700dffa6639286b98bdecac1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h136c5857336c43dcbb6ab905efafca7faab82b2b949f983f42caec5d9318d8bfebd41f2e80e6cb198d217ac67729eaff66a1bb338227280a7b869a2b24150467ec964a68473d387f7cadee1c6c21ce4764a33d5ab82a2b2aa3347c6a286de369f2a496631cdce8589282ceeda9a69aadcec4e0fce2a92ab8a5dd6e23e9b224a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe0d2218e942e55a85c4d0f525a1b865ba948571d87801c55266c69572f8e559390a33d1b7349ae61bab379848f0fdb99b455a27f7c009b5653fc0604a685b65064fec8a485063edbaeae5e74a52410deea58cc3c63512c90f2e4def6a0814a15af7b7549407762a7b4f3ea85a7df6f0709500deba75c60e10d2d2c92df330a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f24c49f7153c57ab5060049a1a1aa3b07abdee4b0f0aa9461ebe63b8e209457cfb72c2c1d01ddf8d5c126e7c2bf573324c0aeba00c240f462fe87b58e9a40a15ce0d6d7dd245f9d2aa880c3eb53d0f38dbc49da96c7b199f9666e18fce0e0f67f08be5e50201436ec5f74d6519fa1b88822436ecc16236235fb0f85edb4b376;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18cbeda463cc6bcb300e9ac9b82430920a2c2529007ba769b4389dfa97440d49dac8240ea162d799353865c0d3738f14b91089a08bdccbbbb571bf1a325fb795ec6454b4b3e91bfc04024ceaaebd002cb2f43b3522a486c2e701c73cf5d59c71184db9d40b9359d89529a1cfef275353c6c661bdda92555468ed342e1b547233;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88ba11b545da29017033e5e843e30177c4a1bd1e95777428307227f8a4102f75520c67889e7cc8ebdc82a9826728cff982b16353e0bcfbf9b24f97c5a793e843eb6eca8273ee0964470f1b615eb073a340b68ed971b9b6d8c6f70ba09e452436cae5f4dd11fbc37fc9640e9b4920f527403d185f2baf766f8dbae387875eba2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd75775c8a9b09e91a0268ba23ffec88c8464a4e3feaef3f4f400ac75a26bb048c2c2871a53071f5a3679a1bd5dfa8e61c02afc597a665b162f98bcf3f24ee7080f02108e6065d8755469e1bdbd9f9f9167ff5a5abcd8a5c75dbc4290629e73765ed39eaeba44f542255d004504b31b68b1ac378a4ec77c1b27e47162a89e871;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h644633bebcfda5fddbd65d3b6d9f29443001f34952f493582b735b38bf5b0a90d44464b59dbeab9fbdfb0ac02d98b232da2ae213ccd184222f7f91db5240600a5b8842e8848b515227833606343c6c64e7bd8a0935eb5d048f89b958b25a5dfb81c48e5f7eee7e41351f69a20f316a6003305ade6afa40938ad018b1c181a2a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8283ce8bf25fffac343f0496d285d751682fe470a3d8e5d0ab7505a18bd1e77285f2d32ef426c424cbaf6d5801e9d33733545cf40e7304aa39a9581c0fb2b08eddf74fa45b42ff5ed2814e7fa662b7d48b7dcee2a3488e066fb9f534000882bb40f568d57b9616f50990455ce4d69a70f13a50b7ed14faeb82d7caca49a9203;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ed37840e9d9a373c98370711d5eb4c6f971f3dca56fa94c9ea3b79f0d74e361dede123e53b72ddc2b81304efd766882d93ec26053c66994f0955cf9fb48f22ea5d0e08cc4c6f257ab59547e7c13e14a2f5ae92a2b2dfae475e14d5e6c74a9cb609b15c5e692d3023750848ce9bd1e9c4d0332148b02da30d89fa61dfb5f6c3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9eae1de4fbc0a0994647cb5dd3f3647b4f265d206676b93c066b6808378c675bb2a7bff59994e9f9e37714cc8978b6dcbf86baa5ee2e965a99985c2dce759a3933322958d970f0530cff2031e8ba4367f1b1fcbe1e9f76d3c8e0915aa36230c24eacba7f057a0014eac5d891fd612bb4749f25998416e40dcd9e030c7efb0a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffbc3877b86ae7dd60e584734469bbf422764f692c1abde99e107947359034c2248ade02992668d470e30431b6089e673e4d2bae52e3701d237bc7b763745f6f0a148ea2240c1cb49155d31c8782a9a730ff3eb74935a1453f62df92925abe976d5285ac27c558424d5fb92e6c9edcb31b67007f58c1483d22f7e8ad32f6eb2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f33db2d4a2fa28e5f2c956ab73d342c50066b9cebbeb4d486bccc3685bc0570fa46b6e896dae2572c471d81c2a44a3e91a94a2f47e58023b22211ef9b3812f1604d06882a8f1a73bd88c78d3798ff54e7d0dc2bd33788409f705fb0bda466718b137dc9b0dda88d5a65c5195da7ae350586dc79456eee06e486d950913cd9bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73d2c782e2420c5a91140272868f423cd0dfa4424a70f4633962d0e83da5c6e19a613a49345a0c6151b4aa702f0ece4e33743492d7189f4dcb58ffe1e614b58e9f402c6a45bde543c6752890fc944501293bdfd29a138f1a513f60de9126f47848e8a46e240d54c5049eea1dd6c75cda9862652c1a6d92af6d17a30c5fac283a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48073c43446218626fb53eba9100fc09c3d0c4edb28f9133d8cc1b8b25ebd326054843b1fdb1f1a696a30a48d78aa229270e83612e17d3408cfbcab2a18571f6226d97bdd6e03d47d2521cd4d10fb36732b54be84a805d313c06fd4b21464f79773b77a8d95ef7c71caca8eea6ad8ffa5148b6c75c4b244b116e56608235a165;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd35ef4acd5e1ee45e5da6c651b1e2ca52fbd8c8a094b88839b31de3b0bd5154ba2cdef2935265142bac3680124736e4214dc1f8c6938c3dd94fdf9c89d084003f280f83a37ff2477136ed28ef7c112d1cd93328bc569bfddfba3972a351475a59c886977a80c2db08ea9b8b0708092cd09235bebd4ee794c15b48e4301c688d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b7d85aea1e4050862b9d82652f228e4800705719d39aabc65aa7294981575d9441613344189d7617580a773c52974478c5900eb2f9063a92bfcd0cd9f701801e6f8f41207baa148b91da9604ac149e6f0249ba4d1cb958fc0e5fae8d1c7b0896719b9928eb9fc3d11584273f5f803b160f5b4942f4223dbce9207e584b2e994;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd952dbf7deb94e56e4efa0fb3ad1dc5bd11c0f25c1e175c7064db35b56919ceed5a79345e97d3375ac23f97025a16bd4d48ae9d8baceb7b29ebf25d2f02c9d06e319731413ed644d4247ea7bcf016de1ba7dad2af2c382bf6afd2285d1ccf79c28fe06405948aaf20af0e42db0d749750fe6c9ad5f1692a37e50f3e42ddd06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bc5c3c6a3020a2feab33c27a3b3c4c1f010e9efd9225c8cc5fcc65f224b417522ad4b6ed9f22841889ba9521e0460ab222748c5002abc97b4fe17897e168d9e1a86a5dbbebdcaccf2f96e94af92a1c061553fa5ac76b7a6d274db0ce6a34db50e6dfab6c9694be9c929b6370ba83a8a8e8cdfb12d00b40597c9b6fd4007048b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51c48ab8334fa170fd317870b4d7e311ae836149f27f9dace7472726718454c1635d79da72c34c42a36652c4ada0128f95d3d714358be4255486a3fe6cb2869c0d0e4dc5bd3c6f1d4636ede011526c02291656b01195ad7374b7559e369a28c5ffd6857575233d75e4d7002da8795cd40cb43af518d7945c4003c3f5f18d3102;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h474cca2141961ea1ca0998bc2306b0fa0074735cb7d52c8f9c27ae9109993f46fb24b47e6b18fce9f17db0646809ab58de1c988348e33bc262170dde5293bc6bd38e917ca03efc2f5736a88ce52ee40015b8434ff3d6f572d91d099e67dec231ce06664a1d4cace1cf4edc340294319810136a965083256ecf6afc3f4413732c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had3714b89171cbfb9a1ac3907be1a6cf2efd1e7c7e3f0b6d17d157bf8df29649b1be3f98d5745f6c3c4e4a1a7815168ed344e49fc285f46c09a88d39b6363ff9d8600df5a397e1527ed62201fcea839eed1d5a33277b2671d319eaa6028bc0a06e9a8d7a04dc5d4eaf5b8da1fa5dd2b3c44a72562974af0470f5cf28e1db03c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a625553651d434b54d070fd9da3210fa84fb07aaff74ceead4169017747eeccc8be9a878fc57f86c66af32f31a036dfff9d1931d8faa980932100003658c6b7831d841d1d6ff55c5ffbb3edbe3c506e90c0ebcb9154877c8e708297dcb6c2197fad3db78d27f103054ee78e568483d1fb038e5d6a57c7463296273edf8ceda7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1d385b15c0354524094dd0f2b943e698e529b52357238a0fe204fb953043a66e2d40f7f0a63c7e290b04fc27f1363832f9b3ab86aab852a0f2fc138b34ddb7ad12e574f7b468e475d7d5630a6c0ddb543eea85bea8487b4f404f92a7fb8eea9c6b5033b0c9dcab867eb8dac044b56049abfa0b4deb3d2b67702bf2756abd99;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54f751d0ccbeb95a6ceabe9e984091908a9387e00d15f6088233d9ec716b0742b9ad678798a0364e47b969cb4a85a94fd53eb914e604ede531b5d50c02b0150f9992e2ae07d4afcbf06e5239236d868f416197ae69b3370a464b22c7066c5bceaeaea9e4e546a06325fe4b2fcedd8364372ac17c86800971ae9782f9cfe24ef9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a505f0739fcfb3f64901b4829aa6c911028c37209d756a812130252fd0880e362f6904777965d89f7177c5aa081d77dcc8928a01a11b04be7f99330b6b7388dffe03ce92db36d533963be24f8c90d8ef99d7ed55c90df01e49350deae710a67be0e2364ad6d80a8a677340a7482c5e89274f52d7a62e7d76ab5f5d21d630b92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5433edc8278bfb7e9af90780c32ad6354cf17c44004863aeca54283077a498628dca9e341f6ff1328d1498d4a163c246ef623644977d193a42085fbdf343f72cd9c3f8c75168b90e1ee72901f82563c1c8808f6a6ba017393a90103fce6a1d91623da30c1262ce46e99d032fa97acbd8abe2eab2e242b6b43a9b03f0ad84647b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a2383328d5fc6bca00c1dc3b54114a73dc50414f30665b2a75710db9d6270aec59b694187219a1ddec61937c3999155cdca04960b3031eecfbdea89534e15cbc247f6dc951c9ef7c2afd1f5b3eee83e1ad200e7a73c71e0c8e72ea1621a191542030c372423c97e973348f4e2c8eb44d8264a99e4afe6d4310651f0964b502e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h820cfcd6ae12985f55355193844a55c1fd9fb8030bb38d6868c24bef0b4e77b7bd6aee6ed695a4831bd8498a8f884caf732dbfa6d89d60781ab571da88f30b772d6fadb98169bcc4317ab9e824a3bcfc90f23093d627cc1ab2bf9ba3065bf6fd1225e1954f572cf3312ca12187847889afca99f16a54944c8edbb0a1bedba460;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h886e14f6b099f64f8fc32935104fcc1a09e00763891fea0f07acd92f432cc453d687f7e490e79a799825a0c49cdc74408b28fcb56c9bff4340c06aabdbfa42190f7aaef4fcadf3509a3a50c6d1bd4f5f79cfb67492ff9e7dbca13f25f0f059211e6bcb64a4d2995885237ef8ce8ac62d367dc6f5197542af49b1ef5d336a1a70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4244732f86362310a3369c400cf977429926b083a0060953c53817d1756856eb1a672ac6c8b4ff419d9f7502813864185f76e1469ff093e13b77ebbc26e9cbe3d63eb7d064d1a1971f14abaf042d829b673b2280e975ce34c2ea5aa184e0aa9e7b80b7ded1eda7da2aa142c51cb8388febecb87e3f9c71a781ea96a77798244;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h850c3ae2f0a9724857723a1b07000d671767ed0673dbc8ed7928dc69ba9fca09f781d220de16e960b450f2a8eacbb8e3360ace74df27116c0b8e697be0ea238f6383216bfeed79881bb3002bd2809e52e467416adcfc62bf2c807a5f4fa6099bec7cc833e1efce2c657004247f1d0a628280c1f466ca17e668d2a23b66fc47e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee84ceaba61d1bc5a2e70a3836200458e37b20bb166a8023c0c9793ade3f33819eade92f528a9252914fd5401e1f713a2e20576ec0e72e814a87624998e0c5580c976383e68552ca79f5422e8bee1b5e3c65bef486c6df3ffc53a4422bdea146f0b9f6985f1fcb5793888d0b73e022b99fd6b8ccd530e67a62509bcd1644fc6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57fd857a54912f52b7b455bb87ba15ee96afd32c6981095529a31d089bd48856246000648e5480a4ebceeb0432a1411581ed7ea58c115f5d894b2853cc3383fc2654d65da9d9a50fd140bca08db2d7aea2b6bab1aa696df2a84d9e550e431c3e81b4cb30e131844744a550e4b4bb609e60daecb1f972349fe78ab570834694b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab379eb0b4e01173eb96cdd4bfc4828f5e8f466bcf80d1da7fc343b3dcd784e0ad134540607011b1f8f329b0eb1a8da7d49c3fd9f4a8a5ed657eaabdfbece37218b3e5ab84a4c14ebe1566ba12f8bca1f5789dcd09ce65abdabac6fbbb3368ee33e87ef475c99c23c407a5d90ff3efc731ff95cb9ce10137a7f2fb81a4d641dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9adb68d44229e23ab715f8d4fa28ec2a2cf4e37eda30c4532b5948739976d78666dd1798be421ab61844f2a6d9963064e448005e924a21ebb6f4834d3e3737b2226b8dded12eaf7edb127d9e073fb308cc6291ef9b3a09ce8baca2015331d4714594658aa6e46cfd2c0758ada481b7ad7af42e9398401934dd5bd6a1b7b4443;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2444d751c8b84244657ed4a45a03d9092e92767da66d0f53cd4427251243ccaead77320d3fc4715fc68cd49d118d6c12e97fa6531e7d91118a2b822ec05dc6fed4f4182677ce7c2e7ebd0899388a41365601988299c4ebf2da581220e2d904218e44362c9c79e3080ec4e5c734ae548e762bd90ac2b6141b5b34021b601dcf8d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0753705e26531bfaa98b0f5b1fe87fe6f893263fc15eadaddae3e7b3af9f3bd8b80fc496e5582856ef9e2b0be342b325831067fbaa2227e84b364f0f81739bbf2d74523674b994ad597e882f8e118d267f43e8c8811165857a506edae83978366c1c629c4483ece87ee92645e48cea0ad3aa835b684ff493df3eb960794c879;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h587147d50161226f04a6d10dca355aa95347529be144f5fa5ba62c5e65093f2f505333cd34a3e2f629aa20c0e126fe9e1c976415b7d092324c3907123a78f2cd3916bfe25ea6c3b685b7602b263b287ec1733532d70e153ecc7e7f3b1ebfcad4f958d62b7fadac372efc58946315aa0009c2023c2fe75e50a45c4bf5832342ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38cd68373c562abdb22bc9fb7366c26d2b4fb37466406eb9ad64c264603a15e575b0979635f3784024477607112b5d207a6b69124e6fbca0b58b893ef5dced5353c06b19565bc70ce3725b1d7753dd516ae06ac26e6d9703d3562bad535b4e36fd87553010652f9a99d50736129ddac4474484136a2250636d11b5d15ccec405;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h675a55c7a20d5eb19dd9cd3f25b823607b4f257d298b11744ca2856aff5350023d213c39bbf226e512db5ca825491eeca88a3be06afad571fb53fc75eb39757189071911f048723c1ce11560a7e278d9d18739f2271b2890d995a1684a95afbb37a366fa2c014f8c38d1e2f08d78d44bf2d154f1f2d60217df8e74162d180c16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed567cd9120a7445784b2e35014830fa70b09771c74540fb8bbac22777abcfad741f32fb2343d731e1a228e2d0f98b877ca4d39b7694b8d975a8539a7c9c2e928b714b513eb7498b2baa6314fd6b6912e90e50b64265fc8ae72ee26e57be6a434742632d54011e97b1e9334eabf9181110e8f1ceb7dea236225a647e26240c31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc264cef8774673d929917631e3a35787458e5d27276a27af18fa4ecff05c073272afe4ba11e1a7bcb22fdcf963590e65fdbe4c4b8cd15b1e2b12fbf4fafbe1166b5d1eb60f4dc459e7c20b9ae9fa2ff143ad5f060b4ed0b39c4c9d16ff384f8752d8b69b848b430a07346b41e4c45fbe56a63873cfaee0f23b17725a7955d95;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30e0d5415939f9fcf15eb99760d2ca52b2317fe68dffb47e0f9a1f179fcb4f9c6d4af5267235ada767f8be60acbcc58c6ee9a109e0ef3033d4c03dce1de1764d5eec9373822ef5e54132c0442f6b270744b7a4c52ed07cdb7d4c826213bce60057e363449fc8311c6ab8782051bf5a1f76e80d25af7e878eab0d9025a58ff7bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c4ebd5be4bb616181022577cc34bfd300e7758260bf934448b3e09aafcd10648dc8a5823df903c9c10e9b22c2d2bb1001924cd3f558af213a62f4d4f9537754cd95c7286f1c3651e4c756b07078032feff1e2721113ded801e7a0d814f7fff36161f36d362ea674e6497a14dcf7e300ad70b46f52d9abc975e9296b9a711be7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44cc1825332994fbd88fbe07885961e12ca3893dc79f5852e325c5e42796e84f3a9e642113a19d909320ad9b27d4f7c076c9e38be5378b11bf376ee60974c64f1de4d8810020426111606cb56c3180beb203a9ecf4a1dd49451c40320388f465bf1506a543fb16a05460ab3fe7b80a2f2ac7b9fdede0827092d0f348a9c5d3a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f91b8680720a71f6def6405ee2dd42f0b7080634daa6aea1f840c8676a1c05882a7e04dbb5e8038feb829718c892e7d7b485bcfdb78cc53dc40e5ef44761897a010f0e192f15d866c1c495229d3cbe809d11fccf32a95f79e9952d036a5119a723848db9285a003556c53e5d18c9ac4b1aced1cf4a0ba04a801db9febe576d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcdc8e2e7cce23fb788a5e05cfe1b898210fd37656ebaeb08b577d537855748c003739bf2c7c0e0ae3b461bcd14087045be3860e78be9ad80a4e8f12a5a0a145cd9affae639ba9c3bd5f1b21a1cd4babc275326a27aa53c80be3d0dc65df19528001a076c6f99ee2132ebc8206eb20aa21734e92cd76fb313bc85f7f9e6a732b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bb069e2166097f99958ee53572b88073b65d688b2976f5409e83037e110fd3b35841d99f3b3ed6a763e765d0c9426fc9aec6fcbc3337260c6fb7ead69cb808807ab0941b490742694896e7b863e1f8f13bb13cc76813efc1b2d6074a4d0a3c35bd56f41c96abc3fb06e5ef1b80fb0cd9537e0167278cfe16b6d54a853777879;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64e0b9fc4cefd9b9639f5269eda13023add252750a14f5dc4d00dcdaa230bd08417b6d162c3c7d304312d321a74d9e12579d7cdd4bef37850bc457b01c1aedffbd0ee1f766ad8e3ce1b331ed66fa283d116ee6369f7981f3ec15e5759fd7be018127f13b27938043a76a418a8b1972680c916e3fdbd88f0c72713907a566b327;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfa4b7dd6ee5c3d73b290621d7ad3f032cef53f5a655f73f31a036d6b19309451fb1fee927d7dcd8aa0fa7909be0242741c3f78af10ec8a36f631fd324d7a6e6d444e685eb43fafa5479f7162fb27fbc6d9d078220c64c6a90c469d630fe2c9c45cd3c034cf42dd98e569cf09ebcbee3a962941637ef1c3499f302c7dcef692e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b09afe0bf0430b7a1b0142a120d4f37b9b20ba4db948d27bba4573f5cbfbab6ed02d3ffc3fa56534fad4182f8bbf6fbf834c40b5b8870d46b888cbcccee857e64f01a95585c5b05370159abeea0f4c87a28e3a7b812dd9567b31bca4f8c438e9f14cd94a34a0c0e74b68a49a0a4f40855569d96ae9ab0819d9d9717540dde33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36b93f86adb2466b0c079ab614d030fca210ce33547dc4ed5ef29590c8d6c8ccb862cf3277e4ac13de9be0f2b7f42b20ba766855703e7e2e5368d17c36b8cd53ae1322ee81642d2fe45f5656c81b728228b0e472607c24fde55baf8de28c4cc5ac2949d19652b0aa03ffd55f9b8d319578d90cd52cd5c70353663694b6b8917d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ee03b62740f4ef6f2292532cc440c4bbd1d8522fccb52b70ddf8ced8385f4ab9aa1f01951e3aa893a6366e72bdebba3d38259b6526da0d0a7756e8ae6a22ddbccbb426e782db09424c3a703ad9e16f2210f9b8f8d15813664dffa38ced96fbfe0c9b1443e003abd92f7e8822effd7501ed1291fb486620b616d34ed8f412f0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f2a0e66c3b2d9a2802d71e9fc7f5d038f58ac3cb32ac3b155729491b5d6ed460b5db15aa5aa4cc9dad70e4299b317bebafdbf30d15511d9be0caa738680e117d29dc5040274ad69b751ab7d5b3601ce9b285a0660c9f0756a6c83145d3bbe744bf39035419661539990ec366145366baf5c26581f7c5857d0b0455aaf1bc149;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8916ce547d751165d1fcc87bb52b83d129a111b4d38d986613e0bccbb6701e6a17414b8b21cdfa723ed6c91ab121d1b188ca4670ff1dc10cb8d13aef9a1f82ed7dbf62d8b812701007fba4c876cef9b8035fe17a55a21ee3290de947621bdc482d3ac11d5bae9437ccc9cb47e9731357e95c762c80051c3eafb79851d4533f4f;
        #1
        $finish();
    end
endmodule
