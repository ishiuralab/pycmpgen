module testbench();
    reg [16:0] src0;
    reg [16:0] src1;
    reg [16:0] src2;
    reg [16:0] src3;
    reg [16:0] src4;
    reg [16:0] src5;
    reg [16:0] src6;
    reg [16:0] src7;
    reg [16:0] src8;
    reg [16:0] src9;
    reg [16:0] src10;
    reg [16:0] src11;
    reg [16:0] src12;
    reg [16:0] src13;
    reg [16:0] src14;
    reg [16:0] src15;
    reg [16:0] src16;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h79f5507607e7f00a0fadf461a05466fcf3f27912864c2601d5466fb69d1b6cb9051077ac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h933570349ce1c9cceb15344b74db5fadc3504556a722efb4162396660c893f268eb9dd19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d36a6b1c619f5dcc45d97954ad83b38a42e6781a301a725adb26ae26135083e7b1c12ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1af60a0fcfd817ebddac7767402a52ae6602e7ee0ad9f6bab7a99e97f6ff7fdbcbdcc90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d0261bc592784d7b0c589baff6ee3eb8d72cd3df54642ecb7728e35dbef50ec631cc8e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b4307d092323df4b028b5c90cddeb9d8654015c27e20bbfc2d109ab640181751f4364e30;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb78e3565b8cf390cee16cb340c8021ae4bef9fdd8e0c5252dfe80233fd3c919363a22a39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c765cec91875cb8a1941ce66b8469851542803bd6690cd09412162011afb001711661657;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b9bd07447a23e2ca9ab9c8a4ae0acda1b777c15e0a90856e5468ace427379314b2fe6926;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f07916e4664133c5f7f0a9ff6703f6c4baf30662981630b081c9bfecb9772f59be86bd04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e07e3770c915c35cd5290705e0dead13bb0f82a6fec9ee8198146d700e8f3b5e1322e12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1541ec77760ae249aa0d05f1c9f7a9ed87cae321a9079a544a729a4a53c9eaddddb680b53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h495d43b58fce923a670055cf7c65df06d8ea53bc6581c6944359c1a4a1214bab16b82b37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b12fad36103a69a2d2be37c9f5232714a35e2af2536da02af9c750fa1c3a00cb6b38901;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14010857fe6c9090d4aed17eaab0e74d927cd07e7de1f2677b162b37eb2566b0bc7d4e691;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a90994fb954e39f1118fc432184f565884753af1b7d74d4a0bd1c9d89357e15e323ac0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4dbc69059fd36e955d859b4eab72e0bd96d3eadcbd3f7550784c322ce98cbb9bf143e4d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h618577bd0a231ca831de925bb62192d4d1bc1ef5166c6e32489ba19442b629293d6576e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1440f29a72871f4ad9b4c7d95b01ad3029f0b5ebfa1f800641a4da9c0e803fa11f65dd3b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd46914344986cbc03c91ef4b5d93593be15503b89d090bdc97f76d130f613e2de1e3d20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbd7654c9625777cc027cc5fe58faf6eca68ff5255abb99aac71ca5362f80b96fffa0f22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a534d1de52745bc001e96a0e8f075bbd0072474218d1a86433608f02153af2f42a430df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha4eaed0f49e73996345c71f716bfbf5c38ec6b8c417fbf6b6007bf9e443537191d3b78de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfdfd99cc162e3a51f48529ccdf2d9f0590561ec9880955d5c430106ae22017adf3e90744;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h845239c9d6cb92bccc1f6e507261277817f3fd9fc1f983a4a6b5eb485677b04c1c798cca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60ed6c2c2fc07cd5ca744315fa961fab450cf2ba697bd746b864a6d004a64d635a8fabf5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187877b7646b6445ec2abea7a590a19dd6f173ea503888ab7178d0d99cf6f9a49a2b13dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e63915ec5e8dd69c33bb2ab27ae7b6a797e8da0350250695639133db89214055f8d1d09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5994f46fcb4282d0d07728d335857d02cfac96b2b48ae97ee3684911dd6e3b6a2257132b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121f0676781d67093718f2aa44c584e8c99a99290ebd046604133d4c8dc241cf86b4043ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h55754a20eaf2dc7c16ad699c460cc0f48a305ce82b0f81ac0c02e525fdb3f6ee6830b7f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6faef7c907fab75d0f4aad2ac514f93355e21e4ab49b72b4f3a64d482b0692363c19974;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6de1b26c1c6f01343d474eb226fab4c50c07f302b85ab1157c4f317c07904c9d0ad72f72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h27196345127a8c8ebe610f31d81098bd13e9db2dfa1f29b79cc0184988107d6f7ada57ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ed40e0158b7ec60e050bb7530f2f6a2246c689c5468dc394fbbe2b55f6a00c564b388a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b1d60e94e85e0965816078c54ed8d4349547881406748bf8c05d8f74151f9938a72bc9d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f0a373581f2a9ac97a5bd623db600266ddca30d1dbd9a9bd3ce5dbea07ff9207ef1f4bf1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175d4dfa7dde67cae81e4bf10f0a6d0c26241b3fbdf4bd9400f2a32017fb02a077f29e2b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2c53b646bb3a6f3fc6057274bcc92423b8654df704be30b5b21a78563080138c3d0ff9b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e817cf1035184c0436df90a52de0feac65a30cb3a6792530b5ed45ddc5729621f90c29f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h53cf3c746cff957cd7d90fe8807b48c4ac61b1f4b44c33bd9932790bfbfd931407cc0e67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e40ec1c36d8b4484289c1e6cd2d2b601a8d0425f1cdcc794ada74ac623c7edc08b8fb59a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcea8f3841cd1a6ca1daa8fdbe88d138fd63925bb014d2db4356c20ff8ceb0016a36d9d78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e98818a8506805fcb584db965f631250418f634eec97710bf3e52307f7fedd3d4089c9cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194b8ddf141228412e1a3879172b39186357258103b04f236524d4805c6f3ad2ec9610b5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37e4b9d6ad73d3faaaa0bf4abd72cd993818139e25b649376fc80cff3389af8b6e6480e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18989db9725243c9fe4aa597ca869024bca4a4df2822cf4e787358d464ffcccd802b3eba4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5501b353ac0f19a86013665154ccdc71afbf0ae44fa9e9adb8d7e110f64c954ecf95ffca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d0dd26a359a251e144ab3d9eb94f197a7007930cf977b0b60b5f69c21e0542758db9ede;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8330428e55f3d6a538eebd4083635e44c7c7e0d3b9cb9de868ee856dab82b37db245ea16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164a4e3976c9c80e32eb133ad57610a3d6c2356c3f2a37c6cadc137cc5f67b09cf9d6cbdf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he94706dbe3366b056f41b83c72b32778494bdfb5cb5deb422881b4c4ccc488f62f7a2bc6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba4dffd293afb4f80b135c4781794041a05eb81f0e97407a431c11bfcc0512418ac8ba9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d828b65084a47e673cd825f154a3ac5f09b6d1861874f99c8a694563ad69624966ce2645;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2957f605df4f3a4d2daf5b7609dfd6aa9185fc3a5a53f5a0e2ac5517fa5f38019acff09e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h834b4170a897848154935a051dd46eac42ee34ca106ba6ce8a38f49b5bf4a5815d1fc274;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f026fac2546e5d9f9ef83c2a4e60d6ca5ea6d935b0538c3fabf4517ccb8415703bdb159b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e13e105e4da65260da0c5dc48ffb77db3b36bf9de0952e364b7323c2d91c2ca2fdac79e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c5eaf284052585e0c900f7f6dbee473ef9b0f05198a06aecece512000e6b4e9a405f1e9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1047760653a54c2b21d61b21cc8f332d1330acb79fc17e55fa569cd8a5e2c524899a6fbae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2dee911280897a2eeef4ca2427bace8fc4c0a425b81fbb189744d329f48e51911096dc5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17baa5d0bd87d5c0c6b7766a695fc088c1375b7a1a21ad73655f83e35f51fd59eb16759f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h857537eaac8e8c4ba033c703994be6c610484afc39bec7410d6139938e5d8ac1832f6f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf98704cea86fabc875a10c4031425003a90dfeb594577c24e73c7f2f95ee1932c9d36d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1780ac30f7f33254d748b2819fcedba88f72816407b488711b988fabbcb53a8fadd8cf5c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3df34dfd9300aac545a655228c9373988da188cfbed760d98b5331ed4cfe8f39fa887802;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h270c70307fa2aee294069a2d25c64447206c03ddf8a2b663961ff7e43f0993d7f4459499;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105b76bc265ae4244b9a65bc3894bd9b6fb6a3b685d50fab08a861f0df00d89d64f7e1ffa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cdfacd031c5678f8e5cbab8b7e1ed83b9ba66cdaf48e88117da77a1e248f4d9a0cf8e1e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h673d8eacae7cc95fe2ce5f395e88884d480e34c8a1a64e708ee611d4e02c4e4bf1b79a19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h393b9372484dc9b9c14dfa48457bb934dc55d33ff210edca75956d46af61fd529f65fdac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf8e94c266d3458d29670fc09f853d60a2e463ac4275a79fba7f5840c4e6f6f317e181250;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4f2d5591194839070c44939760234dd70e4922bd292029fabbe95b7885acb5c1678f185;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7fb1a2eaba7842429d2ef842204ebd1e4c0a46e140ee702837eaaf875fb157050977ee64;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48e4c13ace475a60c3aef651af9460501c94dbb53b3ded58d29695dcb46679dc2c8ef95e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17ae24a340811e2d6a35c3692b4f26335a70698dba47f6fc18fd1c5a6509a74bed82eb4a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e334660c1513d598a34ac1215ca3401d89f0b45d6a175028e8acf64fa0826ce2b7e21361;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158211fa23dc939186d0da339ab1ef9afbac99267546fed6f72d3e69d2e4afe243c954ec9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187f56eaf0059ada550f2c8083bd8e1b2038cc5e7bfd5098ac44bba20ee375e4f0c4a349c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1688a5585d33966f5c415d7a97d628c0f5c58b56c8346d6e57509ea1f566962f98801d386;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8ab972d1739e8d2fd1ac8fb78ce6d1388da0f53b9ce99b67ffe41f2368351e7e6ee55d8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e46c76782a304d69e61c5f5ee7a8967139e31bff6b1b300e736d00032babb978dfa15cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2afa83baeeb839787103980f21cfd62b80be9dd108e6527526365e7e690168904468f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4675fbce24edee746feda32a093277634cb4b2ba89af635f9b109861268ba244623e323;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9833e76cc8b8b6c753489a0fca9af764b0532d3f46b6ab4ebc8e02ee9de55b70ded84b1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he86ff124bcbde23afd16875c8a4897487a1b7f460c11a9b1a94a5eaa64a661f9f6875f9d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5d75ee929e1c0fe35ea771be0b811efe8c78df5666267ffa43244329fcd19b340521fec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af16323568508a11c334228fecbf15182af47ee979374914d4e8e1980a70caa3d87199dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d19808ad4551cc895ad5108d302751bfd54026659fc618bfb9df0284b9e8b89a420353d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97040aa3b979b26c649809a0559d4dc7715e25fd9ccba9d9b56387359868d9ffef88ed8f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1180798f23d6d12dfb2c468e37d0186a35ed440e43bf8420bbca719274d43a8a8b1d11d83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hded72d81a02b694f7f662326714d2e948485dd8d634720c097c6334945921a800fbcc241;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h936815e6508d104d095421f50b43ed04a3ed1687219159a7af7d4341e9bc1c068ed1c54f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1efe9849e9a52912a6455b1b1461c7725acdf42ba418ce1a482055af7b993f37c581af369;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hefc931e2be5ff05e9eede443a451742e0d0e78dce50440778e1f4ad5938ab5cbeb1a1550;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5c12b7f5a17f5085e384f88a0893df81a6aefaab94ec8879fccb10537ed057c9cf6e987;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f81b54d9b343853e23734006636d4d27dd663abb3c2e55fc866e2115680b0c7ac83b6dcc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13dbfc5670e54c3196493ddb225c07389a8be7feb86c45a02f489f3decfab1c40ddca9d0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f185d735b18e9974b0cb774ce454d949dae0f6b64f5f7790415701101aa82f1ec9f588e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff13d9198fa22e44fb3c4c79612008f7534e2ed758a7e00944af333f4e1e4fa8d5dece5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa5ae58e73c78e8933b4c564bc895344aea21930fe43951abecd2928364c3d78cb5e5484;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fa42c4959c6e16a02b76790459a8a21b6bbee689a0b1e2e1947f863c93507779d4a6731;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1096c3d47567af9efe655fdddfe19719d25c6afc0c1e0d1946c1d5d134778927797ef2a39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47bb15fa201e37a36442b25f0ddd1f1c92d72fca522033fd26918f79dcd1a8b912a20fe1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae0b4972e6415f2e78fb4558be1e13cc1a2129ee23be39c60f9cf5e3b1eff5a72f535b7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1159a1aba7ac9d9927921bad8c71a5e7025ae1555a41277168a3385b2abceed95cbb84a8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h890c0d5048fe66995e1609449672121f52ca857ee12afe1e68b80dce4fafc2bbc6027764;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5d0664ce818ef641fb36386bc721107f640dcdf8eef8a108187ef2586d75f70306ca56c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fd199e5d0d9b5f2fd3c39142ce52df6f45d901e82747635590ee4907fe052acc3e687a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2868d6062b6ec9c9c134bed51282ead442233112a9af9e9bc90760f89662e9cbdb83ba3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h459216a7dab6ef8800f00a5834807d8f70dbbdac1e45a572eec8a1c41c045cb0aabdec73;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7238267a455902a4df157aa3e38eb6a26a534d76a2e9b79bc21a56b1997b963f797f8c2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48f2bbe30a622540aeadaa0a0a6ee28a81ff70aea49a69b0bdbad3147ba31d259ad189ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h173f947deb61572f072bc6aec4bc35b988a29f38b60a748aba7b0b949fe9787d4d9692a36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e82f5a49a539c9799075461654b659ff209d4ccce0df4e9efdd9a5d395e31617f2863cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee9c7b91b651ea28c03840fdc0169c8608bbee70bd533dfbe45c23ae007dc851f0a18a3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb87aea562ce7fe72ca4339c3f9c103ea6b8a08b86091ff2acb9e40053bf7efc90733aeda;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187394ff468c1a555e8d4d3c059ec34f38c59ea2ca0d71c1ae3b355c8a75d9dfce22271da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7632737da843360bfe5fec2237794ea5d5295aadb741871621310b55b9c68c72fa91c940;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ccc0a621ee7b6c825858da57e0428deae19d579b9214814d821992d1befd0ef27a4227c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98a63aed9a7bfc78a2a7dfb4dbf279fad7b159dbfc6eac43efd6a65cdcb826c06b2f0eda;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h186914cf34125c615b991a73a0a0877d1eb75532ee727cc66ca1c49b0979fe6d254aa11ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he09e27f0f499e5de08c0ac7108850f6c71fc327013b244c63da0b8cd1a45584ea80fc7f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121b112c8576cb0f94ce49458052696021fccb69a6ab2679adf5a76f22117897fd5854be3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51d2f71e922aaa04694a5b1ee4c61e10a01587f38199912a6f81d0b9295f0a6870e49604;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192ac046b9b7750b21acbe2a570af1393547cfb8b409e07e0f10c03ad47025f593cc9ad1b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a6dbf0a06910f110cecc5b4b6fd3cdc1d80b726700e65aca012daf224ae5aec0f343dda;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h253ee0839c5fe62414c7032f26648568c76d1c0fcac0cec7750e667acf2f14e579998592;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha8b19e170650914bddd405d3a064aa5823e494cb1f0d025119e35f5be8714369341741;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50d6464a7130e490d77d61812ace1cabed0d33412abeff1c52df07e9f04d130791b57f94;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe4387c4d7e4d28aa601d4cb5be29d116382f0b720f4f02cdf09a9d2895683cefaa212d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1952d236e4235c0f151bfa9b7c16d230465f4e94e0d9d794d9e754666e7f036a0bb16f77a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1cb215c7141602e52ec424bd2e8cb31e09aaad97858cebfef223280765dd263d8f20983;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140fb70f71cf64adaa0ded4e7e329ec3d60c1071b05cca86f24afcc4f7fac1a7f2daceb74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11718235c2b3afbed9a8bf8490867951c2ed032cf708e473315dc7ce27cac3f9fb1b7c9fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1255b12e6b0195927f4764710838d993ec8ba360b575299bd733def7a2a294836f6ec15c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d21faf214be403d580438562b6df29d36980270150d33a1ce493ba54beac1a449d7e974;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6ad4fc961cbd034903446ade91f4f42f59a59c04276cb1158df40f561d4b80e3b9e2d6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1721192f3b4189edd916e4141154ab94f0f071a4b9fd36fae072c8146afb6e06acd7130b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec8e08d49bac2507c154c5ce588ffa68f515b6a8be09faefc5df8888ddd955984160523d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h163ab682a461ae9ffecabd476fc24c598a831451d61edadced6051b03e634c21ad3988df3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f79387e50aa575d30b9d68670b3caf565447c300533a09f6d08d874840b1d0b048bd5fba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c61bb2390ea9538536dc610e212d37e86c3b13669fccb6896cf62ca7bc702451ca0d80d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153e6cc24a73bebe9a3a83c15401d93ad2542a300758b14d930d213b3525ce97a71a4a3dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181c5d5a29b7663c05ae29bef59b9c962b1eb9238b3687432969de34c6f3dcbfe7b94eca4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha88bd9cab0b5a81b52d7be87f99ad720aa192d8dd4b65f505d018ea36534f0358679be63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1928f5211feba7470c939cfeb63a6d1d26859439218f00cc93559ab2cd3315be5e980bbf4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d194583cfacd4f1049fe9452f75f447b22a47993c5795c094b82f5df81b56203b538cebd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3c4787fd87083b0fdc4f15c263fb072d1a88e4ecf69cfa90108af2da0b91c606007eaf2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15dd151163efda313733dcfb9e2192a7b55d8ccd3ef74427cdbe82e2ec403f3b8c00205d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62cceb08440eae312d8eb854aea17167fec1e4b8478f33bb337e52ebe1fd01b942650740;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb176d6f213ae2367d4fe5904dffa53d0e48d903422a60918b5dd75565202289144c11a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d9d527e08fe1100bad6f21cbac37f28343104a118f8dc6f3c933d711248e1ab05cda7a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb1e5dd26bc8f17f150f3435fb291632c174b8197b397e6feea25b3a082fb4e49939c8a74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4d1446aa0af12b44a21ea499a920185296b04089784dc0550c3ed6cd12282094057cf31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c6d0d855f436ba3235636c0e31cdf864b2bed78a82a2c26c2841ff645e46c50cbcf9435;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37d0380ee7b8f49f331ad8c4f9180fd2bf825aa8b91127ce8ca12f53de26bfe0e6f483bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98a5d4e8a79ffb075f77fa0224905e64d67028457242752cfe0ae2a9f052a97f4e9712eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1225b978a07cfb02eb2f4f33ed68e99dffdfa684c9cee090c7563ade87a3735134757b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h816c8ed93bfdbf28d42145784752e0342427e1309a6012255b2b19e59c14e74a5d13bb50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0399c65ac8f9fc04b4370ad923ca28db9dd7bacfb5e47a49308125b7ebe0f342d950cf9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1255414ae2a9f5fd996ad48a11b4d2176611932cf16059687c01397ed5a7b361d53a7573f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f3434b1cf9ec4f9f9219814d62a6f46611320b6e434e73b2d549385489e2825b43523be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab12b75f859c65454284e5ea0b9c61c608779e876796676eb2bdb5aef8852e428232f360;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h387951a5e5af15fc74f44a0d1be1268a7bfcf47c70230780389fc7c932ac205b62a3b21e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c00cb9476ddf90eca47d9850106174aa833957af966d20e72f41d0eca253d3ca88b01d09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he636111234732cc187a4390b1900c38b34fba3ea6effd7967c1e614330ada89c5b59eea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11670d112bca76b3379489ea55ce6bd3db3e5099d74e1de9dd26f9c8ca74c34e57dc8dc46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he937ba07fe574ec033fef0dca5d3237f0893af6c6dbe5f10130f007d45b217f605913005;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5033aa905decfca2c5916e3768447ccf5b088b17e8b227e6ed9a73b6eea586ae2a6f8714;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h78140a58a779d893c8c02be9429baf57ffba68928e89955003eb4a6049aabd4a961651db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8debd4b8b6e5c3fe06fb1177e1b405ab7cffb228a5ae954c3154454e2442ec7d6dbdc4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d87cd1593c288394cceac85afac427f715d2e5cfdcc723c5c4f6af0dba490500814d03a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cc35a9de0c60e58e331796c78694ae9204eba5ce126de650168d16950cf2340ac31efe0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164469ee433d820b94bdc74789b381d30ae6884c0dea633649fc5adbaecf0e75961e6cd6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1d8c3bbc778edb84e3e363720b755090563b90306bb37b0847527802d75e911e7648c18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d9d3af53b1fea565cf7cdb685ea36df4d4016eb0a8539f5d663e0d12a321b2c209b1d54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h99d73bdcd2c6839842e00b3110d518c80ae5a9fcd22b27ff37b27080df90871f4acda288;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4274126060b3095221f44d2280684a5a07b7dc0dfa35f5c6ae496365082125004868f4e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dbe5e7b01e7a36ac90257ea45176f98ffd51cb08ee523bd6512aa946d33f62af5a33a24c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h927e812cef25e99e21cfaba02f931b92d8e330322f3027749937ac4fb6a82054cf5d1d83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49061875e74d01166f0adc8aea334d332471fcd9cda5e335239f2ce27a86a8f0a2b0be1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f9d1f187c89fbae290ebde577d13f130cb279b7f68835c1b7e1c1f2248f58610cfc9e32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc019b0ba0e4965ef6c0fde8179d0e6f848a31f63b99c44e689f609e6b8c7c61969376ac6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2fcc034d02e9804881079bae00fa8e2258547fb103da3f77c0925716881f952f7ef76f1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14fbce516e641bc6ffbc2dbc57a98c95e1ec8b128890a345b1196299b1a006270be5004f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b31bd47b03857a8fb9f2b5a5067ef9228f3532ce1aefdfce171e04211f5025621b58df3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109819b8aa54a7e17aee5ff3c7463caba2d4d0b492b72319f54f928e5bfbbe55fbb8b42a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115534f9b0b3dddaa97ce05f678979323ceb74b972c8755a9d7ab9b05c3429e34893fb071;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a0dc07ee1f7a3e5bf2f74518aa1c51510ceeba3d118120f23c38c6b3dffd1590a412e76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d4b4a1e8513b4c82e8abad3047a1ed97acec857d37d3f7307a819ed17ca806b93575045;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8b182278570493bc9ff7bbde1ef30a8b6bccd6cda8e8efb11d6a2ab63b1990a999509b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hac2c08b82adcd1e3749230304d7af59c5076930b1f26b2a9623cc864d53f2de6efddf904;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bffc012b8586cc60b76b23dd941c8a38573e105cb2ee7263f2529a726c48f441a3c3244d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134d283431c1ac010ee20e35c0f917bc3de8bca963a6149a0169e07fe75af7bdf700a2b21;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hecdddb59c7d2b5e05d9fa3ac97982eeed303177554a6d1891ed0c4224acff5c58e0ac914;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha4ec5ee0f69c73c329a028f12d4c473e388ea5eac0d133f824e1bb8416ce364e6408e107;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2f6efece4d2b3437375bc75eefe083932a45638d636076fbbc0d9c3211c0660792705598;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9abc8197bb5647d26551029e1086ae0a5f07a8a5cdc8f2c459d2af4c86b527ec0ddbc530;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6253ed554d632f2747ec95acf42d3b54f437dc032526b0cd23512c1c29793cffc7a44c3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf6b6182ad959f281c8904e076c55cd4b5d6780885942c9fc0b4e73bb986c9dca4747e69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91fe3890220442bfbae01c849abc9d3c2c1fbd97a655c9489675129ef64a8c29bb36e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f998794c1931e264efdc6992b7c86ecf29c167c8574e17534d353d921465aee1a47f138;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfdb3ab53fa3007837f775012d35dee254c2a233d501c34dae88b5f8fed25183c2c7cc8b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b4359995a9f393f3605136250ab88c84f354dbd301d00290ac143cfe9069f57d800fe38;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hccde43d2c0338368fdaed6e3d74963102ba0bf8ffde8cc12e5cc341be30ad11a01449fbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1433c47e58500005a2d6482066d7edfd3adb6e406f2d893de14f68aca06b790f62deee9da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23eda48888676706aebdc4b2d23cb318468eb580939f7b68d2e0856552e8eb1d5a1a78af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42e283704aad17cdafb22251b4f5c3fdd77a9d819047bfc5146320c21d9320883727db58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51e802a7cb515c215bada593bdc96c2f304353516819b89bf4105ae55de65de9b287c37c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fb98414caf5a2376184b9a21988e3bfac00770280fa689c453d6c0ead97da9daa0ec5f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13660a4d5a2864771d3a410823e7dceacf93eed69d8829ffb73c12fc2436b64ee59a0de7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa6f41c0f39cadf542712c5e7d8d4cd6c6c482eaf197084e1fd6c918231d69c440ee1034;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5324496ef0a74250a15c3a8f9296d907902f6d777ee9a8ead524d987515996fad40540a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11493112d628ed1156f9e7573625f55f3b80fa8919815baa8605ec01eeeb4c8511f3aa4c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a670daa7b5e56150d05c03eb34db5022d03d97ce693dad03629bf371beb0196e951197e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdfabfeb31afa3998472b7cba095f694c1c960f7af9dc136094e1eda23d1d1c4c2f332fa2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eefa147ba7980dc6bf624543103305da671681f0da544080643b4ed9c58e5ba42d60bc1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b9368fc938fc3264e83012ef41bb6a87d1f6c6a2b96b394df7c321aaa6a51afc9d22f4a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha18a9f27ab299cfa5945ee1f3bb999ef60157db492e2972c71544e4774fe0a14661781a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154d167b64534bfdb19dbaa451e80530610d681bc327ec569d102366302c58562ef2b78a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f4e23d5be347e0efb23013e0b5509d7c8a540dacbb2435b9fa4ce6b8054175d2020b8c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9e28461cb4f0ee22580c9be4a6cd77910d81e08cb7c15bf650ee06e5a88ec0f5f3a2cac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc578e8f5853d2ada4f80ba9de1b000b2807e13bffa266b756005679857a2045bfa35fe0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16121144968704cfa7050250b1f7df3f61e97548fcfc54bb1be65d3dce7fbdcf4a7a77e0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12187a607d62911ce95d20c629d8e5908c2a699be78b09326b97354d2ba7062d71fb5cedb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a5ee60e0d975aa245e17786646ae57330ec15a5a5752973eb3a2e4553a9f65a5212c203;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66ad1f718003a10d147b230fe6b61a52e494e3b8c72255a70e3cb95e0bdd461e46847b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3bcb67a346105507249a324e818ad579dfd9c6519099acde11076eeae4bdf4ba1d48f7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb361e7f2c03b4807fca689695d2a852fc0ceb032d3e36019dc55ab7a2eaefaa039844855;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156e2f09bb041c24c7a92cf4fce812a57c4112f139cb50136bd693db95a466d0f9d2f394b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3fb375869542c70a6350cccaf258ff6725c380cbdcb66e12d5d168df4ee9d25509338d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h120bca8d77c3a78a583592f3c42c62db60ba7ac38ac041b33bca8f27f619454c918fafc0b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbb8bc07e31f1aa4e8eab618235747812f3d231426dccfe7330d21607d833d318796bc8b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e11c5f1e9c1c81918e91f0ab5123865cf2ac3a39af8959bf05607cd9abedd860c91498d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1acdfd5b9941d05f173205f6c4bedc452254bf451aba720b82c2e9c9e82052a931592556;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e5fff3919727dc7667355b6cc85d588d691d48a9fac83a92c1b15f2fdd92bce31a7c45b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1530b9930faa0b0bc40379c044a4948f9dc386e5a77ac6dcfd0fc1a39335f27dff63e40e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6f5cabd6da4f2c5832f66f135565327a24e16c8c3ce9011688cd8cc8a33fa8330c5c4b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc4018337514e8c01fd8bbb9b7b271d87b3aefd08a09516c60d4b15b960845208dc4d0044;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd675addfd5cec5efd6c1dd511bc36ae66b96f8c126765b3b68e97b8a78bd035075dc8fd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c88e8bf8c8f3d1b1292e2a4867f9916d1fcfa9ce6b3037d642a2decf96e1400e1c939d2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c43dfbb4fd31e8242b73df13292c4642a9c759a74f0b9499f97b89bd0fced10afa3870e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1414d0fe09f8f4027496e3cce6927a2cdb4b02f6705cc98ee077cd30e07e951f2033c9fa2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed4e15786dc34643e820f4f541c366a70a308b8b8a559334dcfefb7002e21ea071a8a762;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a0969684443a13d2dc5d40d8a1aad33bcfd7247888728adf37ff5e616197d9186b4512;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c8b950e00ceaa9711904c26bd57dd9da190996ad485122691c1b07f38f4ee36689758cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfadff85ced7db8601c3ded376a72813a367569299e4380b3f53869844f69827612cdf447;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had9a5ca1039574cf9da3389bfd375090d0c4d245023cb79e0b9b4eaa07bd6476aa47e83d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h126c183ba088044d48efb0b98202abf1c38cd871dc52f27f1820847c679dbc4a6f67162da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12309a8757bb5215cbe76026f71ed9078dd73592deb5f6e19f2eaba475f9e6c025eb337c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf292dc642afb81269c66d9f80209b7854a50a1b12b3267075ecb93b31c8a09b848a5f263;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e906a3338eb486758934c85c485d54edb5532cc6fa15de5325bcb9f784872526134739d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h56d3b1420adab06db227136bcac806b24b5128ab9602194ecdee101c1fc10663f7cb329d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8166c6c0a536b2c90662917a3e06ace4744cb61a9c9ac407a06484f2d04eb39eb14d283;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b00eba0d36cb8bac782d964d3711e9917c55512611e2c05aa838075bc2a612179c71141b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a50548aa8d104b23d93db1ee2b5f40a61fc04fc93aa38d2c0c28ea17311bb02ca04b61d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86371c5ae318e87322134aa2e4da831e5ba4cb9d9e5b2d082cfd9e4870af7e670f661d52;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbd09e8e7d0349a136e7e93545f6d710be8403889da43c04bcd4452317dcd2b8510ca744;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c8206d8627fda03d13ef7111c409b3a397e94e228ee9e405a1ac49bd80cd86c7f8c659a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a96a520375bf13605b75cbdf1f3c70d61294cac6122e39d74ae266c820ec9412ccd8235;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc68fd340a9c4ef0eb313958384f2a47003c4af0536aa2a4cf69ae0a971ca35378830c39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heed65da81b2e4df31083ac30b23bee7e1a80d1ba8c327cd6d7f73aff1c17fb3fb94e1d95;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12be7424fef69dab72e21f4edffc797472db8e0f2bca8bf3a6f103e8ad1268b5dcaf70d62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h790d82c89b3d9b1ff48dabbeab556a489202f38530b4d8560c9e2c7297d21602acca3326;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h96db34b1a01fe5a4fbeb65d397d1264eb0a78817d839173769cf51e8aa9128ac9afa74f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d7c403dacbec01677161419dce5c6d0e1252dcf2c69f642a6b217a0d6881558cc33eaf8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f5d13ca101f7b8049ee30b7da7fe970fbd2308cbfbda800a82d86678d72f6229214c8a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c61d9342e1a909f630df886cca7c2e11e4c8bb8aacbb96b55cbe7b2f83aae2cea4d1e19b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1237dd6706ed3ef4244ded2c362d5731a02f4707db982863b0b0328b076b21dbc39246118;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1acd0363223ab4ef014c40894bb399801bbefcca7dffc9c83ac0d7e68ede5b04a6851067e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc61710c42e6a2e33e84ee84bdded2f6005782af2d84ae468474c0907f28cdd72d69c2948;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h106bd95e2df167be2c1dd8e846f6accbb1455b8f98b20214eb2f6c4ad1b13110a1e8d9de7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h79ac10da76138c0103700de2e67d8dc638579d6391e1e44a4a7e5fb1fdc386d5ba34c9b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd690290e60473e163e34411b8b835e7361179a4791b162b2c19658f378be4be96592d028;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd6948d4be94a2e637918dbca12a012724ad615afa2b42b03b998f023cd3d76a2dab1696;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17bacd5362a8682147989a5bed1731c9b8c09d263baf28593a8c5947dd7eba15635a9094f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138b6ea16f5ea244e93657a0ce3ec6cf4a927bde18c7951e6e0e2d413a8bc971695a8c825;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcca76b9fbac6f2107dcdaa43eec95a1cbc61d2c755c02f5427e5dd61e8b685de40cd5c0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h687824ef613e4cacf78fcdbf21ce7bd6b9e3effa6f88bee8c0a10e90c8245e8e38899be0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e154e8f7e6afdec227a578b77e7bc02b2e70720cb45e65545680bb2227d88ada9b00cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd3b1c54071718ac2004d6dacf73aaaa423f4c6815bb1481f58d366cb0e536417ebf733ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dcdc406161c637805226008bd1b2f2cf2fc716d6fab2fcbab7112244eb0165e315d0be3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce6b6a1f7aed60631e6ab3383751feae1a8c52719c6c2d4cd6ef97164ee8b919568987b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9fda141682efe016c40a30df980977a55ced652b2c9e89bafb554c2c332a8b37950d4299;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf1ed0ee6f110101566d611be5fe5c4fd22f94285e15ac62a06bae20b22da143a95b03068;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16fb446b0f842d6cbd400c37cba0c145524eeebb239d1acf86b47a93e5ce9f4f043a3d9a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1365dd50a44d0c804a7aaef0257aa226f7adf74f46c8cdbf7630b3f7c32a62bea09dd748a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107a80862a3fa538e38ea0805f1ba63e6f090b68a78c6b7fb2e742126b8f337682f39ad12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d64c0f93a174cbe27ca8af52a047b8ed81b4830b1e5616f54b4a0a43e7aa1244a602a6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca75b8e8cecb3b8ddfc5e098bc4d216982b16e28c8e72f6f2f8cdec0cf3cde87a823ff59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dbd14e9b805b0c28f6a4a4f13eee1c53271384bdaf0587b70f326b8210e77ebbbdc2f366;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5edc8a028ae9f7d1f303f86c38d52db0d82f28f2f52eca1d0b87af2ab3847155f001198;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15971359890eabd795d35d8f5e083b07a528d3c7ad12127d9002d6e40d5d7414c0ca276d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2657624f551df8bcd1528488379ec90cba72148003d7b17fd6e9451ba05a470b282d4c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2839929faf8b422c81f1b9061386938c6a2b08bdb9ca8953af1366cc17f8888ef722e3d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ec878a662fa22522bfeacde6301a78547882c35b97e589cbd6d8f0d99c768639a34528e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1108d325bdc0afe7566568ec5c2f3bdf45d3cc4421e1a3d0342aa52a7ed4ad86f43ba1336;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfdc274ae9840068f11be71f52e7e9a77f2749eeadcded859f93837a53bf00203576afaa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4c64b8761709a0a002e985523247973cfbbd07c264acbb627d962245b174ab021c44ad8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he5e1aaf586943764fcc3bfed370518e9bdd9fd731bced3d1b84a4ff2d5db5d189c83ff2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae49c48d1251fc115809b2f214d5e3499e8e8daf415d24d3dd4dc013e7aeefd0857df857;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h689e02aaaf07080fc51a6c8cac0a38f5b029b50c914d89352d3f228c24cec055b789f72f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f25927b97120bd01dd530be3a7360124ef7311f5e7f9576e09359c6eee3d3bbeaf864dbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107e126178bfec6c9af62a23e7d07db258d42c8b10c759ab64e52e532c86ee750cb30c85a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a748247c297ea1996a9f3fdd3b5d0ba8bb64f7f894cf82b200ad58be4b077b8ec2feab51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d11c0a14c20fc73505027bf8acc5f8b93910034e308f343586d6b635d65e9a24ac86f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h68a87d3cca2c8a4d464396b64711d5403d2fa3525d512e3c44ca86bf67751f2be8692658;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heee938c0482aa9b560fbb4d07f1d74115026d44c562eabb179a59fb1fa076bea8188a095;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he6821623410a076c7c9a89f31487ebbfc01d19f4e39eb65896cb4bef05daa920fe85d33f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9c119949e6cdbe06820cbe62dc9c240a86e59286675c3f4fe2c8f1d557bbac327ebe264;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ee59ed5bbcdd9bd0db017c613ccfcadf06e163a8604c8ca8bf90ec7763bb82f206116cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h193d00cb9e58bba60d7b473f472a8a35518ffafecf26aefdb1f3ddecac2e684674bd447de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bed4f74167cb24afa4e0d48518a177c14cc5464e1d2cb0f32b28a3aa60efa606e6b994b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e481c96734b00b0eacbc9adad9d431caa492f148a67affb8828744059e8eac8494b75e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcbce35463460f0d3c36ba30249a8e6d740feb33b90c893ef9c2043f7f128470b84edfa81;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb47580b39e6efe42ac6a1bd8e18819d35f3ce04af1ab53797c9623e5d07ad4ea42746623;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11741d540cd848702e46163df55488fb040a3ea0fc2cfbaa4326b7899347a03ff8fdef889;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca060ba28e5f5e567f25d52f67d59a76f71fc5eb87f36f21c597a72b3d2cb6b24dbee1f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12fc7e35709d9509ac0cbe2d45a94094a5e1281707fb5b7c667e81255262721abb68066a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19250cba35246dc6bf98494fcc079c60877bd2d517668b35f4c68b63f5af9ff5045d9d3c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b78ef87e932094c2dc9d57bb45252aa1e36b796a0822e564db5dc552b58d00a093ebabb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1007e21f4f5a5dae11aa4bf57121ed02a5c80e624a83dc56bafefd53726b321718c8299e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd0ecf473c853953366ef0c7a0b9a0dfde33196835a62ae4c8dc2587b857ed3a835ae905;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a44fcd1b667dfdf3ccf901cd3af2438a9024bea9740b8b2ad48f14bca50a4553bdc792f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1933784fc6dd3428cbf4988b093f8d5930835c9bd24946cf17df897f4475d9d68ae81b47f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1054f2d2163bb74626c954dc8f564748c3d26909ce090b3c86f47d8d5cbf91efc40352a20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha5870ce126c222e4e989e96749e9ed2f4bb06203419e1ddf46dd3ae4b937677b9a55b725;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b97a58fa53cfd64b9cf38a7c7db183369b95e96a4db676af7598b193d7d5a67108d12de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2eb62e419c53577df0f3d9ed614f010f61f85955245ffae6abb6dcc7ccf4bcb37e8738a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3224f8265f106415501ca252384354850d15a06223d7accacdd1420b261d0e676e444ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b501bb8c472ec91b795f46373cdbc28723785b831865357686244445ffff887d6382af5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdeaaecc19bff98def934e41cc5d18529ed8389ff617ae9d093d421c63a29ab6d88020d32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6af1a6f62eec991086f0b3069d7a617c61f65cbe2a3a1758808fdb80180df9965b373865;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab039fae4e8cb4167cfe99d5fd4426d939c455d2d54302e27c0a4c0dfdd5c5db83abb093;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5805a4056f66a7d9711a56103aa770086f6c6d32044a0f343954b098f87637a5efe4a21b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134b4a3473811b95a31cce0f847147bcd7db16e3992ce0008cc9a5b802573199c761b76e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199fc82e09746b978098ede5bdd1aebb74b48c46b9bad5d9321abeec4c9f95d4b0796147;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e414d458d58f18e1c65107451cfa7f10f806c984d6d23bb1c8e33e0562e6f3882bffa03c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdcc199b7949ec39a4a641f9b15544468d691db187c09c9bd41906ccb862b1bd091098d6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba14862b70bf8ae988e04251751531fc3716f3c7e75543c3842d917f370130d7fdeb8881;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha59db00aae91004bc8b8ea6078c3c0b7039a424e60b44f7ab4ad8d2fbfeaad7705de539c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2dbe4e9a9e587daa85a3880d9fc5dff4b247087d9cf793b9455f959f8dcb87429835f37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b813203f38e9262e2a7ecb892e19ec62545681c42dd6c01ac37c543fc1b78824bb4e544;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d940476109dd9fff4fb9338a6c94a674e4516e2dec6b11c0607ccb70305581d3db4829f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14adfd8a59ebb67eb2531e88712ae0724f50a5f1e2a22511e8102d543fc94c92738145f9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195b75bcb4aa54e80bc00c62ae466a3c80712eb91f151eeaac7f814cf297677647d5e25b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5e35de738c810b0133106c34f4915955dee40dce4d6f1aca6a36e197b1c8d6e8281a09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19502badd7931624515025c119d1880577bdd37e928dfd8b4d3a841570810024d3c99ad22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe128ffc4fa9ac5687356165c7bd9d193503d745ffbfdae65a010dd828264306a00fbc87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20a2da93aed246b239a48aeb989652e8e91658eea6414c9989fbaa73a6159498cfe3a0fb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5870df80911a66d89c83d6d4d4ceccf182c479fb8d9f1627b537dd3b3965eb634a27079e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h196c84bddd950d2a02cb58f70dd3c7a340adc3f18f92dfdab0f01b028122e264673851a95;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50c4014305785dbc810eea340e34831b83b41e077546bca51a57ec7fe2d6002218a8859b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12acd68cc507329aadfdaa89f1aa26ae86116e61faabbbcbb8eee2b80b9b8dcb4385293d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1706d82224f1b3291b8be5543909c83b3eca1bfb489cc5b64f33275165dd2c8a008f113e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d201b3350d97dfea13f9bf4515d271e278140c7268b90eb742790496b60b86d2172ce028;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8430193749cd8f9cafe90eae42f8ac2d75709f2dc99eefcfc581b9d0a85fb82202ba94fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6bafb180e8fd3d4a0be886b962678dde84e42a20174095447a5234ceb40a588ddc6ec47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11823db9db7bfacdb98506a85e38153fc729e47e9a4adb1b13292660e1410cf96041d21a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a02801700959ee6df03aed3399f5d2e2d6a229addd754e5e7e267973af71be21a0cb035;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d968eb435db83fd877d597b2efe22af01384f4bf4e73d8b2bfb835fa2509f039a2e048d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f86e3b5ae8914b473fac1e740665174461f16cc77d0f0232a1ae242111d9fc16e4beac2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc13dfb5536c05f54447f6350e1abb2dd5a7fdb5cf8cdc7703a1179cf7494a6ceb7cc37c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9280b46df6dc1e9a442d300a07ea9dc092906e04224598108675e69354db92c0022769b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc24dc743af03d60f4307e9537cf044bf637709483cbd80571d693b3fcbb378d5e265d552;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he5e0cdb53924d52bf51552f2decaf82c824ddbd8a76bd0c23fb720186814f0906cd0c1f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e529e39e6b2242141aa4281633f60c7302589d68146460a149375dfe33380d9d9188e1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha86bf4c19c8bbafc45ef6152d11fb73f9cf29b153308bce252ccf7e0edd3d5529ad744eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b4e43b587dd4e20fa155f4e516badd69f6ae4c92396967047360bb310ffb46b54da2be0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162f4e0e81109cf861229c3ad964e7a7b82cc9f4300ec1607f85db924923f65ca9419d9a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54ae7be49323047974128e1345d0b44d1d42ebd89418dd9b8727e9eda74c4ab77b9ae6e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cf4036bf1ceb16fec5e98685f9844a5e94ce2a4f29361e1df423cec73bb444eb09842fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11213995e0c32b11110b2dad0b8265640fbd1fcd3053ad1806a208d65a336efd68dccb163;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff6bc718a5c8a1bce8b8295b55724294e80716e8bbf7d15f6e33a291b0a4b3356f78321f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1baa75bac90b90963cdc410b11ce97be917381e0aa5f5b52595fd563503693208aff604e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7f0d49b330681c5f5025bc75418f9c494ac4c6cb8f1143894b1ae58456ff35044547405;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f0ae0f59eb7fea98d55ba60e9e4b39b2e5060986e1e8f608eee2a58e9b0ffad8365705d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e5a7f56f6818ad54dc5e8f67564f206755f1bf2098dd6d35a1f63ef9cb2e356313c7dca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9930c72599baa93218307c77d8052573132244c55915e2b7d7fd1c26151458175bf6ddbc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9deac003d68df89713d0692f2d0935f0dfac1964be1eb867d61e901b45baa6db06eb6799;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h802f3de8d504eafc657c6a6fa0bb9f7e2f837939c171873fa999bbbeb21d3f8bb116cc4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118f927c0d12cffe7454508d4d359211f8c4fb2e6b2baf0f66e6d416cdc6b54f4d59a1b02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be72812c00886106a4c64e3fffed872b8091f3089b5000d19b29588d0d165a2d4b698624;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c58f4ee978e9d7267f7c5e42b9a17085b58b646ac70d6394f11ff205141ce3d7e5e7ea8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h729c25bed5979a746cb251e2d9b70d8dab52b5c6489ccf76f17005dbc53b52b588d33ecf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h31fb440554997122fb667045925f98cb92742ae143004850d5c91cd32cfa3c08a8b59dca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1816a1428122e287fdc521a8ac6cad47050c9018a213a4019b110f012c4f56abad1daaa8b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2402768d068e93762de36623175d63b97f0b3b437f87cfa208ed32be8fa74e63863f8c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h75e92b82df614530182d8352c870bc9050b6650468fd86eb8a7106557f354fe19da57f2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h418502bed44c03549f801f87f9be3b1dfef823c7f6616cde2b12e49c5e7ae770aaf6dd40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7fbcc5e58aa5939f3ab0095b4acc5101aab6bdf595723e5d749003518ad1a3837a1cca36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132769a279e8be403177bea8bb873f3376c14a48ad29246db3354d1b685dd3545dd4fba0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf941561ba536bb65cc6427baee6228898204d0e9781013246e75eb071b18d4f487f3514;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b275b8b2c5e03e7459a6c1d45b22ff4bf9ded41c17834e97a1bf1126d0173d0096e722b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47a08c8c078bab7ee2226fe3b50e62d61eb25808dd48521858236331a8eb382d0530f0f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca45b446f931842183cab2e9ce9b97fd6308ed957b7e011d298da581b8e56068890a74ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f85e42b8316a31ca2f41ff334b522effdc6abd7f65a56c725de09e4c3fc874847793bd4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd4d30c9ca93a4067d902197c3fd762fb612e86008e02e71cf55c426dd380990f272aa255;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cbba74610af957c795686bce217b43f0e50d95761a2d14178285777799b8fd1890cb5b2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haaca19c1fb4c64eaffbbf66d4c277461d47446cea521e5d2dbf45625fe286ae3b354d2a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10be5871398679a18278c1c7e0ab3e45827e6eaf25a3694ee3b3042b3a8024b56419c47b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b7d45e4b8626c4f81d3ed5ca99ddb2512a90fd8e93a208ac1cc0c54d2a3288278f47a0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1841ac50dece31fd90e0477b8636dccb71a4583655d7639b2478d6ccddf7277b3521c8e65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h29c3c3b0467ae65fe261181d439633080749ba6369ef3ed7962554317d0f89879bb80b8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he6f1a916dedf30b8cc82fafd7d27243fc9e939dd9ce026545101c93b3ab4d7b6ce175acf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e462806b57a6d6d4e48c410a72a49630ef0abc36c5ebfc0242765814d578f6d97ac7ef19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5229c398ab429d1affcb08905cc23c2eb0da941b365fbaea1368e7dacb1bb5260742c6c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a2f65d9194d6b8f225aed37fbc3d2c30b71e3d5bbbd540804393440af10f319aedfbefb7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae511f71cd64589219f97c4140ea91b5abcf16193074b8b76f4a3a8fff56f7b5ea45589e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1080f7965c3e4e23b9d1de37b511bcdb67c47dc4f404da6146587a1b86c1c37d27452a21;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bd8e9a5f02330e70e0a4fc2028279db5da628dff3b0c712ffb98d1e7bd0aad617680c9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe469b61db7fb33f9a4dce2b027a5f46c4cb37025d6083da2b78f07c7d564c4aad30257b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he2a180dffc1eb53f8ed9074037b1e99cd2c71ab1aa0bc016a6eec50f59bf4d2e6a355ab4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2eb3c63bbe76b6796d4045f824f7a52031995a95d871cd2ca1cbc0f4d2e666dc63ffebc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ebe822e8a12034abcd46d9b05f38e591fd231d3a69ff8340d104f56a8566f44313cb616;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1faa543d3e65b4e22c326c50c9dc8b7c5b12d61f174eb3571b8dbc606ad0fce01f576e5f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae78b9ba221e94b99ff5e2d3adfb0f5e156f6b6429403d7fd8b72e80994c4a4e906c52bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1991ff67b4230746be60bbbce5c79355fbf5d1306cfb98012b5b713db9bd853755a58e77d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fdd3abfb274a6d9a390639b56599d7cbb7e76ef945bd78e2d352d6428bf8e846eebd0c87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h551c2e74f1012e55d6b00849f153f402de063ed50640f49e9bd54dfde2a6fb40e69068a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1680037c2fc1d1f633ff6c05b250efe9ea459110dcaf1db2d12f893347821afde5a425570;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5eb438736dcd17d361f978883df57ba1bc257363d8773a07dc459b27e277de10434a5542;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2ce9c55158e17e1de11b0bdc70c2d6017b292017fb00f1520ffffa2a5a10ae481e908cb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1512b36c0a9758ce5ec8eb159f07d68c45f0e49c05ad4c9897c65f3f9603bde3b42ac5ef1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1208629d9ec14f7d6185ca5295407d7c8ce905f70148d65fd08607165095e3e030f1b1c4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d3cb3bacbeccaa2da62a3d94598a1fa21f40a2005d88bf4dc4e4161a2e70c0e31104e3a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af576c8f78bf45e4c61557f8eb64ecb19ca2dbe7187dd29725c4577ead04af9bc5548709;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h552babb7ee037af4cfb042a7389867dcddf3e9f2004008c801f55c7cedd5f072551f86bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4cb184db1377d58dc3f60d32fe83a4a73c603fdb23e42a127fca24132cfca3cb553e2a23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c1811496b53264047a7070df96e6081dee5bfd86910d8f3a2e6c9c672aa32875c23cf60;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7abf0d8cae7777860f941f3e82a7b01ed3c99308ba98eb7b82dcf2546cd56441d23a05f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he6b8bde50610570357d9aa2165aa1fe4cf0f6031e96d20f5d8580a55ed2e859d476a2ca1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h44e4317ebec1f11cd508503304124b85a804cb8a19bd3cb49076b436244fc1c625e39ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144c67a310cf19bfe4bb8c85e117b73308948d65bdff5a2ae9171fca2828b425e47c47a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb642f410410c8be6cbec251e53b995f659059566462bb95f7bcb26d9b9bd028f9776f067;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ccb2465614ab2f3bc0c0ab8f8747d0458ff293781c6f19a61caaa286d9eb60ca408914b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1464f6decafe1cfd862f13cce0f837af4dae0c71cbc62d40a787a63be58d84724c9558a13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb38bc469ec6cc83f188095e4eb09c3defb356d1608c09d39b5fac1a81fd75de5bcdde49c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138aac9a8476592ee0d89637ea8e0a3a40ddf0dfada38997d7cbead9561161a6be7b80867;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ecafc057623d5d4dc85e6b648fa58bd02c54de0f0e35fb916718e51e5eb1daf00d3d805;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1affc6f564e955cb94ae226c90a892a2f9cea8fd1b7f0ea500de2df1a7463453b66c6fe58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he209afd3c9b3e8a8b432daca47452899077dd763a62088752cd8afd0288ecca413b01fa8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17cc96b66ee6523545658fa7a038c2008002d72ba8b4f1bf08c9f41e4debd98ac6f7c976;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d449f09bf0bd107dc9df463a3c83d8bf7d6fbd3084c78a624a1bf336ab8943d32eee4090;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8d0230cf895bfcf6b33d09075db2ee0406cdd7e3e6db0810f9eea0d5de04d81e9e36a48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189df95f5a0488d525bdd34c890841c4c1daf4c9200663a9de96b105e8eeb5c20cb57d166;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b69a1b76d762baa2c7f1da5b5ff6ff10b16375debcdedf6d68360696cafa0c8a6a54e51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heea53b4d4ebf5d80581b3aafcd576c5039665a0b70798f6b47c5c97debbe10d7bd54f7fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebd055b0fe72e6e2c1260b75da5b3aa9b1ba022c977f08b055787745a5daa8d14c4c0fe8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ceedafb32ad7eb069051139eb10e98b403d188f176d44f512a49274f922e8f5851717d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h127fbf28ea15d69d4736d8e206ffc14e83df2ee6f90dc4a6ad7f018c37335fd259ba5210f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had561224234c0d935477aed640efac7bc1015f7101d64025ad349485e30f8e06efa18f52;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6b5e0d33bc0522216e5e6309852141218a6bcaaccd13ba87bf8b1a00a6812d9b49275ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18bce377f391bb61ada9675d07143e0a289f2bdacfe56dcad78c4dfec2645512f7fa70688;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6bde4061469455869606b553ceaa2905bd41afe9d440c7b9c7fb3a099deac229568bee72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59f6601d533b4086cf9b13617cf1bc7caa75428df9fa517741c0703e23fcd4ffffc4d617;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1854f308a797b81623d837fa5f3fef52a146ae7273b636c607d56d3af946bbdf4c81fb9b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf35c3e0295a36182f313b026056b892632c15e2fc3f248e61b4c30d1a1f4baf671bb83bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda0b1350514801fc03c1ea2b41fce487a2de582be5200bd6420d68207095dac218695215;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h823c28fc3f868a36c52445b66e4b58766611036fde38138067968d43e5274b91b665b987;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8fe5b3ea2c949bfef6cde727943dd169f81d995739dab34f40b4e4f2f78875370562a5de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6cab976f8f494197ded126a5a05740f61f37949ea467a4c407b270a2afb34771c4180a28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h915a6271a43e9d5dbc01838eec2207b9321e12420767c6935ee49ec97a8e68955f4baccb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h864dd4c94b36ac73f71aaaecd254dda5c4b0732034266a2af96955b5db0db4d4515364dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16fb1a4601ef25ff0811013f6f31270dec2d1f62216e1b1d133e471213dfaf5d9bf110cd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113a24aa170705fde397f3cdb8ae1e74c2e9c7d46c2b88d8698ea2a6e9927f0b8a6d3437e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd2d288b4565d90e10412dcf1f519418749b2ab1f63fc30cb95aaa30cc5844927ca428f7a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h96016c7e6dbc29d5c67009a05fae3580a075afea519d842b5894164f00bb2c96564174ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8856a7bea5c0d20310e01c504e5163414eac015027519a7e3b09ad8896d11b19b40543a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b80e5855a133b5c462c6cc097de652128c0cf5b034a6795541b75be4e6d4f93919014e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdaa18aff1ac5430d686be27bac5222b46e4a258baf55d9343751f37606dcf2b6459010b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63964d6aea1816daafe5c0aed7c769264e7b847cfdb58cfcbb08237e9d38c8eecfb67d96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h917b23f9179d63883c4d4185ab2d6b321cf5fda3bf297c79eac939820a659a2cfcae90d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10beadf2038ad4335aa580c4524de51ca47017b74fbacf274916e201ad17914d6e999c10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha62a270062ace4bfb31f6dc59e25e7f8218cfe3b8ab181fd3b8eae5d204171deb88cf9d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcba22819cead759f46906892190e1ca4843cea42b1e5907d387fc65a14576ce92fc6c088;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd7f5436d9017d28bec94f3e3cd4ed5e09274985836f5f9b761147d3fdb9e09ee64f73bac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38df98892c6c2d64de4fada464b2d0111f960e31fa7cf3d0dffaf5e3dffe103b49d0827a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e85c24399193c1dfac67044fd9a1f53c257ae622dd993ab66e0e484197cdac4fa872a0f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h655bed5f487379f7a3358d6f26e5a46014690abf7bb5a0a71db85243e81de9d50ca6f77f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd9dbd435c36a3fb4d2d5a1a27c367512e50351ff6d1e92d88745e1a03c22e2cf2540431;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c28873fce55741598611bf3dd86ad0e04be004b520f51e87f872dc5d9283cfde7a38282;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec1bd8254fb4cd04e163131c34be6a481d172499a0cc3d28bdbbe535207d7001d7131458;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14feda5283991b4d03749ba7d1f3cc2c3b11ae67f4f91ee1d3ab1e3dbb2e3d320905c337b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h130da8f08535650ca93e975cce9e877fa2edeebbea41da6c5e28029d458fe212b72747ffe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16961c4a6dfdbe8c608e501809703e5d8eebaeba4dc4ef65f8aa9ab6f4e6fe46b059d2bd2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1033af95b2d25c27f3f88925e6e3cf94eb922b68696be3e4bf29242e94d1c7e37624b9894;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a2f2a788cb0d35f19e5bb7613ec5817b413053e4a2ee0b386055aa17ccc285d3ac358b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h161ea076901156d1fcad26dcbf4a5178682fd3f1aeda11c452b9884ac23d83ab219d22048;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1381e8cf7399a55c454ae319591993e469f731b92db05a57be27d809cd71d3aa605b4c0b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d1a94eb0e39a5ba3b2dd9cc4b12bfdff1ab1d7d200a0c585d7b3fee7c88e82bff0388f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb375ddc5b6b2c0d1f284e62f12272d22dc4cc113aaa5aabaf1dca86e8d5ed7e2ad526170;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a27bd2cea8c31e050772dd225260f092bef8942b35cdd06fafd5c84d6199e74e778b04e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d2956be36861bae712d324ae786a26777c46f75386533aab01d39d3933833a5e5b836ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6780bb8a90f403f436098843dbb4f0332b1d5ad651872bc153a6147d546b31d6975d33f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5aa11c1f4b6dca6d47e668f8c86b89d67ac14eed42c2c234912616f1f88addb3b8c76c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74ea68db3b32a051a235039cecf72c8540cecef72557b8d41ba28adfbb8ae819ce6ac42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb062b81b11bd03141692eed18e5e0bb7643566b2167b7cc3aade2cf0f0a19874d743e819;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11197e85270b80235c7f8b73307e4cfd7f5a6d733e8ecf8fcccbe193f946678a024450cb5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h103fbaf0cbf7e97f038ad90cb8f6ec97e45e42c3d1c9f6cbaebe2728c11cc18a326fb31fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe6564c4adbecc034877b47f8a59565ba68b5b2834c749b34434228d431c8689c43916ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16071bb47309052077b9562d04a28e0056d8fb51a44a3bd3d7671e62be360069545124aa0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf366621f1438db298ad824f8cce2f23eac5c19deeee781419377b3396c91eca23c064201;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13bc3d861588d0d657f253d77722c87052b9f1d13d4a5c053c5fd2db9f2bedcd838dfa1b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136e233a93c4e1a3286249bb024692c307884a218a4cc1cb5d5a35796f280696e0eb4d847;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1169d28b526296e4582cea5294eef30cbe4140f42dd536c876b59abcb9d67f0c15e3eb0b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17bd3ca6a4ca4219415ddb5f752ec10357ec9b250003382ee0eee4fe540c91ba0f5319a79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192452d0f95c095f58f347c38f7a8503e4e7ae250d1a582c39e8f63fe6f09386ae096b208;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1836de5b0f8da6792c2c637bb3cf4f592d940625153b74242fe3b04447d436f71378b1427;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1447d10cb17742e628181af9fd3a40933efd19c60a95b8c1c5b60643f5bbee5a6832188fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13650cdfd87f27dd385b5f3be21c36784e827f4f767cf37b2f7c881b0dbc11154df48ac15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h438cc3a97febc8e29979339da52827ad84db4d999605ca92d79179107ad3224d08929c90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebd0dd5379e61efcb495db92c829e7693afb11f612b12b0ee31e1690ef6f2ffa0c9a46f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee2786c0470e652bafde3404eff41e641077a763b46b3fe8a2b290c37c55a6187a60a557;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5be04019743167773ae4d2d37b6e3752215f2d134435c22bae00bb2df41b2f8579569e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa8b2ed95a7ad198ab32c6a333a612c4c28b697da8ae6136ae987ef6f2184017170242ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h897419d791b468e9fca2969ffafb53f8d35ca1ce8af37a88f94c19720b12b6d3d217ccdb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6418e316cff02bc95436e92985844b6b30f762c70cdb2bbc54f1645b477529a87ffb5b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100ba9733be5a6e10b56fd0a19221d8fa7ab8059ee5b8e6de42b72af4a57cb578b84ae2a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63f11e834214ca42b9ceed9b17f495159538e949b8791a88c4214b149faf130c26a6a0e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h685d1c6e5f2234ed0ef2c86097c20cb763783f25d094e1131418be49bc7b59a2fc2b875d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb964950a9ebb7a23002b926ea3428d39f3ba2c1f81734337a00718acabcd91d6f867bab8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66ed204494defa604b6a3a03176d8d60d82db0117c12aab61524a8dc58c6fa3d6dbcaf3d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190c1e5346dbe9359a765bfa1b7ac530dd3b483bfd2ba24c9e1c25814aaeffb85ab169bcd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19df6c09ce8d85423fb59834009ce3a11356673f714ff5f150e2fe7a05ad69679509b954;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d98a78dc2e1e4ecda45c54d5c953b8c4b46589cd3e2e4de2e457f4e5f8a6ff5944c778b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3cc6cbcc2cf101f9f0a8775666098ea16b94f558ee4922479d4792296bd964e268ece7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e928a75156a43f1cc67f6d634d3977e643dfbff017c752173d3838c3b3935331886d5f43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h102b168c65b12eb6c3df6f6fc707d72ef904f50f9160ed042105c27feeb4806e42a3e34c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13bb892246b9d4cce378b340c118e80fd38f1ed366fda70882cb0f8325a8950dd0c8ac022;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8cb618ebe81b99f3010dd433bcf7ae7f138ada4f0078f57802ef6ec8b1405a359f57d224;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140c6ab393cf056c10061e385bec5823791abf0904a9a36549e0138b0238f6b72f17ed093;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b578196a3f90f8f95ce85cc140e43fd439eb675e7141161a09d2cbaf7bb1be457bf0590;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1639cbbc8b4fba82167fbf8c0ab0a6d909d665e20862a6b6eb07ef5e705141699067b1ec5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h34e9ca0de89ef124bee74d2a94331a4f276dc5df4c45546cd392284327a365a99eb9f0a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10e7697f3face13f404893f1fc158a5207d319abc61d106040553fcab472c453109185fd6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab1dbc06bd6a8a02aa531b2bdf6fed4802ff36f079f2f3881430a276a28db15b93088630;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113ed599f26df22c069dc28628289de7fa48da50f2306b54396eccaaddf9eae21063f832c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ec76e82319f46c469bbd0ae8c33da51ea5f60ed305deabed127a795e127d56595582c58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h529d513761ac03687fead872c0fce5c283ba6ce83dbe69a568f8f35e670e4239bd08b4ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c40f8543218762d8c6663708b1c77836fa15242ad15bf4f28174635d3315dc0bc7046e47;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153a1babb46b0ed86c60c39807bcc5a0dd4347b18f12cc535631863da9c1912c0f438d2cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c93dccdfd368e5e8cbbb010c78b81bacd0ab05c60731b7d5e8ae7703853b1cf7d93741;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc47a348b9a7eecf878f4b898efec11b66b31cbf94e068656bce96bae805a9814ce51c9a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc1caf97ad0422995a99ea4b3394bc3b52284009578cbe989adb3f93a84af6c346ca608b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59b06bdd9b8e8f722f91e07b98788994d2fcf5b7c509a62e34ab0b5c0fae74ca42acefac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0d75d47027c199539a1bb9c5a6f9f0d2f4f3a02fc0841b2be2a8a95c49b37094beffdc0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h53ed46f909961f00177a97b5e89935324501be3bd75769b2e4ca088759ce315c3cc2a9c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1758fcfeded44cebfdb96ae75b24f213b23f1d5963534950ba472784d9b4929b81f2c90fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3cdf1534847efaca79770b60bddd40ac7376175422353d6b8a1aa5a3bfff3be7973ba969;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h83d72a13e1cc113236db96648942f87884c0559aa29371f82a097592742c3fc378be7490;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d53368542aacfd6c0cf167b245ac06f74750e5fdd4fc01202787bf12f15509321b58957b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb2f2cbdac1697568272bbb2926278704e8c6408a43ba2bb0fcae10f0293a3836227f0238;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbdde72cb9d791eef02f2702cf5f6b914866078033d4d161a0d17f3e0d7a26b9e43ce1c56;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e77435d0d114aa23a453e83973641be6fcea718af339aade13c56d8dbc3ac3ba19515419;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147b0d99a97ae98144aee2400595940afc7eded599b22831b5088f044b1af57dd6fc35a85;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aef741d882879ba0e183fe586c7875b9626ebaef9836e5ba304c3966843a94cd0fae0855;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a2b863b941ddf3b2fe5978e9dba98a24b5344036e728d7c2799d3e3a5270531389aed4fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8ed4dd2250edf2981df236a7907a0e24fc7361c3860fb718526a5aeed7cbd925da4c3184;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h827e2424ba44b5bb2ced2b7c084faa7b5d46fb74879cb43b9373b9bd1cb8849743f4bde3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8956ec892a9911b1d572dea921d6101cd9beb0aedcc8113af32064e64995f3fec2c4ac1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec64e634d26452dd8286c39fdc707b915d9abf974d49beaf8ce4ca44009dd64a01d8fea3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17512c0fb7c6051f165412c232759ffda3f5ea23bb26dc05e81fe82087d5245769df0dc3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h178116361c7fc58524573ac6ef68e3a3dac4de337ebd9b4d433434950295b897f9907d14c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1894eec170a49fdd48208af2063738329825cc98d284ac6fe003bef7e244f7f8a50d499;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h70604a94fed03a7000cb4d3fd285b477ae0cd5100169b60d7139e2f1ebe9a327aad3ca46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfba24d716900c16128b646062f4740bce502f5795751f76b281953f2f6c8084a7bc58b02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h895ff006ec7f7a2e48a7084d91345f9362392f99f6e09c1594ad310a8cb1ccfd94d95cde;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1796f072739a44a9dce592d72e2bbe763bb8f5cf651f35bbfe0119aabace9f94ee96d3a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h442ce35001eb008a4ed54e84a6237c9c6a198dee5bf13d11d59252f224b1b99a280718ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a9ed4477e9450402f67676852cb4e48f63719f73b261e13c61a8bcaec8c3c2fe8d3ab20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5dbbb16761bcbfb032ad08597202edaee7b8a2c3e8e5a0044bcf5dff4efd0cd28ac73c49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ea99460bc4ab06f175177c972bc6e6578bd44ded876b00b41ea1d1a8c7745e1209fb9845;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c06d7269efae0e10a3e723068e77725cbfbc30bd402504071e486ed7278b2ebde67a112;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8665857744bd922f7e3cb265463353c6f8b63083cb2debfa363f2b01011b197042f6d2ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15159d4cd44e0c92db55300741b5d242e3fb900da3db569d6209b3f143a3d6c5e2aabcb02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7bbca7928c04b9549a67c2ee1c4183fa0b8e7eb93df03ad5c557caf1c2eb1b776e643667;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h29c0fdc287d00dc855b7de023de55e277b78b19c8ba7a47780f593ddd60b59d27e222065;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c88d2c52a1abda181529e5cecf1836bdbceabd1a9be7284de363c7a0af721b809a9ba6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1558638137a15c0cd35c56942da63a6da54b5d7e937e1b47b66ca4ede328779997ae58cea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3d6dad6ea61b179049e64911748f2f5ab92dd9a29e17f6727acb777dab0240a8ed18289;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57c6d145a69322abd7453b4d9fe9306b6e993c77ac63c0e251e35497d4a520cb0ca99b4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1134d0fd808b58e608b9be7119ec96d81eeaa0e18cb1dc4075c4a6f43d4ea7a26615c34af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd61bfbd80a9080fd8cfbf573f99257f81692d5957afef9e90e9688ce7d5541f824aa019b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a72d86ad355c64bf3269e9552344d74d6e6aad560df560e14a2e4df9554561413dde5924;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6900ce082373c0b3c28fab6f67ed6cec84e07ef5f605a7629ef61691e72f09ec581f0b82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a779fa771f2bb6a6e7090c25bb7fc2451b2268be4c3d47189ebdc752f4c5b0e33640794;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a584b58aee4b1ba2e164d19a0ae2733e29cfa67690968516f2349ca4ee41d36e87d640f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e760f389de58edc0bc71060d8ad8ab759bf5e9623d5bf8002e4890908323a5c3ccbe8f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c891ee836f36929c7c49fee4389c22cf83c7401050b38cf6be4d44f53b89abbe78e8fb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd370fee843b2d08788fa7408a0fcb98acddd3e827acb325def52d69387546ccbe73178f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141b89f749e4163bdc5c779e519bdbb4a4c10dbe0b0ea92ea2655b2f71dc1d9f80f667669;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h27c90843b57f0044715ad0d4dd6b6503aaef9be5cbb784a01cad905cac791924bfc593d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haba66dd9c66c8385e617335575ef2c4a328f634513e0a744d56a59a7cab94757e67dbab4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a43748d0032e248061f39c7f988f8bc437c082355266d1db2d7629a78daf89d17147d5df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e2853a7d13d227ffbaf06217d482700427cafed3448a64cfb77fcef021b861a646880c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187253ea1dcbcd015fb0974c9f02fff96ce277ff0a16c15bc86baddc6c7e455aa5f418327;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e62bce08b90c53479c0e29e080b973aaff125860e479e80683cc07cc5cb9e23bba06be56;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14073a175ed8daa096579cf10d00c4e1bb51f2eea6bbb908bff93a4cae4337d0b344b74de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4cb0616bc5d2bdcc1b41815d029f564e026d4358e4ad60943ba4c7c77378aabd0b8c17b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4af9b558ccb1bbcb6a69133603371f710f56da7e90ffa2f54c900f348c5d40a24b587318;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h367ff304ce5e06ce7fb95de655e6338ea33827bd14b6fe47a45aedb953bbefa9d63303ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7ac7502fcd82f57010a9bcfaaca6d1592267b4ba3b362ef3bd93a62fa5d482f1eed4f59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he86ae99fcf9972eca42fb35b9f733d090a63a4bf4083aa7581a1baa9accf1456a01dd44b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c13a6c714f11195e944ce13c3cf70431ef31851e053ec194cacfe7d3433df03ece4a8b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48d65968a1b3a5e74e16f3e221bdef58978d2b470110aaf3bb3da4260f0c333184e9e307;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f1bd7898d2e4a60baf08d4df5d2c9bf3a737d97c380e1c76d6f97faf10bdbc1a21f0eb46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cca5d5973fdaeaebf262b16d8655955e191aa0f357746eae825018921ab054ae42db3e69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138102e241fb3bdee17ff0b8ef6c6918154adc1128c831d64f956a8eceea72498cdba630d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9df7526f4f97face3d38a643e64de54d53ba8f96369f976859e2e9ca3628e01047d71b9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he893a3f256dc060dd435a415fd6c602bd0888a7c19ade8594e621f3a0e62e1166769513f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea783ba3a605fea9deb12172a05bf287a2f8a5aa4bbb27ba22d941c649072142b10d9755;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dea9eb70ddf09cb4cb24439e8620e45baa97debda8c5d72a7076f225196f13cdf5441f15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1994f4a17e36d871d0f55dc40c36efbc3e504969e19c10f26d0b4db58717d4be86928783f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2429c74a9692272874970851e59dc292bc5a84e3e9d06319bb4f73c2a820d9774214a19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8e018106bd3f106f9ba60d0614b3be800b457fa76bea092c52be2c0a22332d154ffbd03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fea1510303676d84b9fbc9a2df154259d34982a57e6659457f094f8b924d4b5daad297d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d133eb5664d126d2bc24d4da49c0400e6f10ba871d2524538167a38e5647953860fe4abd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bb8eebf0b81e1ea1d25822a50cb8ffe20efbd2215e2e4dddc84e5b6630df847a5ecf372;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1761cddfdb5f903bb34a25efac1c052117d039ec7d451a22a55759f425070e9d3826fc255;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4fef4c83fef0527e3d258870a992908a8bf784acdc19cae9a63f98bff1591d8e9460cab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6047b53c12013d98a2ca979ff8b6e2bead8ec4cf8b1020c14b120ac8ad67223c4a1c4b0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c085c41b917dda95a4caab220331993c23635ce1fffdf5358d35f4b525308100eeafee00;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d3ee0a5b3d5de19f316f797f768599d6ddcd5acf8d82cce8cd4f6a501f304692db3452a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d5c818df84be59084134790fb120526871040c152f6f3948bd543f213cb0d8f1c27d29eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b372dd6e2e9c6eb838d30cc0571a65be76b2edf04b71f2cc6edc4cb6086147e2e2dd30f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6fc4edf9bfa5a26bade976077de14693fb8d8f2637332a43d8140e3a6be47670978c8a32;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19044eeca7025261a2a5d4e9eaccdd6f1c1b644b7f2a74934bd4aa2f8051c9e0585c8b973;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1512e8f5d937657cb3024bb7874ea1c2c6fbb16a07ef4e856acbbd203ead57496ffcfb0cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10638844a2e7a296b996a2b251432e482b8f6bb13afa42b7bd6a04718899a473af0bf982d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c018c2a3b2f72e1d5d6c2f14722783d9fb385849c7025e80c3b01dca4187a413e374215;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6bee5bf081a9da820ecadccd2bcac09e43c528e2c68dfe32cffa2fded04b83b4473b93f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8bf5e26c4892c1ffaea08be45faed0d4a467d0376d3ba363b157a39cccc9297111aac88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ea823fcb9a6e6828d4c8b4f8964dc0dc53538420055612a5e3c66f5b2ead877a353722b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13418cc2b0db9e0b5d3d553889f2973aa752eb62043679180b48d566631269b3b1729bc5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7647e0a4eaa778b09ac33546a5b60a577666d19dbb4a1b8940a248cdda56210ecbf17927;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12a2ea291c54fb84da3ce20c6abc8f9cd9f31a7173859063a0e1bed00aefc71cd6755c86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd452344f699e972a582bf4f4e7968412bdccea4f8475ec0b9ef00ec664ea4e507331737;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3d30b0d84eec6c3dc31cb03c4b57dff6aca51ca329e01d26edba2092be8defce3825e944;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h31ab902b75da51de83ebd1e5e1223104f52fb70b6ee1be7279ae1dbc0427b9b79927b5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b7ff3c31bc286f0261cf8a8ea47f8371840cdb3ef0cb3945a9b250ed17fcaa4c7601318;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd4c3b6c7fd47e35e6de9a13095962c2606bb916036ae7f62dc9f026dbf3b291608b4e208;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76b83d51aa8bf8dc24677b2f186c7847f0824e12f3e58cb49e9d078ec92f4976e60c15b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba328dfafb9ac4866a634a548f7c9d217fadc093ced69af44d7f713796253e8a17626271;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3418006c30711a1a83c791fb2c7e813600650b3595abd08a1399422bf4f6e8feadc53763;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e1ca9ef9de7c37451e199f08939cec71c484e39be05e24bdc319518e23f89548841389b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1464c90d464696a6fee583ccc572720f22be454d2c747b6f5080bfa6df49fb994861d23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1106b9a6340730c8c681af43f74dae5d8cc62d7fb853ac4108366a718e8b51c1d5039fdce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c297e4e67028382c55ac2ba43ec9aa2110ceefe99b1e4297052ce559407fa832c2a4526b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bee63e1dba216e4e15e59b9243c296d905e5ac2b8bf7e460e4af0046ed0cfe8d02e4826d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1664f8569bc61ee859ad23a700adfe6cceb00f503823a2d3ed6a801c3d6c63f8dec77f951;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb70f872d8eefb73709c875e6498b09683c5b7222233dfeb916b5e361b712b781a51adc2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d2a74c839c609d0ff659bfc4f28ded343343865daf6560da20e6dc55623c7faa65f46cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b4e71c50e2a4aae7b4fa6eff36bcfea1f99321edb3bd1e4e6a296435a87001ce291e0bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9274b0ee571516c773da074c699b11566ff074607cf391b966d7c7b323c769969709a1aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1572039a8d3c1a5f5627aca09393fe9e567ff499494a9c66e0c07c2a736a727d46fb1294d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62922b4a51c7d9316458952215039197f9b8d54cc80d1fb771e8250a4760577e688ac6ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h720371ad834c8d6b9876216d64693c3bcba23b7cdbdb107e9bea3379490423b736b40c5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67f7681410856912a47917569fb6f8f11f5fb791e36e0d15cfd13a95544557b28bbba29e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1240682cdf3b76ede304feacd8553ead6fe467409631c828351b04741d84054b0a4589947;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8c4bf918dc27752a102365fd3e14a78581a6a1d1c8b9f7b95d1b25006c0761b7c4d9d8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fcc3ab40530bff32b453b07374740725eddbf0175f89de3f6a60231e71195e0fad6890ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a9347c4cab1b4f295ca828dea48a20b1799f17c6ec2e52e6929e7809ae1d7d5e2170169;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha31ec0953475b770aa46f9eace384c0c642259251ea5732d100fc7a4174bfc5ed4c0bfb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47a771ab79325c65f822dfc96e9d57c56362ec6018fb02086b45a2e897f921449c00473a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he49072849d19985dd8174b140a57b16c4e968e4064e34c30f3c2781a528ee094fd76fac0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18972b02b99f4c01ab12fc380c8c5b778e5b94ea55bfd2e73c0a540e52a87a6300878b153;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1343bd972b9f334dd76c27432dc9a42477e1f9f29d608e2a34a251d53220b38b23a957c0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h108354806934bed96122b64dba1a79d4f1ad2d7884a8cb89f5432dd811a6b136d4dc9f4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf14fc6f7d5fa9dd5cf84e955a34967d91e60b6f15b9ad952276f260f605bc90cab5fdd95;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2e8d93c68d2effeb8c9ae4084c8c0c9b1da69d73905f2fab8b485435c3e62d2834effbe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9db42f86bcf1f71021142ec5e94e09db54d2c82a75fcbd44afdcf762ef5120283764d69d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5791b994899e260ae6f488d8f888c35d3693efd0bf9927be6baee2558eb2e90c3f7029f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36af2f014a3799f0a2a3009f658b0bb58bf558bc0af140cc72a186e7018ba2328bda15cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3fd2c0428f746dd41bd09d3792dbbfeb03ff586f0d9600d66d8d88a3648cd4e0e5334ff5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4500704479993c9a1c6c62a078f943948e11fb8ba740ba4a62b55c5654cbe255ac6dec88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha5c7d950f21a3b5ebd9445f0189d2e4bea11ea3a01b2e9bbdc25ab453c5b37340f018738;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h102d3188bf6ef08bda8c742e6f55493037b4167e596782ce588ef85688b5ea8c22745e5d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h236ab8fccdae7ca56dd0c44898b964b806833fe0275dceceed0014c7a69053d4d20372ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa578a0622ad79246dbeae709c78e1a9aa2eeefbb98f5ac490f1629f23a371b62a47fb74;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ed0b62b3b5bb37ee7c3c6ba1fad932b44198b5dff04dcf18da6944da614e85f05e95f46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1338a52591981f12c26fe0c0d847b540630cfdaefcd464a29d6fd455f11b109959194424e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6520f5a3ecc9719d395066b01fb29badcf5d136851e284b85fb505ded3b9d676f036042;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e0fc3f013f96fa2a8e3a7553c8989be1623a46ed8ec9e277bb16277d9bb30c5f9b87c07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190d08d81e2d9749ed78d7af2657327c1d5d2fb2b6c589ad6c6603811e5cde575014ae834;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7048230b1b6bd671cbefc85b5cbeca86664236c19e33cd93c4d005817cba416508aa9462;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b6b4bc8e5a5d63eb3c45ca247cac9e2fedd4c42ceba968850b036d3c0ad726afe7f2923;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h558f319078491d6d5c6bbc48c152d615e8b41a19bfa237de72b2a6953b1ab8edd1a5cf9f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15db920ea804b20e5d63689a952ab3d1967f6f972601327a7e5431d53bc5f89508b780a08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62e726a425384b98dbb3bd41ec0cacfbb7d8c476fcd2f524d2fd3a344cd6b237953ee970;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c4d4ae22386fa4fd6709bdd09963a654d5bb7aea7d3bad66083b406bdcd80d54b082bab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1750b933f7ebb78d02a0f9e903e3888224cededb502323dcfeb3437e35b5ff4ed59c63f99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cfe4494a8b8604f3b6b15fa2160c6896be43116693610790a517af7555309b3ab8ef80cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4872a969c602dc80f0e81e0775a71fefd31be723bccdccd67428fe7726b0af58cbe801d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h84fdeb6b4f23f09eaaa44f02ced969a07fa8f5406c53738f873530b88c79818996e7045d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h169b5b8de0a343523807f27f1d00f958bf2a1435d2eaa139c24885c98d818fa49c7c34c09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4087e2a84b1c54300f9a55f204b121e17e37b8e98b3e01196a5ff0cda27c40d5a7bdd2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c3140283c3ef482d488b36a170c702dcf84e6b5223207f1a71c69c889a39373ceeaa4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h99734a3102a421204811f64a740d1acd6893a86486d7922e751079a0424fcd011f5807ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf60e3b88748e5587098391d72c00b1726dbc991d7ed05468046fd726c90d59d47734f26c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h241b25386c08b8719736e78a19aaa470c51ccc011c461aabc6f4bbf0fccdbe4a8d1bd6d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c258aadfe7f47fb83d089145fa29f51fd4effd413606010e6358863422576c5c48248fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd4d39e639fd368dc299ba7419e8a22df59c5140286e04a8ac142aadd392fa5c84f75ea2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d86de4483f9a3a3ca2cb3632c46ba6d37750d13cdb600a33eac085ac411c9f673e6a4c2d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1187de5ce5521e6b98d30c222c042d2c45c30931a532237c7933aba0fe863fb0f53eb6a3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h106e204cb99d548809c8ddc0ab6c2e9be0302a4a1ab4c2a9d51188c672ef2ea586f46ea94;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df99fbfb10da793e91a7817263300555f0be12dcc70d3a6d2816e3e867a8e9562eaaa0a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6890db386bf4906433152f6d875b41c02e2e76d044ef178ec789b5b02203743eafb39248;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12584e7ea582c695ab618c901ad45d270fda0e28f3c9e399d1c1e2c69a4200803dbcdaf41;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h483acff699b548fea43fb9519b97a022b5fa7fab1c7bc2899ea6e9b72587c0e50e994ea5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb17e36bdfed08fa2d56c5b2bd040f07046f247b0d08135dbde581bf98f840fe951ea8355;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a0b94e6ed1f34a285d91923c9605f4fe08aba751d36c668485799125740fc7b2a9f058e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133a1bed57bffdc516ccee3ececc8f06043f399eb07571276b0cc660cceb80babbf06460;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h360f58fa40903b30957415e32fb70ff6a74952d147c18e13d137a3abcc9b5c5f06b090c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea7473f8e8f0ba0fed0056eecf610d742fd969a1d1d5542c8a90405b0d85c40eac6ca80d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b78b6eac65c0d60d954c2e9d07335c8b01e5b96abc54d8df4583bf32069db925ec010e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e0f6a315ad6f016d4d35af064809a49ee97ae229f16f62a6e16f3b6ad3d4868624cc27a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b31340669cbd212632958c0de462060e4cc8c07715fa0f4ab9359dd881b43e14b3dec6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6e0461f891862db299d01c9edd9bb8fd45a6e8fcf91721aa8fbfbf3609d32b4b7d03b27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h271b2d8fea4d7b6b384aed03f2bab7fad669d8acc199bd2ed2cc3260c779f2e3d67d99f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hce274267ba0633eb30ee4aa9faed3911cc835b8f18b8543c935ad96ff6f81038e305e865;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1432b931f22241d5b171b00687f3f962b8ff8040dc9718f96f0e6c6d36478f3bc40cbce72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9489439f8bdbd0548141bdf334ee28400af1aad6a20127eb605582bcf57c4abdbb9941d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd33a0aac9b0063ccc81970e03508f011aebb93d0e727f9271e39dcbd648d360c8bdec991;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7de547095f2684e33d0a43db6a704d93cf74a24d988661c2c264e616f2418783ee5fc809;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b71fec7ff1f6d5eab8703dab49696d24dae21f2e9e02fdb93cd9aafdaa323ab1b38d97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13c5497789efb454a40445b11b38d86d09d87dc5afc726143991f89b7006c1f3ef85d0f16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3faacf6ba9eb3fc515e56056010ea0d9403cbae460e3c18400caa84ed094b16c6110718;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4480779a3f21043eccc606c601e9c1011396f9ef5e85b72c56a069026401d913df29668e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b871a28ab596ec9dc1870f8f56696eca920bfa24e9ee359e9ad7fdadd5d6edb2915aba9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16433bf99bbfe9a9775b398a3eeef382a75ced818fd8bd7f28e5ac038ee9432f2aa374011;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6780e6896e29573a270f8cc59c92037ce32e1463b3c6e83d03aad8fd597c4d90ce61e045;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1253574e0890beafbf3d1652d99e0a68c66a6d2e02fe0a9fad9b0ef252fcc1648e976dfc3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8cd9a2f24a43baa5ffdcd6dd6d61319fed38d33fb3659a1920afe7d4cd198e1aefcfe847;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a14d9a291c3758a1f3c4bc8106287490e24764780ca5d9ba94f3e227b0c9e9c92d9cb3d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h795965c2cd2b8e70e09ba18ff16003b33e211eec0294f07a76c5b03ef6bbdd4b0f7faa43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138f9768a335ca8d62d3ffa31b95e7f75461cb7e39f0d4d01abda47e4fc4986860c98385;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h374bbf1033011611b9f179bc752329e8964f74fd6732de5c232ce141c7a7bcbddaa37bb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143c2bd9562db5847afbe5ee53d36aa07ccfb193897260e21459a54aa328244712cfbbe5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4fb5dcbfe2aa976d109f017658d7f9899605ed687bbc286c0615080ce4d0733168cccec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7ab1ce56d30011809341b306ddf66767d03c92822b9fe347ec6a04743e1c4aa6ca9ad60;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db610bfaa11d4355c161bda4b62c92df0633312906a6d17881f24013de37f6c0cb847494;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h484752b060ec574598025fc97afe75b4c16232be6da605f3c3e16b630ff9d9035ff2d8fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h186364936bee6df6747e454ba6034bb3cd6e408203be9fd9923732cb189dae188380c7f53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h674c6d1d8a3d711ae3dedb204a33f05024ecabc97c1f7cec6defd9689796892ef014a4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23cc4b1f14045c65b2043277e0afc27a6aa8ace1b9075bceaeac004b614d894cb7b18002;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72db40a2d2d6557db18bdeaa19c27079c0b4682c71f9421140aeed0568cd9f6d36908055;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha39e097fdb5708e332d5f27a893911d52c1cef811ced7cc8cb37972e2227c53cdbc79fc6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h68d32f235e232b122601bf237641ff50616e856d1623ef677ebf7f9c1d5bad19473e88bc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ae82bee127c74e15ad0da8719ffbda814905abeefb571039aa89597c8713c624be3c25e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dbafdbef68f164eb080e1f2bde52b3c2d3f98f4601031265dbcb6ba438ddd90ff192a764;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2693a81149cc6ee64efeabf8e7fc474021ce54e39505ed871a88a0d57658bd80dfcbc78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h752a473959727f5eda6bd3597f1bf77017444b4a64b5c55849ad9d1448cf32176ed7f56;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137b4372cb91c70e6eb0dd2b48079b60e5779069c39fd4920b12da2124c0c71afe8927988;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49b27a119c69f5af75e13b480c8bd098c40f429e9d65d61af1d3fc165380eed1204920b8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c03aab4d259bf2c7a381e4a00212abb086f386fde23c6e00af4bf180efb95e6d6b07dae3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3df29c9e5a848acd507f1ef39a752ff7f1290f137cb80f00d294e7b34649277d34886f16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1154e210de85873a40dbbfd14eb675f7003a21c1990af0ee581bf5bd164605dfc2fee6c76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h108d1aafd2d9c46a3b633bb38d6c17c87a9d0311c09dbf67f27231f06b78d1f8778d52b0c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h969630199603c0167d83aa710f6bbbe06297a77b285748f2b2660c96dcd1230ce02768cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dfb97130964a6129b9b2911a4a9fd3f4e51d690e0aed44324670b479641d1e2f75580f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6966dcff4189ad50093dc24450183a5201f2fc278977a26f7fec9c7f2fdd31aa0d52564;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h754c2ebcbebe30f25eaa118b2978a6c8c4eefac66ad3a8fa81f8aa47eda12fedd90d671e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b651310a9910da3f97c1cc1af50948f1d6d9c8662cf05630e2ede0cb64031c236d1865b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h924022e2a3898bda85ef523dfe4a18c90070d417deb9529321edbcd831ce436b25b1a206;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae49ddf74498bb3b7694ff457f2f0e6bac04a4ce93fdd243dbf9c3c38118967616c05231;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1873d6d77e7a77fe067e21651ae7d8d353741e8c8fb301af412e26be0ebe0cf7b7bca61d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ce3c727e0aa0c4cbc110a1efea030cb8179928b54c83cb774a6ed0d57493493df131989;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d54a89a0c9781dfe51a631255bcfb98b095f81400649548767c84f7c232d4aeeec14dd16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bec8a37161ea41d3832039a4bd684a0355a8a77f63b6d584dfcba09d6f3fdd919936835d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf286bb4fc0ed38797edaa47cb3511b85d3ed19f71d54186420420d464ccff4c93d84432f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ffbbfb0b4bf320fc928e115a942688e0f954ef5e5b74536c6dd3b5a01d8087a8f7bc34e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cfb5eb1b46f870b82c0849ca5b6c19b16ae04d40045f75c1c21cef3002cae9b8a5ae0860;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7109eea107faa9f60499f5f368cd2c02e4d49d54d2872b3574b635d5ba71c941b657ef49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h108d1bf8b579c88ed81def88d107d20bfaf151629823cee30fbe33bd542141413dd9d3a3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45992bd5003fdf6a3d2a9290727c268797937e165cf2da2e7650f26c5c55b45fcdc7f06c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f04b0998bfdfb26b6222feca250eeb844cbf2e522debfc9d709ce40e7ede413ff38bd7a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c32ec52fa230c661f952262a9d4e36c61e2388a6ea0367350999676f794a3149fce7497;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b27b7885e970d0dad03484818b52a6638c1ca0386e01e4416c7d854a100dad68cdcafb4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ac89a3400feffbb1264bbc253e3dbf397ea829ca0e853cb5f0c7980f940ca3d3295fff3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c9ce3d45138d1f5f02fa84d579b94fa4ac7b59e566f3cd2c96fe7b42ea71168d011f80bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3fd0e614f08a4960d21c23a397e2b158018946a6f5c219d3138815cc855ece06adecaa3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a3441a9f68573c3cdeeb76d2d33c5da25676e59ff077b99e1e029abac20cd93523aa539;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f274a1db938c8fc1ec4072cff4cea9dc9530a1cc1a8dd298ba485e4a772377f3b56f42ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9daffa103165a4b667407f541b22f200335f79287e864d2c875f1b29c7ac29be21f0461;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23c8066efb312906729dc6654d17040ef2d9b28bdfe3c3be82a8c6fc43497cf1b3dddb39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he6df4ec8c49a39ca6f199fe600bf2b0dae52b52027a36a275133c70b78e12a3b4d55d5e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b522d1c4418b3af108dec457870e1c0ec5ba0aab7a7e27bc08eb012877a10c64b9adf20a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hede73f8f20641063bd4d2307ecfdb090ac582e77bedee2121f8800926b1adaaabda0b9fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b8d6098a579ae347d798a747f253f016254e3c26e0b90ab9a6d349dc0166795e51c0424;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4b1797f4ad57e7a9bd72c3acf4a882add30fecfb13ed45175c10cf8bf7546bf065921d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7cb855cb8f8d6b32f1de6c07ffc0c2375e0fe77bb99bcbb54435fda1a02866c188004c33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fdd23222723f39dfe6064dc052e23938ab3364e16d498e6fab29c33ae2cb27d8d971cbc8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3142e956c144426ec96e9ef85745c2641c9fe0b3dab2e938118286356308ff9d0edd9e7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117431682cffbdd5389fca7218e308749daaa8cc44d6eab5510256687078d7ce0da2c25ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b64be02c9a307e970154bcdb4efb2c7dd33f79e994cc3e961b45bd452cf68871eca7325;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90c1f6f0223cf83a8f5fdeb0aaeadd1fd0ec1d7a153c710ff417a59517f0c5835bcac064;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48a72145034b4f307dc15933d8c05ff73917cccd67ce679956dfe35624ae9a6ca885ec3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10513dc4647dd8fa443ef34f49ba64df72cf49ff033ba608b3a0a70499d9c1978d726bc0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d7e5d1fb2180e6cf80932c9d62b7acf2fcd5da4184e4b682c69300c395543d0a5dd969;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdfea07f35c635c29f95cfbc1737a6b4970a2484340e94c443a1a34cb18801cc6775cc2fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16126ecd22eb9826b129b6479eed19031463d8fc21c0fff20af8b84d0343c8c09fcd049a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b90c00b6d7cca320f9bc54fbba9f5d35ee34c15b245e1bea6d79795d503d603f7a7a5bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18458b0502416fde88942740144236b31207d129e33c435fd6e2ff42e2942b11b3b36ee4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdb300a5c48e9313fd62b84db4da85c81d914ba0e6a936b33d3fe79468230caa85c0e5e65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h176be5e69b6647da98e1cee940b4934c1104eba0336517609d68ef14a0b9761f91197bdc4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166daddbff7af69a90d6fc46a858e2917e6954181cfa2ac7818945e888cda68860c0e37fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1947b22d7bae3354e56e94d254035e18ba680ba673f0dc5f799b6a2af3fa35c5f378979;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13ff2ff05c7db014173dfb15ab3dc2f0304871354a4223999c7d27b02f5df63ea6e965489;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d7cba2cd003fef12a85df135e9113505af9eea6fdd9d0b9ed7bfa9d1dd588897db01081;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1089a792b026bc8eebe4f88fde3106ca6da91df7a92371599dd677d54f0e2c573b21b4e49;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc061d53bc7263cf30d443008afa812ed289493d28468d840de0533cce82b28297daebc46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3bbdb4808a39c986abec6f22f4dfe360d63a36a661b6eb7991b18b52b10e58ec33d95444;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heec52891d15ec391d5508286a5974e40896abf60d7952310f0df013fea9cbe9d688825c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c443a0668597a19ff6e6798247060380b57b419f9d1078742d5d34751719dc9945a4acfe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ce5fb3102c06509bff8f93b09d28bb16082772e3167cb754f1feba9f400ecafd5eca180;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5980ecd9862438bd858238987f473197c631bc369ffe9124863a6b6549418f8288b3d275;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30a76af6fe7e1a16d52e6a00ba4c3091b77af1b33e797587c91a1340fdc2acaa3800794d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb797e6e7cd6f6b2af28b9a7567874e5e5713d61291ea22c97ce4f25af962f69c54ced801;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h280acb17288e15e9a435546a805631ac535b676826aa02660ac21080c25ef7118efa9eaa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h633cd303be58d3fc140e08d41c9f435e5e8dae5e565c1227b7fbcd9af608c50ff0b2e8c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habbb7a5aad77911ac012b1270b30ba736f68937371de25cd316f205e9d28defad9532335;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1587e3f78cf37159b8bf8b1215429699bb8b0aa72f3b0c41245325723e1167a7837c5fb7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19817172c48d8c8fc4a9725e09e7039387c8f06ab968c544303ee68dbdfcadda110d19241;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eef9784a560c3e456f88ae0a32d1153a4a30454319ce0ccb52a67f4e51160e8591c360ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1199bec6293a5171bba73dbf5963c934fe5bcea73fdc03cdb5f69e46ee23fa56afb33567f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heb6b7c418db1a9a27d186fbc8546e5368b22a9e3635bd4f637210ad41e17123825d9219e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0ece76a9b9efb28f6c1510e1f566a03fdb25d6601b3169de3096d1af7331d2ce5749359;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73a4d2ce72cb6e9662171131599b0388124dab1d875f8462cedc02b8aaa2c63ac1cf7245;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc79514620330dcdd925483cb0966957ce7d493db2a85f99bac225064c717ef83c6832853;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cb16f2d9cfbe1da60c0fd839274862a599eeaf1e9cf009622c923d30e673b2a31cf6a24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e84a47d53483ad0753d542d34e722181ae134c100c480b2208aebbb25b456a9122b43da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h67f51e4374816abdccf2b0168f43ccd94c2370aeac7353054c45810e51f5bd0160aa8a21;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87cee2925c72afc8c2079e6f7841be10ccfab8207143a0e9832e36ad098112749db2dbe6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9525d0d418c9f99234400a509d4882359ad6aa0ff60112fa394e3b567b56a2abbc82a9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa80a13ab2fcf786a5061220fea2bd50ac8d1583fc3ca993769c0a4ab34d4fc81513b1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1126391ddf920b458f6f7375ba1016e44ea099730821dee6446bbb4803c6425bda5ee7d9f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8b8daeea4012f0cca02f347f07be9c64864529900bea0ce2331690586609c0bf9b171b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1136f27e5a16a0e39746df8087a9d61fd19ef6d16ec1cd98fc0973762e1c6cf3086dae5fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5b97263e5df6404d6fe9fafe8e7053d1708e237ebb9addc66a70fe8c4f04cf347e4bab5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ea78da6667933f3e210df11ce70da76d391a32f9cd976c38faedacbe375c37fbe167043;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6f2b94574c7d614ef1a823caa97568e010d81cf92c5e37e2e686cff205417e0db1705d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd6f9d46b50d48261dc693a2ac2db9c216e3ab35300e55efcea82ebc35e4d0c9098b4d05;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179bd5683bed7f0fa84038355d6e485b39f26f3edb9cc9350b41cffd78cb5e7f1e6bda1e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1090d17009f5b2a8dcacf408dfa9468cd7251017617335ce2b34738bfd681421fa04979a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e21b4282283f933545d1ade6b5820196c5ba02a586f3ab91c81816772b98427aca74241;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66bac4be272cc735bc78d0cf912c25de7f92113dbad3ac2eaf0c4718615cc5a30a4637c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2074b36c31ae8cd0145a42b61c208402c1a82b172d5751f40f5dc8785455cdb20fcf0745;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1283cfca919671d710b732c0c37b8a4d070a03e77b8b0a2f1de49bdff303e713eeba08b6e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h157c56ff8cd7ee24148d5c2f1255caa18348d80ed3b6d5e326de68c0302427c049d3eb68f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he484e1b69c44f85ca3d650c9fe2f4690b908b542a14268a086755faa1cd39d57186e756;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfe3ea2be77e411d44d163a72b45fdefd4fa1aedefbcfe56284d60e82718021ddb20c757;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1221a7ccc2237fc9d8de9873912879e6ffeab709592376483831b7443fba23e09de8b8dd5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166f9da12747738fc6d680774d486c75617e665ea45fa2c81e8eedf52f5040edd34a31219;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb8e0491179628c0f0fb6d580d1e0d92d7725d4a6ce0917d24207ffa9ac86d83c1ac05fd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187b73222b878ee0aee7eeed7668a2809204885941da6dcee8cb553fc73e1047d274f5e9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ffeb03b469e6ac2048c82c613e42903928eb96153e5e02cc7466637ecfaf5df478d0285;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de3b2ed4a5d6ac8c2fe2c60545889bad59341e1f97c2a5409c88e83701db2c1ff43bd9a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133d389f9a79996d52e5f0572283d3b75985acdcc2f9baa6ddddae837ad1a12d8e4080387;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae487c3a31cc1889db57c140dda5b9944957cc0ca5db997e11b14262f62192c8747f0a86;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb42d46fbfb2ff9d697d5f340d03ec72ffdabac0c7a8c480f2fe407fe9da61afd9d7b3d6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117d63bec6f59870c8b8d8b3212e5ef58a933b2e1e296271debb378a1c398ae2eb2561198;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h104be9c84d0ad7e9929334a9a401e4f3ded01e3be8e2e2acdc99dbfdadbcdce5087266271;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9956c86d7abb9f027ddd0c197ecbb16a64db943dc7ffe8e19eccf5e2ad9e10c88a8f13a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1017a7fefa77b3b3a57d0a4aa7387a6eafb59af309be18dd7b7b0c5c998ff3ac6d64971ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62567cabf8a6d8cd15547660c7119558b1aa4592f64104d402be1b8eeec45aa2325476e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab4b7adf36971e83634097e8d32b8103e6b62e898c100cfd6672e53c26782885c446ba37;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1fab894049aa81f392e7e3edc851ae311a03b25cd1fd829fb87f213eaccc62cac8281f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h172d2811669feecb9ea30a8de86ba86c3066095e41d5624a8d486715244b2c623e5bea296;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7037436f4615795d400d0d6e790d6dd0847155d007dccc241e641cb74ac7c5099269774c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5235abfbb2d849295935c5fa4873a2c0065bb350ad6849355fa03f71944e362c5f5d453;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137a6349ad8c941efc9342d8a0bbfc296cc8452f30b3df367df3ef77b83fe32ec23697c50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0200d9791a6fcf4b2b14acf63361aaf92ecb67c124820dad7b475509281f6b1104f0618;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h142d7ded93c8211d07e9851e204205e7b8b4143c6587e4b9568926f0345a92553579e659e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6dd2ab920f94a7984486ea7e3ff6ee0eb518e833aade459a1d3f24a0b333365f7dbeeddb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h157c59106386e197fd12df7f5008ce572ffb5ed11e4e4690d0e6f4549b910957d6defb272;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1688bd9ec979689b41c3f95c080575fef79d877c9679ebd90b6286a375ee44e7099afc740;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed5cd61a81dc5af772b373705fc81d74f13ccce6026cb9339cf7ab8b0a7ddf21ed3bb1e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2f103686124162c03b08bea5450c0024b256715d9121a1fa0cf73a6037690637521f725;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1029018abe42be365cad98e51d0495de2a250deac3e9bc50e5f8bbcbd81279849df9c5f84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cf3d1cb662b763a3b8d09f57f18e87b99e69300fec1cb90ef9c153542d35685c6a801b76;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86a7f15d4e9abdaaf0ba229a837ac9a2fd3fc6a677a3bb98869ac8aa95e071a6e6e78243;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf93d146f8bbc6f161f355633adb7a5096c83573f21e18fedc86459fbc3ecc06ec1601595;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189add6be887fb13308f4681750dc2ea1115e24648ebda68bae81655dd4d434f2d5621469;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a580dae62f1df3f2b5bc8850364491f563eb83c1ac22faee8ddbbe2fd8ddc8c780b32dd2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3cb0e02e1c09af663e79ccd90987d4e517896db69daa34e7cb7374094f62c79b6c0cf1a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18337f2047ea19b2a964e1a8687dc529ecba88a6508b5d0351d22ede76e87bb102bf4654a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha8d2b999680dd94c847e87c5c9566b3078906e5f4ffa91847008436d0d4d86d912b035b0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12888d328fa8dbbafe54c5db3c34c94c9cedf934c35c2cb55a0e4be8c119760d05733530;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f0d353f1b2d1e6804ee3649202b810b1849182f8ae46fd94cc7739c8dff58e2f57838188;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c658d40aba94600e111bcdec2a59b10706ffc120e24a626bb80c1bda5b5159a11602ec63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13675f455fe21bb5f107d1401d1362c3647f7e158d42d72ed218fa4f3ef456ef0a705116a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1958b6460f9ffa75cf9cfeb10c70c2dbadc400e99d8894366f780612231734063754e7aa9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c72dd36a7ffc71342097275ac6fb80ab56d8bfcabc8ffe4627ec8a6a71e21b432ad5c28a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10865f5c88f867a0537bd5fc81428afe3190174c5897fc55089ad0fa0f7656019435a653e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h96de06772b19630bfedb306a8f7243e499e04ad142d11d270d706c8dc83fefdd2eef026f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62c6162de88497d111c6d8bf8d0b0b53d8b555b4a21efea89c28af73d23ffe6a8ff839e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1adbc0bc62c889029a6b12a8d66fcac2ad6dcd12f31e435de4d75e7fbc7a5d0fb6320cb56;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c78b48ffc4e0d89ac52f225aa5d7c558c07d0033109c96b07b1a55b840eca54fe496e048;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1751dc525abcadea5c0b2792bfea4624650d835820e30f36e28449e36f8f38393368f3b4c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ab77e2e03a1ba92eca8d9ccd0f46759a77aa13f6bdee27081e13a46474084b42d0536d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13197cd5e6a032b0596d611ccd631000584d18ca4f48c026830fe7400f8cd35ff9b17e6a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a19be61a8322f4499a4e715b7bc0ba41679082eb9aadf40f6f98625014307892ed43ed0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7da0a8acb0a3388889f9c23e2a5900edb52cd51ad2795da63f86bb31682724a0e3bd516e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ec70e085e9e990447c98b869e8650a68013f059867b4f7e16453ac4ea7862e4e1e1f70b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h997f47412ed32dbe4ce5f2a0e9d5db0b33f3d51e7f85c98d69fdef9396433c7a837f4b62;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0bfd62ccc819c1a02642ac52c729cfb83b72535338ea7403797c22acdd8583a5895983b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec80503374aebb606d9992fb27922a6fe4e310262e36a796498611aa2680776383478d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed78d93a6dd182b77431239956fd25b1e66ac27cc807f7155ec9328fafd2d91a5978f98b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1c47a019c8beb696ec0ee0e4c607b1065dcd017493b6f3906fd541db404f63a4f65140c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62afa1cbda16ff776b88075c9b49316923889ffb1f78b8d8fa62cf7da6ba6536ef022900;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4224aaf6bde2bfcdedca3b38f6d8c4e7f05e9d6081b05b49c8bf0d8e7fa5ae31bc1d739;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d746f2406e58098fdfa0408dcfde0b797de09a1e03b2b35f5f24e33b3d5e3d7dbf6342b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a64107f7094646c9c677460c36f62c497d9e310d78e45e74740aacd8ceb9162cfca7dc72;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h178d6d0daf1822a2f6410963d8ba1ed4d759303b9caa3c2f895ad38396030158f6ed369d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b4f667faeb08d93cdd7a8b04fedad5b966fe43bb8264de9db9d252f39d869c453658e098;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cac5c6d950044365f2b4ebcf4b276807670a130b91e4c2d53618d3773267f37998b9b9f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd55067f11128cfa6cf290c425fbb19552c2c3b30f44327f609211b1630303ac4b38caf50;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42bb4b2edefee1de11dfa96f7528506db8f64541c0f70217d572fa963d35e09b8fd809bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ac0b810a1d88a7e7e3da887a5f94b0de71fdfcb746746fc440eb044e481cd22450deb6b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc394c2e75db52e7b70b1e9ced38b22d942b5015aa2fda9dd5f95ef213f225213b4af2cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf2eb1811d1081cbc6a9b7d7dfa53129aff1220efedf2bc525211a20eaa7d1a80f3a3574;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha4213ef6b8ad91f4d4bd47e7793465ef92a9ec4cd892411dec7a9dd79934129bf84ea029;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b9f09e3553902ebfc462ec62ae2cd52d006b2bdf2ce5603e1fda3ac1858bef094c7e224a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179073d18f0e16934e0b9236031fdd1fc4a8d0f45f215f14839ee96b09b1dc10ae627ee7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8caf7849a6a2a3a125f4b75617cbe37da47d00f46f9afc5869a79086d473bb42904a1b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d8e99926bc16a6193613cdfaa6fecebc4e80dcf18e7d5bdf95893703c0a60ea6431015a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb23a848f1e24a47dba4690e8ae7aead4f176dda19882c868e6b7d870fdd68de58c4c072;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d8d9bde96561d59cf958cce098c2bf325e9b2e1105d9ab4c7d3c582a06fef27341f3d19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da23b2650216c4d8f915f7ceb04d4e7d3c0a0da83060f51bcb13f22f7d38074f080404eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87e0d3c630f0b26603248f8748df01a12dff80e3d7b7809e0e465a6d83e63b7dbc5c827e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7cc5d310ffa970d1c3b2cfff472c7f55344a8c380b2ebfffea1ce47cd431af5488a9562d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4e3fa49e9d7f9f927a2b3ff8c5688db5589e8e8527848f2dcb69916657ef5af16f6d1f4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d4dd5ff8d9984cf3ac327105e8c7b0f880c4500918d194c2c750f61df6e8377d3be965d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6ea00202939d9361f4cd5f3c8ac2892ae3631035b78163bb73412982000eeca2a343659;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d22cca97abad2bec70419c2bb3b43c6e05701eaa0b4ca7a6482268da9ffd4308da327760;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14f965284eb4503a34b056b53e18b103f05cf8e11f7bc0117091f5af377bd7e6e458b95f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17a800259b11d6ae4e11de00f81f2faf9c53f7601a4f5118fb6173416907819be8223ab89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbaafd3a1e6742e2d6aa3da05f85a1f554f0798bce329ee0c4c8730eda575be7aac8ffa22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60a43605df6b836ed2ff480fb509d8ddab3e3ef842db1f77e8168d4dac729770bcb5cc88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a12c98d933fd021c231de7bdae98f82bca93e74b46a085b4c530e317f1448fd222102a75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7e00ca745fc9a020b85bdd219c66445e30b0a0dfd4f9a72889f230fa4fe4333a28f6a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12dcf80814e76f2b9b72819b02f52728a33c23a38c20f4dcedb7ee944b4c8897cbc0bba9d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h70fc7310277e998d03f1b2fa45c306660c7b92f242ba354521571a536d7e105479e72cec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d34001f9866ffd2b4bfb81e01ef79b8b941cd55acdd8bcdd509b77114800797d0c1ac6ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb6f308e806bdc7508a82a7bb173907ee537827a8f670fb6210586c9b340339fa7c9b6ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b17bbf46909a5889a80249b06d76ac4d30c127f82a71da71c0859d9560760b31aded11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1764b3be644c24806de4651f495779906ede9f83a09f8cae2fd9700346237eff567648575;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae79bba0e5ae1437519e7c07dfd73fec4f9f3150386955d4387d8762cc804484a922a38e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h449fad0228809e49e2de1f78b4cf32cc6216606d5968d9e8146714480b18f9f60591c89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b5b61111fa6b9939ceefe2643438eb383bb074c9a161f6122bf54607ecf3e7e08aa501f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b7ee70831d7d49481a41badef3c1745c0ba98210861287a9bacc46facbe0502f32ee518;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd478011685264d4305e2acc457fe3738e5c937245d33c8c0f3ed9de6c441dfacf19f023c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1894396a7ba471f2333eabba1e71bded6b86b45d103c83785497d9ae21d33a47a17b8f7ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1908195c0499f64d46a8250e620ab31f1399f20f262f9ebe9657a167530015469f06d17ac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebb930d7cf5df33fa7efee2b71a2b79cc36f72196ae702850925273b6bcd4d1f0ea448d2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65a997bdd7199e7e473d8be113d8f83774be4deaac7e9662bce5ebf1babc056ae47f131f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162a95cf240034a2bc862922ba761f77e71a953b9140477ec7d67c072cfe54df1cbea8daa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b0a07b48fb1ba93bfc0052acab5402afe53f910731dd3e4f986d4d90c845f0da2655e02;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h79d9d57f682b8ca085d049db6cf161a052530f8f643db72bae5f61e8da71381f4ec8da15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfd11b2ed3b9fb83ff9c1ee0dd3f4b44d33dfbabeb8ab5f7d72eb4c4670f20542a33bbc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc9e3e38edb87d46b81234896b194d0f29ebfab76e65f61f6966a26cf08e0692a23a811a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7e4d69811d0fb2c796791e07aad6bd4d478d50cb4ec36300d06672d915e9bc10f43dd3e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f230ec6f63e98678b808abf2131523ddc94be312afad86e9e465d509cfe878ff6014e854;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he30c93ee55d1106ae5b5ca876869904332922a9ee9253684a4f8edad7b6eb344f7b3ed8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f371832947d39dad8cb215ecbfe41fae6bfdd9723f2ba3eb26dd9a8cd74266edc55ff7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h323db5306c56c0b25bf22de3cc72bcedace9c1e55414bee57bd3f99183c0e1c23371b2ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12592af0620d42c37cbd86dd83771207ca4d25f45147083c0391e3090885934da7e73ea0d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb67c53c9bc0c54fa4d8c8e17362e5d5f66ca0d22f8a3eb25ba9f999b920fa7a9cd8eb420;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12df6a2c80af8a28f4ad623a8cca66086559e462e5a8eb1f2fa98dfdbe527d408c5a2986b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h316ff68c84e65f1501940928d889096d17969e7cc329cf9cf8e62c16f78abf381ff2ee7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15feca0ecd8134fd888cc66cb6c1cc318b99bb61ebd0ccb22eb57730bd23ec41b8bffcf22;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbbac4851e1168e4c53b35b48f06e1c8c74822e4b4e2ce77381363f64539a06b6350ef08;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162842274f62cefc470c16def5662bf6d5eae91c0f466d5965eecec27118b1d45afbdfd69;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff21027dd0c54f6eeb3a6d2066673a10f8acf77d6499e7f4d66cacd9b754c0b0ca0dc914;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f36410f9c0d4c21436720efea4732b63fee535290b55e1b144893fd357ea5842366e20e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h33c5c0e899dce6d2d24ce5cca634faf90095061ca4d2a93360422c056c4566637485f4c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde54353c11cd2242464798d72ba49cf7a0f9cff1308c0abf7f970ff7e2ef590aa6de79b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17dbe26004ab10c0bbfd9282099ce19d75d3afdc069387969b5963d656a4346be458ed76b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ebb7067c651589eeeeb0b273f9224bb07bd4a79e20c055b4ba489ff99003665e66e35b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51637704b760b59531a0b30640bcfb87275d638544061ce9002ceeff1c1461a279bf0e54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3ebe7038610a69fe648e2c8504700a9df5558c3e3cb7495c3feffddaf3b6776c7aeb5c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8bfb089703c0a4ebbc8e679e60a70eb4a406c69a215f77ae03a4344105d72346c242aac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bad2e8e5a551b14eb31116793f4f359f788c15fb1c5f84460c6bbe816379c8261c45df80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h157b0712348f3774b5a3579afaa1b4f7242da1e002c3f07cacd2b348d0e6dfb91d629552b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6b3656ccf0de935ca99cfe4d0933217c62fc4fd52ff8435822a50f8b99eef56766a1455;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1365c6836623dc41c6e19a49212292c9be612c2c85ae2b10cc84c8b44cac60d297baac66f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1223f891effb778961ae52427af70f409d6d9a6b76e088489ba7129adb187b96e782577;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6aee99bfb19eac8a2cafb5b24fd3c8b8a242f084625dd07bebebb717a63a27749a25b23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aaace6249375c3e3965590a612bae6b74f1b3311886e7804ae0f7b3c25aacae975f185fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd926d8c7f15d85c7b22ef8d89603bb85f53442ec001fdaf0c1677c42959124bf7140258b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8c4eb038976b019bc04ca9cf0aa1c25027a6cf5edad21d92f0800994ee36c53a353ea8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a01a5f20af69ffbfac5fbe165960605f40ff1448a3022f1df61ab195422471341d2bb0a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a5cf3ba0e533b03bec8ae6c1bc1722966eb809ca9e600bc532aa7769f0a01181e53a5f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed61a09d4938c59a9c12fdf8ebe45f0fa4805bdcb0aeba497ffe42ef4a7eba29acbf670e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb216e4e011f11322fceeb9acb9133967a97f325c172d49b26d37f1b75d7d4006bcdb285c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e329ccbc2ce32cf1c3dae04ce2df17f24363e925359f026d9fbf0bc23012b9ab4b1d750c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1184f8c237325d4cfc3b12fbb40b37c828a5ca55d647948b4991edded8a80dc799c947148;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d93fa1e83fc9e257c5a2cef999aecc8720ac0bfbe986902a7bec5508e10705437e8dd4af;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13dda6a07c0504793fcdd83bdb52bf469ab1524b26422ca26258d7dd2bd16f519a22f7e92;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19cf8fb1142ac6f9738f92a089a2205e7245a14c2b0e2b520e82b4491ca0f622712325820;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69d851ebcdfd1a87bcbf47623eafa6cd91d35697f258cdf9a9122691a6f34fb8f0d3d40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4ab40f2d282376909d1a376109903781ae671bcb5d6190b6f66d018ff3131380a2052ff1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf167a8b5904891cc3580b94681913a251d8284ed18d70f82bcc93ffddb5852c12adb87d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6809b39ca8f2b3976df9a147bd2e60e7e49122754fa4105c974134121253234e9a18fbfc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135cc938013731f1525ecb27954ecbaaaa95878d3237ca99fe219ec9cdd9619b966adaa83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h40bcc6a62f3d43ddac632eb67e060014030ea28e84f872b974d21d463b0447c5dcfb4200;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6334721975e2da475d85d5eadec609be5ed154e64777cf89f2d24f4a0f684bf3a895b8f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117a0978ebb17d6607d23c30633d156d414d70dc3e9a2da73abc16c3d0e2aae8c8965fdcb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8483b941b4e606bb6edfea42cb3f26d5a9050cf4de39ff8a4cd827b30e7df2dbdca71f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h25ff88ba1ecf7686a02b897ae1f7224b3860afa6ad869cf8a8c9dd6845270123e55c6215;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb6b1877f5bbc78fd024ac1b4facd3e505b2a4eb89376b3904b6d64ace22565d1fa5b308;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fcffac84a5de5a06ad419e610d60d9909b1347ce68b54f99b914e8b0e7353c300c978d15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f15fd2c612ea22b6dc4b0ee577b0d47d5af02168c8024a6b8069ab8da5ea7b92b2ba1d5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hded91895d3f4e464155162110e386b7a5b4886ba2bf1c8d5597bce35f86ca7c2ab8240da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h839be76a4a85cb03d3ed1f1a6f99e86c3d7598c7a1186aa4af142e8877b3f3a3f8888126;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f072dcf09e87ea9b50e3efb86e73fb1f6c5c203512d5b6e607e2324fcaddd7904664a8e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f709b542e35879f584d5216fed04bdce79c90d850ec7f21fa431d7e8112a2efcf0b097b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dda58d5061304a433a3572541fcf6b0071c3b4e5ca506e03ab1bbf24579556fb94bb6a25;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1222332ceee8c7d71796ada10d5e269161fca0c008ad349d66e40a3cec6b50a5b8e736d51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c657630f309861670aab7778d8c0329ae5798dc90f47be6fcb61aa2142097358789c8b44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11560f6d4feaed185bf1d3239b9884e6c22e6c832067bc394d20e327eb0784ceb83cb31dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c20f09edf8f4f4a8e9b2564b93f7e49880c5cf694dc18aac9505692d3369246b97baadb;
        #1
        $finish();
    end
endmodule
