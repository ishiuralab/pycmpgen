module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [27:0] src29;
    reg [26:0] src30;
    reg [25:0] src31;
    reg [24:0] src32;
    reg [23:0] src33;
    reg [22:0] src34;
    reg [21:0] src35;
    reg [20:0] src36;
    reg [19:0] src37;
    reg [18:0] src38;
    reg [17:0] src39;
    reg [16:0] src40;
    reg [15:0] src41;
    reg [14:0] src42;
    reg [13:0] src43;
    reg [12:0] src44;
    reg [11:0] src45;
    reg [10:0] src46;
    reg [9:0] src47;
    reg [8:0] src48;
    reg [7:0] src49;
    reg [6:0] src50;
    reg [5:0] src51;
    reg [4:0] src52;
    reg [3:0] src53;
    reg [2:0] src54;
    reg [1:0] src55;
    reg [0:0] src56;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [57:0] srcsum;
    wire [57:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3])<<53) + ((src54[0] + src54[1] + src54[2])<<54) + ((src55[0] + src55[1])<<55) + ((src56[0])<<56);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdd7022e07813dbe7c7734583e604848a8a0d5f728ee1015255507d3f16725b15d0303560149a5fcaff11624d18e07612a1b6ba35abad6d6f16b6ddc5eecdf967deadfd0dd0a5053b4c7f645c624f9fda0343737567882c8bb661094107ba364890166292df459a8931;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6efc9902533b7d47cda1b8c02111dd5e98857828fd4c66754bac70ee1a93bb8671bd00b9b8c2a37714796a6b1adcc9ffe8b4afee0c32b15c59627f7338b007c9149a297ff9181d5a6718b7c7342b49cf7dee989ffb10acb721cde185f68b0763357b281f13818f0a34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eb09e28cb65029f5267604890f37606d25e20273e0dcd35edbeabcaa5b31fdf2eae53540166c753b4b5a177b2d8b77729bb3906ce26d8d2446fc010b99019873501dd22971733680f651e38e15b43d47f0fa5f83b7ce26b3a7145572d413966c5efbb5728d3c203c97;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d6b3966d3848a38ae5d63b3afb9b319d3f1d41aa0ffa0c5b4ac185af0508484f1d2c229bafdc9076c828fc45cdb649bbfb6fb00f5dbdbf26eaee1882f440d330d3d150bc576a58ffc5f1ac0c69190b631378956e4fca8f51d71fb3045025cb4668d378ed37684b132;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h896eea10a3111e44575a1f9a50e9e8a8b52dae42b5f17325c8d7612682ffc417d7feff5ca3daf14c2b339c0f754caf9bbafaa91ddc2efd51f2100af988d6709fef99af2a83547bfe9f993f7a626a99fe6bdc05bd01bd577a7efc97c79845739aba201a8a6b0f5656a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc6ae5e05fe7e20b07f575847e4cde4ac0ae28d45935df0aabc7ff6273f163677462d31e1129d101709062f4817765a88c64d67860c8f312169e1f383fac005c27a9b6fa76e3664abe1410ba6efc4aba5a2c2f95344093854d6ab2b944d83a33934e3ade3f31299cd1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1602b425f69178cd7264c83093bcbffe120291aacb519f8496c84fa6ca6e59c7de979ddb3f3521f1348c64e175aec1077beec6b197a253aacf34e1461e08fbf0e18d71992b9630bbeb278a690f754635be3325fea5cc150b2b5e23c4ed37648ed4e2d359344eec3cafa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3aea5e1a10a885d85dcfce81c3ee4a50499c798351806862bfc21b8b21f2cc6377718cc59660227c501d26a25916b51e49febd5368b659a699cdf151332630730f830ba1c960ffee067133aa74ad218c35771dcd0384ea2b433674719ba5be0993079a3158c24ed555;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h986f7d33afaecf17820ab0fd6fccb66b22df8a42a14fcb44cb6887d23a3819f3c353214f6b87fdc0896269af716b4683ccca2fc17b762d2b6f457bab440b02872e04331fe502db3a2fe33141533cb086ea81306f389b1885fe8cbbc883805792823d30a0e6c05cb73f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha52e024970f06b5aa1bd5858a9ebd2b725cfc815e9f1c4420a6ef17c2bb9a17359018c3fc739c151a0130da22e1d87406651eacf775e5670128306888bc0f954f6e9510bf9f303fb00bde8eada5760efccaf04efdca2d3aaf74587475947d3860f8ea59bbbee07ff37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9046ca42f0cfa8c8cda7a11bdd279096d2d10fda3d87ef4ed99e254b0d2870f91b74ca0ff51c5d246a8a7e45860b8118495f4310fcaa5bcd8de8026af3eef0caa6c9c47d8f1c523ec5d07731cb56f61afe9f3316aed557c83c0b603120187246606a503e14d79cacb7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eb3e429a4c2f62bec967ba8dabe6ff4ede45695acc798a578c7d7007f2a51ace8bcc6840c16268ce9c28799bba423eb52d08c2779dbc3c5e850dc5a0a062fde5f1ee974571cc86fcb1f24e3710ed031b55cf4a4095834529513d84417fde71197dc91ed2f1561047f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9db7444fd2755a401cf6053d79558b4d5c20a43a81f4f8deb995e20a46bacccaeb182ea28bc68b9c781fde88c7fbb689cbfa703cb6dd7ecf1b57c20f881f6cbbfeb24e9e27589f05ae776df623348baef506d57a7ac3e9971486f4ff3892ef5f6a5c8567f434a4b33;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce8d3e7c0188de91ac8d85886b337aaecd262e0edb5ddc8c06235193306e1c05c6b44c9db9538e2025407eb06c5c0d91c1d5b6890277697bd963c651d89e172158393bdfb7e9e391905338514a2298217f099824525a3427834e2be69cc17bdc767aa6ede12bfde422;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff2cd33fe3ed92fd9cb57c0e3d1d6f15f2c851e9c23551f978a3baa2b4d6949d38197038dda35add91efe2d787e4091977563973d48e897574b4aa029fde75e4a6c8174078a856acc42424adac826af63bd68ae53539458ca707720621cb059dc9b3e8662f4306d046;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96ba22882fa92fa341774558be5ded8646e7597bb9bb39350baad40604d5fb1d2bc3d0bb984e298e42bb0d04c633e3bc7a473f885febd85c58d192d69d5e60a5fc125d2a165e1858aa6d36e41ccde4a3d25e19f28b05e62b167262eea99d1396ea46876417cb5fcce8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10366766c610a8f63aece9cd03ca8d56077cc1503a8217f174d8819c99cd70a76150ea6d40d821925d25592217f1597c4c0d85ef73a7efa648405611b8d924423de7d1b9fa3a7f6de2985f99df5e0bbbf6777c8df37d884248dabd7166f5df4e0c07a30a2328518ae39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8bfe61fb22125a000032e98350fb976bdab1a319e0b2b5b6ef45d981bd17a5cae8ce39aade01cddcded6ab79c03caa0ce860c0d50d5dc070dc6cb8d0de3afe49049dee5cc8f6d547d6fcf9c8984c3db92dbf5f2eba09fb2f6d646ce1874e4cccfba920a29d6d24a013;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd817c541d598cd27ee8307e0ff76a7db968825b9a9b9bca5a40d239b55b9a1c38e7316b84b34365f0f72fdae88f958c9f5a876677ad6f421bca4e084fc950ea053bc05a3c18592ff063eed5e118e55ce1b5b4d4a311c4da1a9ea1d145f4b5a37c330d1556cbdc6e8cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d7bc5b915cc2be554bb26a3a2098d3cc589e06050cf2e4da9ec8829aa16c8970ad8248d145e1d6635636f012b82604fd46ed9b8f858812a250e4bb3a94a4339a114e1ffd0cccef3d6174d1b33fb30566db796d1398a1ddfc86c7d7f8c819260b928cc51b5506e27cc7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63a0d87c1a13d25900173a427a22adf21d8018f5cf95b6f26eb05129a91a1f476b7271a92636aa201099c6a0badb6564580493aa25bc74a220c34fdc381a47de0bda13aed1904b51cfde5de90e01d684a4f7a9b8f7ffdc0e84535580bb59725e6aebe1d300308d57ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hee4fb9fb50d4d228b58bd61ff66830c04908d9b6883118e01749f1e016848a61a1ff387f6ef101dfd3ade2f1d9bcf1dd17bc9203af8bc5f23184afe0706b7c802834dfbf74654cdfe44b9b8720a6056e0f0f03e9e2f159e1c32d8954ecbf047e5af9036c72672bd4af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5791f43586a3079d81f1250fb8e71290d73504e145c5420b31286c4aba8c376238722302f9eb96281e3184f01f2b1aa522e20218784178a91543501c25908df6a72eef6f79b1851ccae725ae0f1e9eec007d105dc61ac534f9736e96b37517cf3828da1c09952fe4d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1564bb6b4717fb82687a1bd314a5bb1f0b9a52be6a99440f41e49a0d1dd4fa3e591fff2f1986552a4916d86a2a0bb07c9a9da6cacbb5ad7cacfc2e2ce6ab0d4903fc66e7b92d1dbb4584d51fbb6eff71be4f816f598737a259997caaa67b76707d7709e884d1329e1c3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb02baf1ce81ae3318b28e54fb6de35b4d430aafc31c00e3fe54a804458dbf77cfcf27cfde1fcfce26ec480397a84312ed972d645df1c98e4aebb4c39eea051ddca98b1d148edf598c28ecdd8bed5c23a983a06c9ac6258eaf90a39078bf48b9d62eff1c32a7f4ba160;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb12fbdd31201594f2a07286451c45793458646d8cdc649dbe55f5ba260d10e2e7cec543ba9f2eed01ad7798f14ea72ace877d0fe39df960a44a5e742adcc80b63ca6378e7fda5c99bccfa63e137eb0895ac4d0421d28f1c1492347839e4dfc60ae26db73996feab6c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19dafe6fdb964875127c67a154ea9824596b851e15538727f75cf55f045241c8e077e29ba0437179aa23a831da33d6fc7efd2379eb8d4d885bb12626dc4e39e84f620254f520eb4197dc5a3e640ac625916d71638e0e64dafdc0bd2766d803e50f3599f4a2444e1fb19;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa01ebbe597271e12c5baddeb51b51c339295912227887f5c8f4fc7eb04c830f81443e0211b611883f714365c0fe0c2f294fc28e9e2274ce8aee422e1745c0ba2ade4874fa104b6fcd51cde5ae7ac2804ae9d38d779512ef8bc9814b85da9d039404bf5568e8ce5fe7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c600a3a2b48f782f49019257dac999c715b95e96cab17a6eaa18dfb436effe51a74fae4452168d0aeadaf2f2045c728ed6a20a3122c4cb7281aa0e8613d1797dde4debe47b8fa0e9bbbe40312a041d8046ce44836a945ee24278760e448d6b12e6f7c99f4f5a3cbca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b822913cd79fd797e96f3389b98f2afb64a1882e33d87683ffe3c38f0c056fa1b1dfdc8a85242b724b36190cd68e3c78315b4c8f5c9b81569d028ec884e01d68ce1033e38e02b11db984ae6e286bb76e1e0ccaeeb683913aef814f86cb9fd0e3f900cfc1df1368a7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h181ec111e2f071eb064e4d82c6bcf619ae8a5b87c311fb6cfc5d57989000860fcb18861a4cdeb75d1a0e22224fd37b0533509ca802576b4476682f13cfd24ec5e286b77ef73770bfa6d6d7b733e765a349c2a590c89bcf2d6271001b5c8adc94d0e436330369f22e37e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93067c606b62d54e45b16ee5afade5756c4cf7337e85a38905bee0b5065f4a3aff5eafdf926a2ac47b3fa530ac1e73b306376a3d426c092577c6baf28a1d064d7ec378e083ff33e93b0a189998127befbbc8081a9eecd83b8aeb8db631f16b347b5d6d28514573f860;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a71e360899d6b1716710e97d6a7d4675014c98db3dbe2f51ed825ebc66b1051eeb3063234aad4dd1b97dc19685f95ca41930cb244d90d45690890bb77d590586321a2550574096d0d301f39f8d34916d23cbf510dc6793acd1061a6feca68676662e8e9cabcc5f465;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h403c06946015b5b7738a9ada26cb5ddeafdb7d9c95a276c5a0858475b646546c488770be200a4f2a7e22d0089abe506770854f5d1774b320c91fb541ba87b669ddaa7383f72e4192fad517dedf5fa76a26e92fc70e5e5c804d224c5e5a69e856b6ed31780840bb4fd6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144824294ceb62ed152deb4284357fb55c500bc759983a6b3edf5c2eda9738475099000f58adebf4e1dc55469f64472c3e7d3cd313fb02f2db89b69e4baa3483e3e89095a0e0fb2e150146d39289b14c0fa629d3a6e03d33c1e8c47eb1a97694f7aa7d2dcaeb0b2cf66;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h46f0601586398a1a72413d685004748ffb35ab62e243a99a05ba986d4e4c7184b2228208e1bc5e78436a5cac812740d960145723a5961dadfbfff5644a88b447979c9661b275893a98b3e4736c3fe62d44eee6ba965af4399707bad75e62297849c5f6cda5864b90da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fb81cd5cb6222c47492901527b529d4ed4536f98294847bcc0adb14b7f8f26cf956470b99ce1071b527d5fafc4d933dcd25ce3d21dd91bc5cec0ce273090c2fbce2547d0103dbab996cd260a71214aabe22a7a7e3db1eb11d93f7c8b2366bab1da40bd1296450a550;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ab64d63c4f5285580637fe9d23edb6e387a078e7a9a13ef487142a87bacebf2178553b09e33ce61e1e45f025346f2bcec3190315bb89c4a2705eee3cad01fb1675c5200c20c47d134851c5240111c77451e3c086cb53e585ae4be0c1c3e1e18ae1cc14c7ebe0ab638;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b7d51e1586d5073a39dc1d78c67c50b59e9af0014d79e0bb53c5844b305fadde447f6fadab0dee9884a8906bd02b5796ff143e8822b8d6ce6ec765ea324d2e2477d1a0a74ae65f2f0228b984be1a5dcd88629a77996072fd1d1bccec17f41ec6b051fb437871e21fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e00e2517fbf50831e0e9702bb0af2629135d7eb257e762d1df77195d082d00690289a9767cfde72d88306d3f0d94032f3d69ef8091131b32e692a3559ed92152b344af8030ac2258ecc12101ac056a6b9fc586c0fab5be68e598a88a60ba20ea07f34de4f28b31487;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc68b4c69c2add87324e14f10d3872106f85ddbceab8268080ecb26588390b98e7a2d8291fed407de7756ec1e1ca3f03907d3e3b1d59b02dd3a2992c0f7e9fa54961e03ef278238b6f2eab0b674078c4e72cae110dc33c173bd92fff4fb6f4c6e60bddec0de9d75758;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b73fd6944a0fbd696a46309d1dfb1b6734a2b0ab14c74579af7f9745af45ba57704c09981bbea713ec995f97fbcd0e652481c30ba110e7461764102ebd537f082054882993fa72404285d0e3a2992d9b9a0607f9c5d8c14072735c0de2e2585e85c81b30b812971f40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101dfdd7c2dae7b98f253b0c8752462d5da7a0de02f25322356f9b9bf2d2140bd39722150c82c241f10aa41b13b8975f4a8f1c3f6c035a1273193d56dc1b7f24a0ead9a933b29bcf19a4036aa2e97467dd9ab73d703ae1d247afc571316d3214ebf1373464a4c4b8d4d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h106918f7c80b0060b93abed583ceb29db4ea625386da257b62a1df2c7f54c9ebd0f3ce0454a46cc8a91296769236ce7970665a25682d6ee0968f5e75aee6c31d8c0d75df25dd15698c1ddfdd2fc6e856a9bed571bcfd2359feb939a528c800f7c1b4a06a462ec487142;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190b0bf410d2e93c2d413badedccec2f45d5ca1d3aa8293ca73bfa60cbcdb91a079a751b1d686a9713035a9df9c195b9e3545684e462fc69114219943139795f2358a9ab3e67b3cb5151cd5aa36fa6f2f2728c645d4be2e289f19169a085b71d5c75e3266a8702db1a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13fafa19c0035f035b358c6092d0157a8ff3a8ae2f5ca02d93eacd495431c4b16b74152b1392c5c85aea6b8bc6127669e19f3562304f581a50aa575f663c2af32b7c23732aba2e73b9d32e8b7db8e743be1579cb2c44fcae7f377793d9f57814663cbca4cb41ec6c40d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3da0fa9de14db2e1e83a54cd0323d52aa4d530c06606b51fa63c21725e26285f921f73e0fbc4188138cdbd0f9a4b924cf56cea44e14280f0e8245eb6efec03c39c2c7dcf153f00e53af1e49edfe72153860c1723f471627f5fc8b3929b7255040daf36a86cc18f7ea1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170210e7401b5e7c8dd803bead54c957a1d1f23dffc9d5105f536d3661aafaad5547a221b05efb994ca8ec8e9cfb3ae4f0f00c15a90fcc40757e19d1e06d354d44de0f9c88402cea8784e024a39a05d81463f074d3e958817d1efa55fbe50d43b93e62c48f3113a2780;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b65553bf408b1f7ce9630e99d75cd8500b2f73877d927c2c8480f9aba6e89d173e031aa0084fdd1adbdace119a2b0e3f7e85d8f3f2653f607b86b5ecc96786187199190419b052d2797bc9ead03e7ceb0436379b33ba8a5849b45614d18cf2a22a66f2d40ceaf1aef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe3d00f2babe5a08d43e8275cbd96b98e26850b0da35b4f0e5d3f8c2afdab8f10ccb1eccb0d8dd05ed80dd02b0d9a6e0ce1d088e409de7c6bb078e1aab493302a5529bd5bd7a6326e3464a1914da36ea8be791572dc83eb6d2285648447c235b36f8a2b781cd9f5635;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ddec789eb61cd6f505f144b24f84871847bcf0753a8a2cc0b0f8f47910ad5858d917f97e93bd5123b9c29d1d02af52cc3112063835491fcb937ed2960c74be7eb5253ef8fdd581a2e662184dd5a0c73c7953ed79cd14b28885bce14b699c9aa63f8a10bd885451410;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe799643120c12c95b87f1116458b68454d9ca5d633c95139deeff73909bb6dbad93af2775bb1d350fc43d028db8b9aca533e780bdf0f386306fae585b19727dfa5e55fa62af0d61654d03682f7e529fd85e89ce0e5eaa959bdd92ce35ab16153b5f99a4291b41199a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h57e9ef3afaa33de767af5a4b29cb80546158217cf8713f38e6e4d58bdd2b281ec9ac4282ba504d748aa88d1f8a83447d4edead33b4af92c61d573b1123b76775d36c1a22cf6e9c8d367c95fd7cda658f9c501ab55efffbc2e036c15773d0eea35da1cfb2b85d93a826;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14eaeb8a09d98e4e51eb45df954d36fb6c3d69b7b1b5384e91dfd99be84fad7df021870b23181d8fc0e2e892de25c518f642fdb90706e5b74de72d5526269fb7ae3c2c08b0d1450aa9f1b28d208476ef3da903b7fbcbfd4e581def484a1de2b8dd9d58bb8389470abba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hebc6d77fd366eee6fc8a6d0d8b3ec01e3d0e4051ae901a08587962258d29228c35245d62d54b8b5278e4a2faca3c1f8b077f3fec93828e016410705ebda7ccc00ce66b64fd24acdc15397ab9f9918b7f6615837ef3e9a1af123a2cf00c801ddb0648edbecce8eace8c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7667b6b2a0f80af38b4d53d62d556acc8d28cdaf97c3e17bbe29450b93d746384690c6c043ba827effd005efa981cf688b07b26690dd24fb4f9471c30bf4cfc9ecc6874a325a14e6901c70b5a6e1d79fa4650e003f080d502db4bb3b658430ed8a96857901f7b42112;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a97a8fc2ed12506da9de7aee67ae17d281d7c9b77fadc2d4bc565df6e063da650d627f6bdf48aaf50f5817edc9997a7edec7bcb46293d83087a4d61404248537c97d3c37831cd1c7704ebbf93234845454558ff5f06f8091411fba0a8c5afc6f04f9050f50bcd90ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e66a13e4312d235d91a3da929004fbc61bd278a6a9cfb1de4b971137688292d51e7b2f627fe2b0f67de08027af8ecd0b265e13521930f0ae48330ffc71c8a54afe488c2d59b0fd392ec9dbbf760a7f303ee1d633727e587963e5493b0710fca69208d0b9ed611e5b83;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h934266665771ef48d59868c2d19b40f0c7f51e4680b432c7e5a558341f20da0100a411a48793f88b1ec6ec6b82f65fe7951ff5cb006135ae17d8b81a786aa1bc747b32e5a14e110bf757729fd160229bbbb50d4339e45d956a974bc78f8b89552c7fd581ff04c611ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb68325184decd8527cf4f51843df4f68305de2e0dc2c03c873eb6ab8b8c6b8201eb4c76d424eb500f8adc26722f28e92fc27ae6c550be04c71899a68e4d57d94b56b39d28b65803137e38b83292ff094a1eff5e13f0935cc46fecd4fe3ad8d6dacec367a61a2ea3480;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha44473da1ad995efa12597c3c9b78b4a6e024d01c641c0e22766dd204591cbd1c7cd5d65e7f973ebb5d3fd67fdd9ce9359f062699cee42fc8fad17318eb4d3526792a2dbea5037630e0f37ffd8ab68504f5628c529f02b627f8f861989631278c6d5a1955daecac429;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16309829b9541a7f4f663488dacf1c1ba269673fef1e22cecd5d782775c29a473d7bddae0410ee95b0b0f63bce34c10d338f05a154c6c41fc127bafdbfcb786bc0ff307b62f582b5e4c86c39eee05e27a1ef85f3732d2b10f49e61590e223746a25b391b3cf0b3bc8c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he16332e432db9dc728455d501a7f70a52bd354f1f404f9388b6cf6fa1f9b2a6dcbed00d0b0af8853e38e167ce26c848de782f1e18f6e89c0995c31c569ab06aeed59d958df8654bb02905a916bec3d68800eef12c048375d70fa670a0acb9030d3712d36229d9f5603;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c0bf0ab9d30fc47cadf971e52be633de290ef84cf79830563fd484f0b2b8c246932bf6b2884106cc2e1a12b9ac16f3a5874da3ee9aae796e126590abc75a73bc02dd3a8d02f82cce182d1723f78e98ac6ccba4ba5dea89d7d75a5cdf5701c0fbfca293570ce6f1b94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he6b5230011c4353a9bfa6fb8f96cccd8cc38a7c8b20ed0304f52d55e160498223411b8471f7b6b2c7014261697344bcfa103f1f687c1786cb9a50ed476dbc567ccb4709d4d694e10f19f3e3b825c5397feb9131709abac07a080db613a2fd1b90246ab4b3e9deeb953;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h381d113cdfe63bc29249bd72ec10f3a2031b3ac8b07c4e84acd257768915c6fc0761e5116e7196b23bc4600f6743a4a2acb66f9d68d6a719c94731326e8f2808d0db8a448a22fc4c6289f8e9b1203fcd01c5f4066deb0a963bcb8034df99e45bbd7f1705a0823e262a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0455b848d6c06dae5e673f813f1787dfe00bde6652a0b4c675c35ee257a0fd5fd9861b614e64def1a6eaa06efff8e6a209df1f8ae00314375e904311241c2c55fefeb7424928115e52a7ad7398d293855a4080951a67702c76454129a91df8b37bbd72726cf7ed5f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1816365d6cb5051712b3dd0024b12fbe6f9c09def857921df0b3a07bdc771c93a8deb09d71f8b63c8075ac2f7606d0e4f478e97f53d6047ae5ac91fa53eeed34eb123dfabe8a01a06169c930779dc92e43287deb02b20ca4c287d1626c2632beafa94901c19b84745a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd7c749b64534fae9927c7a9f0333401fd487d7c99df96616af235f89cf2a3e83377da5593ba5eaf2d6b8b8d7f10d61c2216ac8e08dbe2dbdfde437e3ed13b36ea423c8a94b1bcba933c5d90bd46e3d462588f998e763ed00e55ea43f1e2533d112ea3d1d8deda957e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17075e72791f5949c3eb563665f3522e3674cf5e00c19692f2cdb0c0f43deeae9498fc4e3574c5cdf08d5a5cd067254e72b006665f28ddb5d433481dc3cd92ba51d5076e2e177c3f89367f2ee69890d1499da17584cb94e45e942fa16c6e3e33049f45ad3e6a1b678a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a125aa6ae79894be16f8ad087c7a25dd682661b98560183053562dc7f9d5b52ac13e243381b3e439d681c165c67e1aeeb9b36680107851d4ff66517f33b0a67477cefd80bc471dd7782474362f4355781629522395f5951b018997e21dda34237111fb44c238a19881;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19dfab21f4949850f65638624f62eed04b439774153c82baff722bc474eb5313db3436002b887064b5de1ca35a25ddce95ead9c30b6a5232291dd5a70da73873cc9c0e20fb8a0b4090fc3b0eaafa4a4f520fc40c37a974150a4eb9d84b1cb9420178a62b39756a95f5b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c848d235cfb51dc07e757da775963e6b66e3344e51369cfeafb2ae5a48bf285b0e4763c6c23ae2e6a0041b6585d043102879a43cea9b919ace3be4ae3dd1e053b38a33343c2b69a9feafda22798690e1ce2c3bb68c736b5c6e4603c9e92104a3cecd34e0c04cba0e45;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8b58770b3c73c1aaaf18b45528d76eaefbb478e629094f38aec6487ee77f92c04229589ab0b5d36c565aa3d7e61f05910793c19edea4d8c5d2504dbdfe725ccf0d02b042d30bb794a1b0e93b6ed72402eb0664360634bf8250cd808f1d8293ea5c53a2bbcf50d2cb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba91c063a57e149d5aeedfb5821b0a0b79fbb76916572ceef9e4cb693ebb08baacb4186ea241981c501d00bd559c1ff82e6747d170e3ae374a1af8ae7f2a6e8a2f313acc75a64ca63cfadf2d1df23bf2984ea3ca3ab2138173c885b2b82a1c15585c7671650598c60c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1efc571bda583fa8f4b43b0b28bec5eefb24d19858b85249c83b64a2a2db42905b3a357f725851ca309986de84afc7f98447108f23746041182b97dc2cba40bdb3c4c19671a74a402b10dfb7cffcba18eff87bd759d37884e3bd6c05a72e104eafeb6f85dbc3eff3812;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5dae22fa594fba485a11f1df794eb567fc14258db4044dc1f0520d6073254eeebca5dd824236281d8a51acb28befbe4fee1dab6ab56103c377ac75686f9bdd551eb126c9ba34d6e3548c77bf523e9597b9a8a0d2dfc4f63468c26548a34d64b9c1a02b4808a240f76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d641bcd200cd250b98340e997e41e0f702815b06e1232e29bd7026f5e4ce05b8ed7a7815794a6ad89e70990926318f224860fc2c107a068436d4c0ac72c1507eae32e4dfb2fc3e18b563989352934424d61d7b7971c91264dc9e4118f61177af7e7e646a7e96cd6793;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf21fc6f41a7b82568d915e89c4f3055dad3e1cdd7a872f25965dff7864859314fac2c9c150f57b9318d6fab8b5b9fd262713beda9c94849da1a94866a6df0ca75cca6a105270d5287194ccc8faeb5b5c279583277c3045d972f51408a7bb1c030f2352e5d8927ba660;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72ba5275740034d77be1c6eed440fc0aaca42982435308465b0e7fd9f5e0b3d4138ab1bf3c329d4e1d7f28880182086a9b6f2665e2295ec48c787196a7fb4813273a4b89ff9fe34277adeb6d1d4f1bba5fe70a3093d8fbea0c258cda542def2fc59bfc2f00ea6b345e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h50408c42a429108f397aa1de1847f1ed76c3d8294ba2b66107f54165b9693424df2fe2c95eee923cc79f735fbfef585b34752f1ab9f7f8115a104e3f4effd44c11d9d0f1d84ed198d545cce202db89592476349d48ff7b2e778afcabac0d501a2e5c0ba284dd8c6443;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10882849fafed46fd5c8436eb1b677bebdb50029ee3937d1ff6c2cb6a1bd16e63d27927302a08b55383f5662f2c4ba56ddf6a022d409b0a97957fa93533ea0da7aaa397830f27394e34ab77791a8cab36a29a58f45cfb6904b0854ff6c5df7f45b121293ef64d6d9d51;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7e5a7a954ef60cf14b80233e66ea7c7c33fbac937b3faa403d7326491f0fe5724cca937c5be657ab4b442618dbc9afba5a3d3e162678cb7c63fdff9989e52a10769a173528a478f214c6d1b453bcd8e723fbdef2e2d6d324da1778ecc97c13e12813cb8369094e641;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb34d062922bda55ce5a6e2f16831b206d0413f116dec3b161e5d352746b3112b0705f31a1e5a259318361905cc8d2bd228215ad70c90556babe91d1b727eebff4f44f26402406d2a1643adcc1fa91f09efd2c8f8dc4c334f637197031e5c4a78e2bd6e26925775c5e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb04fc7c4546db76f4e4739a12eab889d68ae506a63cce5005502b970a6a46fb7cc21589485cd78a10aaa5b3506f56d53f5dc4ab695a139ae446122c436d4b258f4b2fd8c92801d7218dc8fd493c11baf91a85d3aae94f43895a42772628923ec55e27f8df6fdee95f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hef26324229b60930cc96d39044aea48b485d16e3a74848c3450db4461ec65112854925e427e57380032581dfb5e5ab0bb50e33ff28a7709dd86998dfedf46da851c5e117ffaa91badefbc182c61f4941e635db7eeada56eba6342b9560b5cb0165b264a28b66a58076;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc4e49245c61f0e33e26c88d40da68da43519b8f96c94d47bb29e23759d91b9e66dd97581642f105b43f83363b89beda30bfa3b40972c0010a20931a5a689d472581cca8c1a6fc24a757ff02c1cffd34c914545eb399c5cf4d3f646ae3ac0babb1ef620fae1ff16f439;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1643143b36ea0a9220b585b8ede6d79cf5751ec4714971403df6e9bc7478ddc66dd93a5c4ab82e0707b61300c9bfe9c3c07bea418cfb47b566f37b06d8821901e597abfd3a68ca088761c05e15285d3859a8387f0feed34e7aa65628670e7c256c24ef4c51e13f27aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h171e20502db92841de54192b4ba82c810aeafd0501b8deb18445b436a3f6839b2023ad4d48579c67ac8cee856111da2007806f13c451da8c712bba74f76a0d7087fe190ff6a72e455530e00322ee5b7c0c487b31b1a3ea9c29b0510284cae8d2b023665210b63c65099;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6dbf84b818b5a0bac77b137158b8acebe6747a4b371d61a676b8eeffcf96a6d0eadcc3b75940bd7a6b49659264a61ec66c75ae58688be3a81edd93ddfcea2d2874df4e5ad2af874cde9b9f17195fee256b2c7348c622f4bf0e74a66fdc40b9cfc0f68f087ce75b0d37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h84cb134ce659ecb73c848bed3f6642b798062b6671f3ab2ae95a5e06d727ed2a3c3f51fa68a386f0965d8a68fa28830197d275fb6aaa6022ea9dd9f2e2bd9d1f1d7aaef8bafe9a4e42369bb2618f064cce44843f3108d6e36dfcba340415a0a44053f9292caabc8e54;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b8f950f0589996276a0262a54995f3269f0f17265f27bd58c0934edd95b33d6584ad0893be26ed5af3ec9b98c3cabb7ab14e8bf59a50f8c6c89c52886d34b4fee653cedcb20db30549fb190d8eb46c6ee701b64e9ba2aca7346a99e503da436495d3e0465fccd908b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b54b25955d1312e55773f1a15cf4ffb6a0deee403646ade0abd2d844ba949368ec417606d420fa9b20f8eb01576c7353a12ae21ce1f2c6e027c00eba2c7df24822416085496388f076ab6d81f2242617aedf8f55642d1956bf35b1a42c198136032bb34343adccca4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172e1d2fdef38ed731c23d99cc5f231457f01c51a9ab077bd5eeb30d40f30d6a18ade307b3a65c1ec6f3e9d51cee3641cb70ec8675379f1e3f21d69fb8002911e1c4472ee1357ef95029820d04264744636c0c072ab86872b688b249c1206fb8b74620a13a45cfc9d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3b7d19f26f9eddbc054fc5dbfb3946de7d700b09e0700780308ade43054a43099c499fcf5a2a9350e4787627910f7d517bbe87a3e2059825045d7f468424e1fad388ef05d0a110ad54ad8177f3b14796be78741245ba98e6c62996f1fe1b44cffc0619da5840669b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14384825bebb4f73ef7227c3f150acdcb174f27038a6deff8bc33b7f18e6c629258a295e65d4fe97f1b20e1a106b95c0cea4ffacaf3a222f33408a2ff804f5702ad1d74aca8b2f500b0d95c72a92e31e29b0e787a3095ee3e7d12e3082bfb4aeeecf1e3b12b6d78b4a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14fdce3b1ae9a13c12d2f3fcbac38d5dc6027c854041b4633e145a9b5bf288d336ca4d707d6f0e1b2193685d7d47f600be474ac9490408e15829d8721cc5ccb3eff12554016a70892f09a0c36a8467e43a52367ad8dbe75100209f3872c85ffe5e897e2f90fba4fe992;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h29bd0258923fba131ab185319f8b96da93474795dfe5b232da3ef2e55af201456f61c191f4c2b7c4c7513b5b9a559fec9572204a1fb8a8ccfb14000a73dfda4105cc92c4e680a0b0a9a7755c502a79de119e744bcf92a2133ee5e74c1c03871a5c833f297cd2db402b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179ff731336a8e3507ead1b1ab250bbc7056a5c52ecb95f912a607383cdcca55e54b18706ac6892dd7236758dd7719175a6b61d83857500914593b7868e032d9bed2c11d82666853ce87364b16d44bb48ce76744c9f7a64bb8bb602052686a81ce4b4c1b6e0a8948e5a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h189ca453df8703715ae470af188cccfd01d228f64438269db2c40498bf4c3050fb77edd92faeb4e4d5d6d5787038dcc30b1a420144a852f06463768f19434d5695bbdd0fab696d7a7d28e8b5e7ea6562763939783d9b41f133584097174b19e8089ec2f143e9b08fd74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h345a8f653ae6c4d2370ba69ba2c835d6c2978cd03d848637f933397715442fe7abddd5f8c19669f65dc21c47c3c207197e231f2bfeacfe57fe3b584c2385e7ddf7c2278e80c89ae42a8846fe10ce27944830bc8f30e6a2797d71e4af0bb371f43b2bd4ebe4fafe771e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17722bfb3a3805abdb20cb58c7cdcf9d90326d787692e350787d754e8e83fb6d332f43c89b13a3ea5f18de41163c6bf30b366e7f5bb99ba2901d726123fdbc64411faa7794d5bf137401c58cf850b3738eb3aa9ae9eafa5b6287758381fbd9b01f00087a17fa07f7948;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1daff496d68e8e5419b7e2a0ee3c0e107a728d670ca0db4a9c490de2947fa884c932238365018a04c609b63be82827a9332dbaaf8d9cc6cd3ff104b4509b1359b56b4621741fa5e383a85a43fd2b7d74d6105c4d5b88c5fa8b1376849785337abfc0d77a1c53d08977b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14469d54bd073d1886fd495878358aa1ad437b34d25c7a52fd5f45dee208c71021ca7438b9ac9ccc511d166524a08d3baee42655203cf7d12f4f09e614140af975ed379f7bf85666c48db683e8819a5a7d121ea4c7f3433fe209d6149c3de58ffd01be1fb0dec4d1038;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193a5e5d7f7b03e1ef1437b9fbfcdc546a5e02b2f8d8e7ed95f17f7d7367e5475b74860be8a1ca4f6f6f195c396ec2441cafed285068ab96fd805e25fb4b7c00c28064bbd693191a7a16fa948c8a978f9ff7684776f60f2bf39f056a1ea05cb2d54cd61edd48099f371;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee407d612779c61074de6745fda7fdb3914910b6ff4753df63a80d25205953572fd03f568c5bebdc98f8d676ac5a63c77aa9e359ff2f5e34fc31c8863c68df1a70e01cc66c767bd2e63a4f6110c9a0a4aae5f6d0c14a362b410b03991c7907fee72550381866ec051d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ad379eab5eab813e69ff246d784921c6c51ba8216c11c1aea39fdc82e4194a2b4db60768923dc3e9347e0684cc8e2f694d6ada635f25849c90d33169b002cd52d5499dcfef1a89e8414d331ba2f8e1c85c80a5f7e2ee27b2045dec0f60b3b41f732d069f05b7c272b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7df5f4b3b9e7d4fd7df974cfa76d75f96d2c712c2b6e24426b27e40626997aa1abc4e0dea1898b963e4c45b6b1d5ebbc735afe2607f750050f31b06d8481a4a6340c3f9944929a5f8fb1f30044b4f46713edeace080eb9726528dd23dae0ba197537ed602228adb59b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce5789858690e18fa02efb3503593152698e25e3137264ea33bf4cfc6163b71f408f6cded7d2ff670a98355c57d988e8dd1472a389166de129f82ca906f6fd54ea6de8b8155daca4314d0f3a32faa9a2ffa7b69aba77de8f9426c02f421d1ea5caa9a7550775df659f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h35d38fc8392ec5c691d4d8f0c4d760a66dfe0755160876cbf8d7bf1b6711211efc62ea932d12a9624350eb39c869894602c412b9e35a3da7d5890f6c30ce7f74eeb86bc42baf5da672dcd3b4561a11a9c0b8195acd47b02ae812c31f5b149628ce29fc123f5e5df3ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eaa4bfb927794f92cd7676c978f3b7560965ffdec8ce9cbfb912c95713eac5cd71add67574c308b74936c27362fd19e044f6febaa9fc76495fb105e03abdf2a9505189c497c4eb2439275e1d723dfb674fca8a33e6b07c3e09704eb6942ac1edb4cc2ac329dd111c1a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c55ba537e5373bdacc42dbf3b7e005411fc00bd50576ab3b2d28e87837e26b269369ba0965ab4f50300701c945ec16796b248a1a5368d6373fb461472c680e98ba03b76021dd040d89aed047373b1bb3de9dae92a94fcfd6fd002183dc33f674983cd91e205a054fe6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123962b3227d612e1e6bac09c90b213825ba69cb7397d4a5f99e615ad76882e49cb1cd94de327e0a6c157e09acb55ed3e4d4cefb952dfc50b5dacd4c688ad9cb71152d07f2a7a19d80740ab4f5ebfadc92c5c3394cb5c3aeb94383d86248da3a8fe60353b3136353c1e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168b304b49ffca1b9ba3a65b9b7fa9d2f7799df61e6abadd05ef0cbd24ee367feec8a394617ebb899fec89662ee90eeff5a1dc5ac58806aabcc8b2abbb4c14ed6899d02e3dfc56bd1431590a852d7708199a091f3547f6dfa2cb492158f27f2485a2a77c4524762fc9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h691b287f41e11f5c55d9a0722f7b1e93e94271697293f7728de7f54ccfbe262fc5a76e4032ed2c76fefd269831f7fbfdcf694337b1a88d05130ad141ed1af1458a2f67fd18d5a16889487fe1df254527d1573facb85c1de0843a5994651bea7c7e49696aaec3fac0f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3ea8b0b434316f5aca905f3f0f1599bbe1c914586dd5b6da7728d5b1ee85f0858ed82b6e450e4c7921fce58e15fe0763104856f161f98f787a1b878987d817f2010cef916a05599b51b65772aea6456c11f30a58ffde4371c17f32463f12e85bb74cae5bfdf84c8d43;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha419eeeeaa88ce7226994332baed269fce30776bc413b8520e79987ec4526a97202573d43139525840b549e5d0d762208b28efcc2a35f1f510981645d3223f40cada21f695ef0818193cfae8d828c541ed53efe2c3ed8d8277a6c440b3a2dd7f9c03d5af59aed7f95c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa79e114222c1decff650ceb89df0c07f0b8cfb613a38837b8f3d63eedc694d58278837f04104c0b2a318d2822b2ed2ba9103bd07dd0f04ef1966a795e2e4ea3168c408502b797318aaf1a24a0de151aa14cb907b60f04ca82eb26c5de361267506fcd7684fbe2f558;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1552a0e608f1f1f8672f60f8f8ed06aafb708e8ca35e0b862961d53a6777c57c468d2dfe75a64c2ffea5752d2f1df9c5a0873d596b7bde6ce7e5132d34e9000b6592ced95bfbbd5a4345245ab74ad018bbb808370b7e767f2e8f4322704a1ac9e92c19f4a817b8a5156;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbcf913963cc9eedb4dc2efba75bbf6d1e060a3d5056bbb4f50728b1173edc1e7c1680a2109d31b500cfb5f6adf731ff915ebefa2cee787c4afa234d50b176bc09460b53984b9ec37571ac3379649dc345957ec55f2f3239792bd81b573a8d08563691293809a6e23b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c21527c5ce3ba3d37cd947fb1c3138ef568c6ec5870946ee44b43ac3d5b4ab0c49260715ed7e7680b94d473ba87dde8b696457e754e3276cc9bf55ee19d2e93cdab373b1452220b524ad7b1cef96202e6b45718b6a878b41df0603ba36f76f653f5ee07b37064348cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183fcf46ca06d7cda9aca03335e9b9fc7bc2c0b83101d333f5b6004759f72f1961fdc91dd0dbda4f7de2b7c98db22714f38eda2858794124c84724ba8eff90c072d36be7e561d109371172146744da6cc6946a08edf6f2cba9c409c139f855b2a5ef0b2a604b825742a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1547ceb3a0920b9ddd2c0baa6f2e50e9106a08d682ecc6bb5e15f620035e8ed90cbfc1aa63d433f93f72abc90067151fa840ce30e257c33fd54d6d9ecd6f9c98b2ee62e8ee10e2ca853bc50f7c84f06056e9acdb0560a0818342a1b381da1329e0bb43f64344c8110a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180f7d86f4286a405b60ceb4704c7ad925630d8270664e19587442dc013474598b38c1f27587c20496694808bad06d4b4d25d0b9a4acd52668978f7690bfcfe95c721a2f7c229202af84661a5008b53c14297238a49aa79c23ff759ec28f07344ab71239b957c528ca1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ff139ba3ecd767c9a8d467d2cdf94b8837a56b4b79d107c1f5336876489eeb98de0d12de5b4eb58b2baccb138c64db603c51aad97c65bf3072e770a28e135fd8e47faa0c65a569c5b8cc274fb98193eee55f340cdbe13cc22abc4d1a77aa8b4ebf0b956b486c5fc15;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf6377e3a62887f1fbf6519ac2eebfe95475ebdd57d118c5c35718c5d2c09da6d3c16dc6a8ef4b536c8b20d891bf6b76e97b4098e72ffa8da3ac93a1afd4463cda08830115ec0aef93ab8c95148e50a5b70970404b116ad12d9213daa9aae17be94b14f497f6111e10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8369d1d2b236e4a59952a8fcd29a415601f1acb4864a6b2eced39d54b8097b8db386f38bf48bd97660850121ae20d5a589d88284c44b38f037f01c442e191136094225a9c2dee4cb0231e28d35a19a3a3ffb785b909b2a1b8a5ec51115dd901962dd40829d577c8e1c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2aca532f88a6e334c8a226e73f823f16dca184655a8438a80d55dd308730206d6d3d56dab9231f8ddf30dc4519be49a6b13a61ee2a4c84bae5f1298f51178d84483834577644478712feaa5677fd98860cb0400753cf0574113a9dc065499c03bf19fa487d7cd73b77;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e25e477226e77a448a578918eb805dc898e361f6bbfb169e9695d0d1154be0d4d183f9298e15d254401ff88c242721fcaf6837c93256f4c3e6ad39f4236f25f2c5f606a5f2a42dfe6b7e16adb82f45273fbca8ed8dd4e7189a758dde2289ee58922855307e3b42aed9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd21ef59b6a65d6fc8a3cb3aa9fe6ada462496b5225e08fa90c694d9622e4bf06fffccec95910af275bcc580d4574a92aed5d9037571ff82864687291dccaafb4f02896aa437ad19cdefba98fc838c8855c89369e1c31cc912094108ae5b5b82d4f3500b9c017d8bfef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3088e75cc9df582559842417377a454a25036f994e86b463817139ea0492b5b5a3958b8788eca873e56442597be968cc7205f8c38f1d4962aa9dfd03133b6add80f5032b8743ee15b75ad076b050613a6478ad65a4d8b396fa01b119957cd953a45de9685815605e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18dad19524f3bf82fb276a68107fa513b3326f0312402e110bce7f3763d381e7ed60d57cd0a1c692ce6f9ccc8c26d7b0d65adecae4f3bb0f95af1e36150c1574573c3068d32e66b87002671e27b3a36148f53aec7775e944f6c1a9cc447c2ec3900128404b671df9920;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cbe4b8f7de5289ca26d869fad533271e2ca6f1a468496a57fdea647a7dc0878a64078f179f08abe095cc285a06bd3b5d20d164473e0086e1bf76dd70d8959abbd27c2696df77439995903b09fec8b58ba76add5af52e8a9d9784d5f2886332b2aaad52346de0a7d8a1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h814a5dcaf487d043bb58343eb6771738d5e27dd3e0a20c7c8f729b5a1272bc19a5a2e7e45896c16cf4daaa3b985b90191a6adf8fe6daed5c6a6cf2c2415e4b4e7378873884594cb339c436018dbe6ab9d4500a2a4a62cf0769749323f0bdc09cdbd0af6d966200e838;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e986cf033b700f416dd7fedef4a0d1ea0add1e32662127ee51e28d39cdad206f1707da346a4a5c47ed2af5444f9234f6bb087bbfdae992a153ef8165e7aad4be67722e943d670eaee01d5728933193cd1e4f9e1dca5da4db44591d1af845bc3ecf10889c48ab9927b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd94c74ff391459fa691e31e286447b7b74a6f4c982b05a6f5ee5e9672e4c4f515d48a96fb8d6fd6f5ff9bd15111cb09611213935e80010974e6d689fb02468a46475ba5dc2bf56800ef66e35707e11a183750719bd09794f410f0865a7e89e013e1a25f32210ee97f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2623e8a8752aeac34c04cc0a5ecfcd7d055323947d72670179cc88406a779dff57eba8afdc2429d9e9063dc16701ef3a116e68d5c245a566364cf8bba6a24ac830aed726d0f7f0310f7a5d1ed3c7009c7fed4053a87b83828ed15b4c15093f6604f10e276ef7d19c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f22c86a06fc26fdcee20f277f58351f6d6024b25122f302889b5b856d0f1f85852195070e8d04c891898dbcbc4fc1490d9a5e83495638264d8f3b715dfcf335dbeb7da5e4a9aa7a09c6624681ee6ee966b182afd5552c7146757b6dd9ee3d54f298e644bf292683af3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dacc297932e1b57485f5c69cfa2adfb53da167749eba9197ea2ce2bb43535ca40656da3666dc851cc9b44281462a45aa4307f2658e69843d060b13348c529775c6c86cfff5ddc9c742a14b04d44860151e35f4e204a28c9102125399dded221c71ecee95010b5d2981;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64b614530ed2fcfd659a564afe887cec4849173ee360fb6dada686946d5d94ac4d5233ccd907981ddd22ca220bb4a256c6ca8ff317fdfb3e240f9658d09b7020d83b6ef80f6668095f31e658c4948c07e56bf7e28e88a404b8840f94e52cb5c5d83a1cde8b299bea8d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdae7a63fd3ad728dd83ce26e33a6d13f865ea7348d2bb1ca3784385cc6ddf2b3f7547bb88c65f5a424ad2c4a16c74f33081b367a6cce661fad9030e448e6fd366104b9c8097987807a42b33ebc50e6e3f298099cc9a8e3fe435ab2fabac14174699aa2c437679c0f08;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha9a11e9047e2813d3e7777c5ad31c77ee74a9135e1afd0d20e8a1f72f2d8942035dcee6234f1932240aae2c79b75538b3e467da4bc717ccc6e827a6d4068409a3ac9927c655100f14df35ae4f0eaa9be11b910ca59ee401d980dd17bf224800e6efc2b3e106ad8f560;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47a934e08e7b8431b92c4b85a33cc7df3f4689ca133178e6b89aa714da03fa7a56aec020ea6642b2391fadeb3da454232bb45ce5687b3646b34ca1b3609595a28a59e9bc973dd81e450c752f81707363f61f9196292e50b2dc65b166a2ff52d91046f2610ba3c1b7b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd359098c914d8ffdf6190127f6406cd0352b402b2feac5a7ac89924e08ae6d319f71776559ba88306455d3a0afbd959332e88a182ba9d13334e5c02d66c6086b48512b05486487cd7bd718f2a05d040563aa7b2da486f29dd1ee7b8a90f2e735e456bf1659505510e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1756bb8428eb3a8a6c92a562636c81268a967011cdfbe6b19297ffa28f2f11d36d6abe28b5d8d2cf979f75023eb4b2f45ef20492a8a814fcd1499c42ce99ac866392c5dad8fb8999610e0b6790ee301cb93ced22e635f8e6ff2c200c5c3f5ea0c629c0f929e1f8557e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f5adc74e7d3ae06c43abb7ebdc79de82786cb6e353db0ad3cd0a5c9b2a142f16ac0b83577abf6832cc37a7034113b82bead92a94e7e947fe940a4ec30cb1034004b1e625a5c148eff97780367f0950394743f8a4261b2ebea373f10854331d1f877f1f195db2e12ee8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152bbc2851ec6cc8e82e18b4a994597b5232ff5c80d98491b5e4adc3c0130c2b12dd72e51dccca64fc5a927522c88ac8f8f65895640de9717294c723370845e45e5820888d6c076203a63e86c89f4b71298a789045e4e279da0d04897aa265c13465914034f0f7b6243;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d4bbd6ddf0690c1a91c6530350196c7c4d60a2b9bcd3f2ff56c62ff0f9c2b1d40ed4f27749b858dd8c431646dad0b186b319b64be2e174a184af60e6cadd4e68bbdccc84d8a8e31acdba46f25563ca0fa4dcbdcccaf55b63a8e139790c84d59a315b042b39f10d715;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f7032b61dfa874209125b6434cf4b0995ed1ffdf8da04e59409a9a11fdb0a631635dcd305af10edc8c2bcb581e7a727d1e9678e7b15fc11f032e7e2e4faff693dca1618ad715efb4c36664fc78abb2a6a8fb133e8c26fa7db9e93a237d28b367938e70868194e6997;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h198a3607a7afe54bc899f432626c1556693e68ff45e85837a5427dfe9ae4f278e5ecc483e5d66f507552aa1677726ccb75289a0a371f2b4580e3122870517e0733e5b633f7e7428bd512e84a614181687aa563bd6b0619332667f4e213a404d71cf0c57fef47279dd6a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5ba41041ec27ab2cc454d78a1a8dc65b7345d3117bd23505b88faf56247a9087233d79634075ffd42a739d693e394c12d1e05da9e2f9003672ac918087a101fca38c062487d006c1b0aefc343b2c0d56d561ba8bbd7a98513c27cdcbd325c6dafd9554f896725fd0ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108be362c56f736ebd933119402b9bac1829b3b8a807434bcedf322c244c1871ac5173d4f1baa3aae34dcc5ed7994f554ef4ac175d5cf7e864122e9769cfab516186cb8e884d31f4aacc36f9fb7ce4e749ead163e315f8ff0c04f7dfa10da4aeaf30a52437302330035;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h627b1da6c063354ae81e7d017c55be7d6aa11cdc92a6f95e8dbefb08491afed08ff4c791e4475c7c93bd344e6d3a7dd8a677fa023fcaf3104ec80066cde7d23f8479197cfa3d7498c148086ebc6a4835b0cb0183ab6a4f7c81ed48cec991472f13533d2af10166bb94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11845ec14e5cafa097de3477f6252bbff7a53d9c4c31e20d6860d28484bb5a304167fc0d00f0796a3285310e47b4f7dea772cfb776eaa764584c049da2cc27ed74e40e3487edd2fbe499bd153e650353942a25e98123edef3d14496db560e17bee480b36667083d5e3a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10134842f9406297e0f67a72f63d31a1d89468841ec14c5edf814bb37764cdcb2d5eb53d0d4325034f6884db8d9272081eab93b0e259eafbe5ca6da29725f353a13b32838295e606ae87d9a067c9ec8a7896ab67192642fcc63e55bad80e680b680acd3b71b3a7a9b41;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c17340608dd99b5bd0c014cc10b90815e8d089b60d8911c47146832df5771624b6a803efec9e2696223ea42f67887b4c9dbe95870ee3a47c089d8b6005461416e481a756a25748aef5e364e08b69a6355f702fc124b883588487e8504c3c8b1f42833ec4fad012759;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44dab4b69c4fd0dae8307881ae28c8069871cb617c39574df79cc62263ead7e0d6be854609986b4fba6ff6e48054f6de3c048e7d5510d6b5814f64115297e1dddd3b0d5ddf64d4fa6c4df582ebfc2ede0e4c5391e1781fa4f421da1ad994e0ca59a5b2621608eb081f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a1ca17aa9443a1fbc38544a674cddacd82b929968602b9d80d4e22a28e6a5e1f0386202856687d0b7d2be82941b251fa7e6c0550486e3dc911da1a5f914cf87bbf0bf5636a3065eb8f51df15bee11ea8e4c48116c104fa29f72b43cdd765de1c781756ebd86c8e7f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h293852d7f4af47eae3f55095fe8df7b4618635dff375188004623fbbdd2c1205f7fc50e337a1d38be7d39982fa9ebebfbf6b536dd436c4cffb5da49582c8c76c036e1e91fb76e44231af7008292110ad6a5abd6df68d51e85e5885c4923cc3610870dcb640f9c7caf8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h184b871ca099903d01724a49af7d268a3d843845605597c220441e6c42e75c2b351a3a1cf845d2c52058d347444409e0ac60277c82b1ce4433aba15c0db90dbaab78b666c3b751add4dec901a8b6b5456b7cdce4949e95cbc1bee77987fe9e67de094662b07105d4e7d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166b00d7a7a3193583fe4539e3657f79a27958a2351f9dc51aaf24038508fe08aeb9319ad0be403662cd8940d04a3220f4bd8f3543efb456ad9fbf5bdd59e7c0f52d8899540e76683f825f150cd68d25dd205f4976d75bd1548266308e9ec106056a595b778a357e012;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22241c890d84de40cf0ac04bcdef25832012929931f1a0c06e68a9d9f3629b9151284922a527fb9fe4ea798b8c1d20a2c59bdeef8a74e813d23bd8a751b9497af4b012463cd6d1743a8b8512c957039047575d05ceaab4f69bb42a755f67f0b1d1d2911746bee34f1c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96ae5d323a270a2b734b6251e2773c55462ab96735cf114008f52b7321139cba42cabbe27965dd00d3ba74fa6b3c3e8caeccf9291bddfe8e87cae64fd11c8774f1043d667b18916dea81511d7bb26aa6e9d4dfacde2a415f2c3641cccd5e97dc2c1a05c54d9e3aaf3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1959f209d30404ac9ab6134d9f61e0e3e4a6ad9eaf95737632a1ee7aecaa08c22b69df3c89b5f1e8f26ec4bb20444254b940046c9a119b90f5afe7167086e7216f0873acf7c1bbfbc440f8965e0577bd131c74918ac54ceaea4082610615f7e1c809eb2fd9127644aef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ecdb430516d3e6f7e24833468c5746abe265bff3720a63250042422d94741bd5ea78251b8a7bcca5463cc70587b64987607edb871a86ad650e9651527c08b6c0bd152f6f36cdf4b0348e8228d7e6d175284cdd4611ac2f2830f538de03a9a61f474b58fad9bc929a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e0ed173ea524ff8d96bc3780f0a4b2366645737d9a8680d0d33487e92d66a7ad68cb24f5f1ecca649c6f867d867975417821d73c9ec426af0810408c2b35d1ccdede756299a7e956dfb26e1a5fafd78a3f593ef07043e1fc6f82691a20356cde9cf0b3089fdbaac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8543b8c9737d6fd6691a476a8e061082f9bfe380cdd727ff4e53495625803ff40065503b3fc51cf4f4e97e84ce5f8fc6bd566fc3020238f9bcf0ec107875fd37cd29f2be9ad82bd0309b516c9d65624521c322888d9cdc8e42a5b3cb73f8e5f9877c2510f4d15f0ea8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1981b5240662d56e52ae573404c1131b86bf5e2b1537e4479fd4a1b5a90d374f26bc8caf1b12e05761cc0aac94349cb0fb66ec855d9f5caec27b200219c884e3e0f079d84c533b4d2879c4779a70d04b420cbf194c0ca9a4f7bb03909233f143727dbc8b1b8539718ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haadd0c596b26e55b4800d4980c7c551a56e3ceef643eb0644b3993583159ab5fd18471dd46daf361aecad319f76893f8dc0320e0c26dabfda8b8c0c1d8d8104e9777ed7b785e8a74e436ba9f201f4f113432ba71935ad6eac7ff01e2d011cdc9f2ec4dae0e417c4283;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h589b0a61047c88da33874e595cdf92f34508b6e3d9c123ed43bfff659d8090b926b5eafec59971b3a885a09d4af00fa3ff655517fef797254805f3416cab4fc2db398374c5650f0ca26ae2255e0fe4110ca001d1c68d230189594b131ff9793001d614b319d9b2c8f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb19c291475095eafb0e2e474153fa1ce25266a9e9bf0d761705974a34ffe935096fbaf4f01df443a4b2fab162ac9cfda4ec10cf57d3b142452b69a44d4fc854ebbbdafa0de55a06cc5076cb7ad87d8e76061e0d934aaf8c122639fcb3a459116aaf97dd7fff55ad75d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a646059dcb1186d406e3a521bc1429f109fefdabaf5137ecfd1820ba038b33d9d38a3e453e81e9fc54ab2171c5e013d15fecf0d9297c6365d893a5a561c09984011094b28711556032798cd7054dea757955dc4ab3e2f93b7291aa49e7ca1ee70c2ea88abaf2337d4d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5dac59a113d9a89489f2d3b99f119b100ed0871b135f48efe979a064f0ab7a3fc1f1f64f09bc308cc04e899807a2cbcd62480987ca450b92f0d58d8bbb78fd05d3a94a88fa3d69cf9cc32d05debb42b199a475642cb85f8ed59e6b4211e043494e66b61ae7c18b5d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149241636a397a3ed267ce0f03a361cc27b091aca7d6f1c9222acd1cb4ab9b27dbdffe09412a67457168d8df92eb3714b4b7b36f5820333f0d42c011da004c5687cdc6a59b7112e3e435991a49e26a9d8edd8088d6ca6ca37745146532e498a1f019d3d3306a0663d3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d567ff0ab47d52008275c6db1fdcc7ddebb20771250d9635b2be44a3eb546c30393e23543d9798cfa695f4cb0b1592ea14c9de213bd8d93379e3b22a21deae020c2c72a8cb9a47c90e43dd12a043f62a2110f9e363270555c78dbf6baa7c8bd1c284cbec50d44e81bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h429ad61876b6d525328a785bf4b79b681dcfe3b73b510b43395fddf9dce319a7091e6f32e200204b69c7e4989704476fc2e4f0d4a7b14788456347eaeb19ee4ac7c6d9f93f5c9728d008beb0484bdab2f71f33c01d32d0f4410ff9d7b8768cb5d21e1acb22891ff736;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ebef7c06ac3e20bb603a193bb525e7fcc22d9ef783519d41ab9a7527c848b56e79695e44b4dca3d8bbed2d0b6ada1a7b67856c692008a00a04b142ac63de29fe08457766b3f186a54efd321ebd369c76543c3987a4387d93918cbe4cd67f1d65db0ea7a0596c1e850a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5da4b4a856e11ddff3d5d5bd2146c36dbdce1efd520fe931d0bbda71dc2dc71bdd9f5db222d2f838125056b3fd9b390ccca056a5827afe34bec99ef9ef6f037ba5a7017e68b6344a07c51b64a22fda09ef2f0ab96dac816a203b722986e157abeb242f4609b92cdb6c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16240f7cd776edf786dbe82352b647d63bb22a4ef8e835cbd34648b9f4287c4354482e01a088ab9103c9b75d5c98204e0e0a93d3ca8f8ee35ad6df3ac0a100a0b0cd4c2311bc9955d1d3ba0f8881e6cf3abf2a249320f5d7a46666b78843d68b44532fe7c53a6fa8e59;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164e7bf7265bf045d63333e3530466ba589c5d72508a694924be80cae38960b16012563591485bae747acf8e869040a5aaedd0a662294876ede2c3545f399cb464983513ff5b56185888ecef6def5b9a823659b42a15d0b31e74a6c716c82c738b299eaa0f1b64746ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101dfc6c36c971643b8eff318ea30773fac51179143791e9f1e278f1b19be5f10ddaf6a2d9351956ce6333e39c5dd78113e7d761b82b20c67b554a11c5c9f0629b03298f3d267bf450527659dbbf591a4415f1c15e63d1830c33b0cd2b4cd10b3bcb801e7187ffa0009;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18374e5ea17188ed1056e4d2b7d46a307ef078959b650de416f0744acc8ae83282d7386a2e82e928aa96e659e8b1a8331c69ca69b09c7fb027a2c74674b2b394ca75820269a490e49903a3c1f0c015140eaed3a9359757224520cbeb7e5750494417037bc721547a38f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5666912fd55c6b4bd947942a1a49598dc576fb5ab6b1e73a7d47685c778e811d208ad22d0ad031ec53b41a91b8a43a8396ba6935dc4b0fe4cf836c3f3ea84a136ee9fbfd50fee491654a63df6ff8f4adf2c8b51da61d38fbf40f58d47b9d16af4c693727557535404;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf60416d38fa5b55329ac62ba85ca3a067961460cf65ff60e8eda1ea545c5b14a4fb92528a458c38e346d3890f22b32307ce0cf3d4ab78769eddf8248d6c4ce2379cd2759a827054b907c5b21729c826c7ce60cebf89a6d57a63266cba058273d996e8f0f4a65f70a29;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf995160faeb710ba29e4b8d1b2c6314863a4f82eecc4d1418bf1cf4c138f5b2f4d9a01270639b9d80b0594c54cfdbbb54625bf8eb5ee4244f99559f2f3cafd831c90af18de5bc4b6bfb40ff689ad5635e17a37af99b115b8efbfc9df1693542817f3b99b414fbd109a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1fe56d970457c403fc72f3dcfbef34686473739fddc8bf450c6200b301f77acd8e44f107258886e4451327429be15efc8310b252b4100952193fcd9fa1a46903758429b6687c11a12f0c3661a8731376b568d55af16670ee9fbc8fb9e2a52a9bdf0d3a2e6431fd534;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd76cb1e262d88dabab87c9cc8cd76b64f8f841a334ecdad61674b6b28af584542e093f887476aff06fe91d0df8e6ad4e375147f410673a6ceb09702484fdfb1c47f0a3ac477a8eb9e66ff06e61f5bc2037ac2537452fca6f863d0d138f55e314ca261cf63a79f42814;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c3611865c6eb2df97e011ec7b386e363a8b9597ec4b8abbd3c930ef6566f729b3c81165ce60a5809ec8f948d286bb6c50c5913859f45736e82a93f8f48be7428b82367db484f0e58f3eac31e547439bc8fbff4dc9da39486f46a500c406bdf3bd1a9e4f103ab243a95;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he58c6d557387633a86499320a19e16b436c375fee63b9433bc944a611bce82f07efcc350cc2eea6c6f434b0fd10c1915ece810de93fd0137b3d4798c5b59958c7eba9fef9d58a651d06cc43639c2a8c5b154bd70494fe416640da79efd86d353a39a0b598e454210c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he2a73c3db66df1607e8336e2e55ef5b429275aa3b1f1fe79dcdbe56bc5024dfa489fd01821e92439cb3dee01b3b2c026d9a0c010bce96f12a872ced10701637f3cb0511fb9a7ca1abd1109a029ea01cc4de83ad3f6bd19af9e778516ab2a38c9b90454b23a25bf1f62;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42ba4c990a047a9bc5c752d583921b27dbbc6e86f9aa5dbd60c2fb806cd7853e2bd67eec6d2587721bc85e05a531ed3991f2b8d8163e249f45beb0e7f02fa421f7b24d05343db5ad4fa0b60f241e805950406c1b09181898014e14e7e446b0ff1265a428532ed53814;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13749a15e9d7d616637951ddead3373420db2bd418e506cc463251c37a12f9d8b1ada4c5ae8053308b7c88910618aa3a572aeee9608b79b8ca9391f7e671a95866465598328241037dde9e35c026ef3b2169c3e9a6db28e2c85fb60900978afa81e3a06ec498499b7c8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79479dd6a500eb5734c278cd0728c64145b7019f2168088729d382abc37259ffb434ea44cfb1efba59e585e7853c7936c5c249e4b3c1b595e5a094d1e32a1529f29d52d7e05af980fbc36a017fffd681c0b22dd1206d2c42a07455ab0eea990d32084274b05feab1f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc01ae978ac8a0cdef2a3373b7015530bb6387feebf85873276f97f0a2be6a4e9c2caf0c07dd67c04cc5ffa3ab6e51cd7513fba0d631be793be25d7f0a9f5e4970bb860fa4f6acaea8b8535e5dbcaf66b31fbcbbe522334382c58d7b9f9e7def899113d2f4abd996f11;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e3be3dc56d1300b7ba6b2d785d97c5edbef23a884abcbcc0ea57980272ecb62db2a8ad4b1a21df027b3ea52de7cd7b77984b1454900647fda7b0170b4ce20b470fe614f85b332e990c5fd7e868434d4d3b3a99cf0d0614bd5aba21655ffc4ce7fdd556ca551160d40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bbcfb657494f44c717c024d7acb93a86c42e4c54f4310ea769ba5bb8be58d4360734fdccd2408c036cc88cce0063287e16c092a941510560230cba66fcfb86221d18f19f00437a9ccf17805a4268b08e246eb770b84ab9b4a51b78c1f5f019ef6ebac24d83d370abd2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee5520c0d99d4962fc2211e49ae9aef772e3b389712ccef0c65c3a106eec6bad9aee744e0c6582a02d0e91ef76cb4773b967ed654536fc8da4155f8882088ac19302f712b1d78b2daafa0d7bd2a5aef38ed624729480cc8e1009db9c0459dea38468d88b164671b21a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba994c2520734b4def4d6feb0a24de59d3f42771ab71e0290234532195dc21ff13c8df11f6d04d8f8e796aa1f75c29ad2c3c48d9f0183ca0239e291a3111a601be9f3098954264e9e2c1f82f886dbe39c43fa5fde37290a4c55b11dc1b4f536187eed1216e4ddca1ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d36eea044552670f583f34ccfefb1eabb484bdf6f1b543c44b83f34d9483a850d5aa76123371dc9fda5215c977307a68125e96d3ad13188852c7282aa34acededd1877d381aafa53534d47442b88b9690a6babee22667875509eef522dad4028dc89fa894c1dfe06d4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21cab8cf1e63f19f807b057b767ed0320e5e8395e0aba586682dc61eca42f3886eca44e37730dd342c7213c96f0418a7e0bcc3cab5f94f2aef2aaec1e55090747d955258793c306a13cf261a73ce4af00ac3e043619a4c058f227c7c87ded75e2643ab8a73c1b02387;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13cfca1278ef464d3de34fcdbd16c19c13a56a9c5126125e7a7e62ff929cba24736479d237aa1367419872dc7ffc9929a4e30330db8bf67ab877f6761b67bfe1de842f84418c4b4ed4e4515df1172d1fb6d3a87135ecfd888502d529f7c5fb228ed2fde0d19c451ca2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha67487689f183f99e09836f26fceb35b10928e6ef4dc1cad0b6a60f2891c5c625b0ce4667986f3c5416fd3ad1b83e44a8f66576b86f2f678902d607298b896fcc887271624a8f7b47e8131e02feea1713b17bd5c393fa02ba4372d07aa6d1f303b80121c30ae17c974;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144a53dd0d3bac5bface317cf3280e6f7a8298059b4882e0723cb860e051debd629d401d331afc56dd661835aa0ac00d9125341b8f49c41801d18960ea49590073aabd979efb0b2c8640896d808def46e58b4201c2a4d1ae810072ca07eaf4e9d2f3e994b3518382df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1305d9e5a631414ca4422bb2544253af3416ac7b042b36ff778c18f8319870504c66483f0bb1d8d467651f36fe9fb57a69ae7ea84c493e6c28d3f9668d122ceca07cf294c6ac17935fb3301789bf1870577e6518a47ed4fa175229773b0dd7b9eaeae4ff1243c2e3978;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha45f3a8ba4803fbd3036c7d83db8d8c32ddca37020be913ed15dfa0bdb3ea630cbf08b29c8bbba955ab940cf1c0021139d28de6ec7c96391f3959c63d685b86bd55b698dfe89ac9eb9f3e79c961865321666eb31a984a5e3b1df7249e433ad0f112394144c5a295365;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4dbff4d22c02dd8102e022d2147e1a02950253e82969ae834d5399d9fdb21bf042ca40c254b502e2e62896e52ef50062c3532dc64cd6da6aea7c74e87caca07eea2aa8b7c1712f6dc2b359573734b88b1761d9c2b1f21260934915e12ae08ae32314319847289ba431;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h97c5336939693ec88695f4b7abd7e9af0cd7445a4127c5ad7d7da846e7d38d8d11db81656ca482cf144e17ca0bb63288b6fcfc93235372562023b6031caf4b11f374592179b2336491d7198a84e2f768874352588c74da5947a40cd2469aaa8420443d700907a902a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haeb86668372ecbe4a4f214fee3763aa4ce8cc895e640fd7170e4cc3b94b228fb62f647a580631fbff061aaec87c2d251a0aa25ee295b37f8d62bbb06a4ba64b7f64f191f48cd43c2003e59f4cb8bd6ddaee4c15fb4fbe5009091d30d0ca059593d6ec7cc9d6c4a504;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10953d498ac467062aa6886a8df4233d1467610e8fa5af90480c5f018e30723ee36433293495a1d99fba13df99cb2833324b1f5d3d30073381c1cb17bd6985ff06a2373b9d6686436f9246057b74f7c7a77562ad77d5e34df3cc076a0043b56f429b1cfae33db481117;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1775a061be32317b05cc424c37d482230924fa99eabaded0dfbdeb41fb7b86741359d04f30bb0085238a4409c756b2e9306d43ee981afdaa6c1ee9d8158c6949f45d126f53ffd8d385c5bc2b3cf515294416731667cf2cb5788f677e2cbadec0a800ce9a1b23fe8c634;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had266d1af4675ffe10363c34a585e70ee9900b9aded0de2045672e76e49d55550a101a3b3ddaff6b3702b82ddd1aef4abfd9e7a8281bc8a5618901dc6847e7623ec5460558e79887087521ec5061e2b50e57b5db32f86571b3254c67e7e7d3f97ff44a68c5441ff6ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb44c241778b36fb3e41a51fa6f3a456782cf2a721365f62787a2cb9e121db61621fd12796c063fdd4701c7fb39cf4ab90a1c95e910b88402afef786a74a572247d5d66694f393c956505eb42716cab6e109c564b33d39e9a35b55ff4645ba216ca49bc131a8e8dad31;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192ebafd58e9c99bcf6d205972de2f1d65b8108a9a40255f9440b0c48f6c891f93bac61dadc4f7766fe2637c2faee73faba6a3cdd8fab3c066f4fff3d8054b48682c5fc49ece1eef3cb124449d54d9eda663a5a680fab747d05e1481c34baefb903991a2771bfbe2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28e94b2746ee0abd1abb767cdca64218f8e99c9937a7fc7e9bdb62cfbc6765884629db1f762ce3db37a5ff9cd28b1bb68cd07f2cd4aed8c254a5cd8fced0d52861ec03c4ac7324ef7f5bae0bb58095622950cadde71e96be763a22ca6f1d1cbd71f8b54cebe100c6f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d0b5e56fd98af7800117b0228b05a7c62a4e7579c7670bde9fd781174b719e3f1ba997869c4ce324b896ba0c39a97a59e6ada0f648de0e05bf9690beaf36f4530af1d447bf28c0b97a2b07e4a8ef5112365c1f6a87eb29ff18a9271417a32591d09d679f90ac2c88d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h639a0c360d2c13ba85b8a13945c28bdb0645e25dc1dbe534d85da5d333deed656125ec427cfaf4b1ba70fc14814aaa69dbd55218b62abdc4bc96d4a5a7d4238ef5e5be903f3e9c5b353a129d35e8e92727f4d579599b2094ca8623ff44b30b29df01ef8c29e7604d4a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd9b8ff515cfba087a07236bd8009d08b384eb3a24720e789c9139f6b170e55182f5f72bb135a8aa742922a3b6a18936e01bb2c51444df546a7555418b4c8e3a685b658cf87cea49066ea574902745872ad53750e5aafbbc46ad98badbfe7602b23cb925147666e1ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16730c333bf58ede06ddcaae65e732d14059213fb2c6c70a70888937a5d6d0a1ef123914656997924679f4e81299f987c6aa838d608dad534eed18f36face6722ad81bdd1755fd3eb8a202307e892b56fe8ca07caae7c3df4fb1ab4a892b1dcd2898477dddb48d2f199;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1a7b1db087b7ae57f009cd8755dac4f907ca01fc83b3bf9eb481bd2110d45f6b58d5b60cd53fbce7c65f3f28ff218c298c100ab04f3fab95d901fbd90257f1401d98e771ed3e81cb7af0954f4ce2a3ce5b62f4991422216d59650d21e0c83ebc00571e8fd647ac9d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6bc2923fa290cc59983c59d3aff9ce0bfbaf7e37e2abbfffdd09925925dfa3d0eac95fbcbd27d4f7c629595adc1827bfd073676360e145ca229b9c8b4c2e90327de3d00e66844cbde25e0e8a8553282e500a5e97c5c48b0c8fe91d7b4d443af48f5f16acaad8304919;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5736deb80b0b79ccc8b38ad47d7b55aaf96f803b5eb5a51a2eab011576b45ef47f68a78e49e54285e85a48b919208308411776a16f4254a303d6a8f7a071c5fecbf080634f53da5483e070e9dac8dc0601e6f90f9486ac7463b30172b782ae4f49d925f0caf654fef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15bb1546dbab6e0c58b97df3ada29b82978b907fdd510e1db438e8b55271cd77443c63a54099854edc1b3b3f143ba3b3d8d2a3d67af028adfaa63c1a1641b25fe6e1991e76dea63d8f3a8ef64cb2ce5ad4560048ab840d0b7e1d77e25f460de93d1a17d8c3d26cc7185;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea9e7d26e02de0ff87a34990a8b841874a8dfbfece6fd927952f45d9e761f9c9d67be46e61f28a4335819e71caa6b8269edee556e37401ae7a943d567afe0abb1f750fe1bb9c2fa3ab36af1f36c8d6fe7407b526fe917cc81d44c95a6c9020ab55315eb7f312a98abc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e8e4903101a6315c43b23b1e8dbb36ba784d5cc312c36afb0276a5ca690274b464fc216c483ea65bcca1b7d8d2b79abee27b63d9a7c8e56d77cda8e3899304a7d8fe25ac560ec08dcdec2899312afb689c1306df49324ca6faf1c5d966a4c495484c88ba6528a9020;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee1bb5e28b13e4a9e56b747a16ff66da8e9104fe12092a3d24edb679b12139cf1fa20cefdb32d00bb200e9b742055e98f3e7c98d62da7f7f7ecf0302684f1d6f57cdaf284d777ba3b7a6fff230ba52d1b2b8112a3a70576deaeefc083bcba4caf5c0805ef91529ff16;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b75755215f7b1c8b4d930e80c5d7155c3b72e94d9bec3b9e458387b0a9f48be190ccc5abc0e927f19e756e3f65483aa3af71f9ce04c6fe86e17add32ae3390433ccbbd8bad106cf1e17527877ef0f4d0b34f7ff961274865c6471f4f9ac19f59a3e3f9c8222ca66478;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd33136d577ec1381710352eb048996ce608ccc2e23ab8531f0c328ae15802921b5aa2d7e86425a1c0a7337149017cb9180932228fa84e87da0a25517da7e1ff3e0ff965e28e7adfdfb3ecd44952798bbb57ded127908863fb5fece0dee1d626c5350253bbdea992d40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h87a5637092c168fee7f25163037cb5ba4f99082ec66d44545e32462687a57dc987aef68dabbed7cc4303000dc8351b201b1555711a260f6619e5efd9a7b4786f1bded173c34e14c5315d33661eee404107b09521d7d666d865d2929088370b607d3767a145287a70b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140f458079cb808fabfdd8203cefb2a16b520cd1cd23166beb8cc893c5b6d07a48041adb3d7285a61c326844f29f3f7c24e6c4b11435b77bdaa6c03291b89f24c626cdf47deaedc4c80c234139f15803fc4e1fe4ba6f4f50ea8c6f9979641a7b8dbf40ef0201d6be07a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba5f91d3a3ef65ed94080b4f812a0729b85624d4afe04a7557abd90822057cb12397d5840e1fd9387416ba84e895ece8b4ffbb7a029f8bf88bdf45d966562092cec1178da1c624f3cf47c26e18871d1dce223c6a669a2f53e925ddb0bf4f88d5cdf51b29ee7b26267;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177df8f5b243225e00456036d35304a4b5d4b36b9d0a7eeda37ff2186b11e2c4150c963d2ea2c0b8298e6862f59634a2eafec4e36eb949609859e36530341ac23dd4da3b84275a068ab6ff8e49e6b07f870665f3cad4e38db8e5b43b63e38a6f7432e9a7ec0db9624d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160648db1a8e2135e18d6577719565cb0b055d18932b4be4fbbd0c8b69a6aafab9dc9f8e8c5cbf22b4bfd86f570e2c082f0c2835e5355a55889af78a4a193c9f25a13294cc0158581f5dbee52321ff0eb290bc9a2cc9305e46cd1214211834b0cfec1c3a2a3f84fa1c5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb1d2bf8799940849c429a3c5562b9cde588e9ba035c5a03193b80a892f246eba8ca67845c662911a4137b73d55f41a8d9bf52d2b297208dd2d61d764a9f00b7f518e59a7de544728df81927e90da24ced036c8825159e0a97528acfc98105aa4b514d6591c1bd3b36;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee965bbf98d1bc2bba9d079546f8f2956437abd5b7266eb1562090a8152aae346062045cdf2a2fe594a403f5ca118a6632e5ba7353a35df3c2e168e18a681bb8c9a928eaa94055befefbe36959693c0630d469de0b5cada9692b026f55e612e6559d5acea844ca90a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3938403ec329b8e9ad8e38ea34bce7ee06d372bdfe74b3c2f007411d6c1d13ca81c0776b4cd2d7bbf34fb34e5fd1b4c25acf800e56b6c9fe88399ae5301e786644226a4636abdefa57bf9a790a97fa7868b7a358c536233109fcd1ca2a1e949392bd0eb6c09299f3e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e9d9be1e9298958c490b4705aff098308dc17746aef972f3251a67cb6bf586682568e2211939a3d5cfdac929db2ca0e46082ce86b112215034049d092ab319d611c66045b76840177c72c229e6e2b7f30cfb2687c61ce97f569ab74684f459c25d6e886efdfe0b516;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31974c00bef4739869704dd4d20263f2629cf6a5a5118c5d2c4b8796e78f692ba00c3c925c936e1785043753780104ce7b3671017ddc4937fdc5666bb0fad92f8bf802afae2a203e0c6f6033ea6997df7b98ac5f7cfac62b33d8b9ab2189264605c40a5c32344728f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101afb4e711bd485d94546c7328e088e2a126363956234a66bb7dfefb423a0da593415c32d55c49c0725b53138282507b37af7ace6dc84392d797ad29653f72821a112759e2dbf745a0c4245f26a168a3c276f45fa5ea9283c10e6c00eab34c4c62b7659da1134af183;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2ded97ec7d507af91505ce49d1588845dc29d87cfc0e4142735fb63c979092a03b21ec3e345519be4d583667c33c2e9db9ebeb9093bb4807cf61638bec59c60ceddee4ab6d5d62c288977563f84ca6e2608d35d2adb2c15f2b5ba8fc333b2ffe69db09fc37b0dc3037;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc618ea307dff029fdd3175c3e8cb8e64ce45bd3e7d0b58b22c2f43c77c9c73360b08c1029c612d8484f7590909bb6c341650044cf1322a538e02ef170eebed2edfe5f71f29b227fca1925b7d7721ba87aee41fe006a9fbfb4b3357a9649b852c5de971efb04d31e145;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hca8d530765af43ad0003fe25526c10d2e339350ffbbeb87a6c9c29904cc5c69538b28a7a7126b69314f225a2ec625056d6ab5c8bf51c376a7fd3628ec790972c5e3bece7307e807ed8b733a2966294f4a828b0d88e1567b15792ff04781342fe0e775ba9c0b4ffc159;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bbd971cfbdba8da0560eda83e45e6dee18be118039beb2f1a5a1edc47f29d44c39a8cd6efffe89c0a296e030db9179ed2085ea6a4250ebfbebe5db2d792e2ca2eddea571944abc28ad945634f49483bbb3e9663ba3d214bd8c93eb06e867ec477903ea36e85aa1b18;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfc4249a85a3bcbbcb45e1c6632dd186a1a356c684717e17b941011882621dc0851356518d278c781c1c3b504b63bb010ed5d41d920f1aadace1ba99ca51b6a1e3a3a725ebeb2d9bab82e573b931fa17b855f9bb1d2f64dd6b679c4dee205fc89af39b03b15f0124b13;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ddbd961f9ac06d8f34cb49b41e253407d58b43c1490a620fa850f56f18e9b54ee83b29e052c392eb6fb2465479f8d57a0baed7799a6aaad6865af84bc1a5bf07924be3c241ce6c485290787d224b86a4ce570bfc1723d0600df1205be6b4b37a00171e2f330560fffb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5135ed2cec42607861b62f361f027eea41a5a3dda2af2e375c03995bf93e02351037bc25ace6825e673a466fec2f01c6628f3a27900da209ee932639ef920cae822347f1a961fb68d2eb7d404e56c904dc5d3b0cdc32dbb8a5bb17a30835ae3c36f00128475f9fc7aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd8d9daf8727d0b853369b4a8bc3e07749df9eb5f55a35654054a22126d352dc30acef19ef98afabd3c0f4fc92d560febb4441e04ef29bf7d2dd5a6a8c30b553375dd434ebfde49961387b23e0eeaa66dc73650934affe81786ab04363d91ec5c9af44e53c064ad21e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d6b300efc474da9ee1f1f8a6e0d940dc6e4ed3b23c76856c63f187d6ce0c0e3c3c4e66f2b60bcf8fcaecf6631f430463fe7ac45f2c4400e615af366a51e83c878b7ccee192e3b390033972ad501fb30c5a8e93588eb97b0582d1ba52b434eefec4a037f1c843d7838f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79de1bc0498043e6af4cbedd50bbbfc7bb7d8ff922f95c14fc005285724ed0fe10fc4f8aefbb2f857e1870a057efbf74dc354b092bcf59bc5c6eb354d58766883db54111e8e8c4ba2932f694dc177ec0cf06676e5ab4cf08ffd2eaf04f70e1325351d4c72966b2a11e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d033e84667470014c10816369f71baa4aee1eb4cb0c2096fbdeb750ed792691e41e9acffb37c1a6c088682bb176abbcf03abae0c6800fa110f61a86ad08c1abe4a7c67967b778a316a8d4dcb28d39d15963651841c495333228246f2a3b36e81b45bc462e6d4f1a624;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haf059036d4f5554987436cea9f27e7fee564de93d37ea9347086acfff789c85833b9f24fc02b873b20a490739ad698c6eedf309f64e767365678bbb26692f7639cd13cf27eba252c54adfcbefbd6adda7e8de2cff7bea69863604a42090d94c27a0b8e619cf9ab3ec3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9eb03e6502702cb8aefa759a9caa3b89e8dbcced01399d207a3903678e81c793549c8f035c30e67631b89a66a60a3962a8af56481651e29a76c57a84505547807c66ec42105eb98bdceb983fd7f7eeb492bf586c3a565eb3f25b7f03adbc1319b7835a8f3e936b8300;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1720cbc6abfa16df0c71d4492288c6ab609860453393de80b19b66fbfaabc559de18a23a1e806162dbb24c6f6b62d049711c6cb8e6a21719da97eb8ebcc103ce60a2092d2b90fbdf00ff86e22eeaa2c127574caaee1eae35a17dc3a7c686661a08dda1eb88d21ecf516;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d42f8a6cfdea1e5540cc70d06f0635ad8e4e3c5bc208b44e1b1b3c552eb1e8f5e7b0e8af80321b28045b3bf7054e097f317edb530f9f56aa38c8f9360fd5a57e2a3e92fbdafc79321a150cccdc1ee8176642f0a3478d9d40b3fe820e71eae141afa04164fcae1eaf9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1938b71d61f421b596c69350170ebda739b574fb196f791f756655ad50071ae978a67455b99b5c48b70e9ca344b74f67adcc420b416477cd6f37d8ffa7e4cb3534e6e4042ee0f78413d53ef8b100e9b64825092bc77487086d3dca9cccbb374a5c96fbc5fff3a1719c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fbb818de5319c199cb4092cae7b19c26a781252236cc6a0ed09be7aa818102f8cc3dd347675fcf2751a76eb8e6726e7327065cae346d6993631e9acb4543ec4552a71243f8f0179700aee802e05587af53ce11ca27617c13a6c69793e32df6b09ff500cd7c0f4eb9a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1567f38044cb55f105948e90219835c525de17cb731938bdb9b27a92fd6be44d8366f03b9ebfd205d96b0fe8c5a77686302de5364d1c4b237138bbe82fa1b6d2189dc68c48fedb23a13d57de88cf6237b813b7438f844d4f6ad63bb424e9b901010e7ca1384476e501c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h178a45c01efa3a197a20c4736a6fd9c4016711d1416c7f5a94d2273a32d7e2ba2196c6d8e5972a0d39472ace642c80aeafd1ddac3f9fc28fab91aa54500c3f87d99869eab98981e834878d8c70ca4d40a3792cbcff87e1daf4d11ffacdcc9dcc5c714b6fb3509542adf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1963895351a4d74791524a764a0895bb9436050d34c3399fd41ebc3873f01f2966506309cd9ea3a264a7eabdbf9292e626f6d707b0c0b5805feeb769432318d21f9f102759d162021db94e5aae190cb876ff2a34d0afc5a58e71e24014f28f40833934d44cbad40616c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h23cfa7995683a3827e03cd532afdcb428f8e93d53bf640b3e8a58183b5ef3520c5eb496deeec2eb16cfb12eaacb5bce58245716796c5f158487522bd7f50a51f3a68299c8d056f0cc8979df912e93b4ff04d61984dccc8562cce117384201f0183c4ccc5cd003aa71d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38462708a4a924557a6d4f79fe1adf90b3bb51468bb7370638c9e5ec921580f61f9770e8441cb554d3548c9d28816067d77e4205091a12d9f03cbf79b8c805848ca3ce2ffb0a16d1261ceca8eef69990035fecc999c5c63433cb9772be38523c00bb9a100a85c51981;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1633354cf8b7e8c3479ce4b8569a90b977fd6ea3b3673b89d2420601030ddb3952a008262b89a2c91b8b11c7b188701b0e3d039927debcf2f47239b3e31634c29de27973c7fe7e74e19c596cbfa330933a5128bd479185fcaab1ff8e36d649281dc5af7acc8de4a268a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h176410233ddd892d7e4319f828efd19d982039d4452f730715aae42a4029eb2e9da9efa948e3f1c66ead3abf09a559393b247f192d81ed801238cdb4c362c26d7a3e0ed395fd06c515778bf37d27afa86b40d7cd0752e536c3a2bbe45c3e5d747427210a9ea82d3df1a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e048dfb9b6a97f106a17440ae4a7217531868935e6ce9efdda31459a98a1264f01e80ce1dd46816cf2260bcc9acbb1345d7f30448b694210ab2671c26c6ee513b5b0a9f03b3356046fb86ec77414a8cc5bc628d3a9340c6dc1c3b455812acc9e1c5f69369b37a1d22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db1629582a09c481ad41b375a25535618732158c12d141d6c6fb467ea11d2752ec3baef19b7d00a14b2eb528ee367b78174a46e6c96d166cc5579c60fadd79e2dcd94e7f9451ccfcb5d1b2ee3c61651d62752084cad9f1ab72dca099ebb425ab72f3e92f9349fed950;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11853d4379cec3621a7a4eccaeae4695b7281c064afa77b26f42322c6fe944181e2c722d1a41ba52e6a06ff77207ef03b64a738e0de90fd1a2ec0eb0b185c60fd7b0e3c374a6bbd2e4870c7f12057bf5e551c83a7bc9d34d8204767983a49ebf220bd2d133590b92803;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d1430cc8c344ec190bd4fadeaa5e5bb92480abada83d9391d7c964124f00cb41a48860cdde6f463ae96bb10045c9384b146be185261bfa576779b2e5575716f91292a9396f32ca50519982abee18b352e01fe34e4c31afdbccd6bb4c17cd355e1740552fc1adef7d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a56b0bd1ec4e54abf1b9aa68765b5ad3e8f81c204585b5c7999dfa6bf46625fa2e6837b4643f63c6ebbdd270599260547aa6a7febb0e5bc28549d326ec06c56ec9a135e4b8256e2f2a8cec43ed79de2a8fc0e32ff335d1a843fc8ed6775da185de3105a473070cbf4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15194af0017cf0a970364fbe4d98864c32332ea2a0f29ff892f5e4dad4c009465477c47d1af8104d6bfcb2e8df70664bb64331af735a11deac02f5d171513b7a3b8d01cfe92361874c8aa042fa6c4dbcb12c5ccc11dbadccdabd9845019952a5f4453fc41d780c95a94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cbce7f12c324a21fa1847501640fe611a1b8d3d15be4570e9ab79fa0e89f363617d74652e36a4bb39810f6a4a0a380e46cdab0da139530cdf5f0c09307373092350c2aea97e1fb70b592d8032af424924ecc3f47461e3309bfd5ecc53f074368455ba4a90b707a1637;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2cdd4f61146bb0630b161d25b97bb1d2f246b32871b524534cb0071d25acd1631259ec7c3292585a8410ae4b59f5bc6b4a6a54bc6b8db4cd2215504b6ecb14cf61b78e9c0b372b376013b6a483fe9df2eb91300c12fbe4c4fb15f37abe1cb50a426805f145ac79fab8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10fc2fc9d203ebb10f1812014443cec43e7d03057d1d3b404242fdfbdcdc41c7c1e9cc1f6b92c8d8c482f76a8cdbedd4137df1e27ba7efa7fc9b246fb2f6927402aae12764ec84fb825b38c53632cc8f74ee206598f848af90bad06f3abd5a737066b0a9b592d0f225;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1720dfbdad7d7ba6107b50cf246b09bd0af31ed2ce287590908e8e3cf957da67f3ddf453a3baa48dc23af3ccbb6c19f3c8e98c9817e4fce7fdcd3abd3be74a82eaefede1821f3d2d2ee01778a0b69d87c24f77a5acf93cc6ee0153b99e7bed73fe6d325e4f7858fda4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a5c52d1e518a2fdbc13cb4351083faef3795877afa41b6f6928b58237b05d565d474d40acc6bc6644b57d7eb7a4320a0b2ebc95ba0875fb2a47921736338a73457d6ddc405f3184ef0bfa1882465e25b334e275b7711b3e062bb526e4f194b4a324b5380196dafdbb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e5195fbd6b9dfa93b9ec14a0ac1c35b390f9af6c861b233aabcf8588f656acdd2bb200f0379de6b6517cf60500b681e22ce3c16867333dd3d984e3cf7467ac55bf952e0de76fb006188289af838d02745c0317c109d2385aa042fd1681365d33fdaea6bf4cc444fca8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1142dee8d7545ccd40baad267a78f5e4353a32db4782c8f37069dfc1611b96d7b27ffad20b2dfab539c90d6d7938a2ddcf5663895a43b3903e74292d6721ca60e6d4584d19f3b3c56632bb352605a3063cd2b81f9e716850e3e03e7417f6db35a85e0d05994376c3c3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7abec1301230a616afd65174f707cbaf844117da5b1cefc80f1c7c12585865147b56a8b54bce87c15abe862f73d4143e7d1d683cece0fb2aedcf56c57922a14acc226a86e5bff68049f805d1b1b235031ed26934a2311b3a30b2b10f5d8a3f05a488368bc1ca8025;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bb668ef9e46eaca64f8f593a98081de69305fc68efb17ff4118fa8c38dca0c6353cf17eba460d4e6dc6a06424bfee7e78b2e61ba6af88f729abca8491e2275d7ab54881c869785285bd08337a18afecfd9cedc3957ba877c072e18bb85706cd6775396cddd2ae090b2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3b36fc1bc42e6492344effba0e0b8502e170987c3deb95dc068625aa099ef005d3421b052f396863ff9dc6fc78983fbaeb49d044d75bb6675dcbad84c874312f8787648b111c8006ed4ced4e855a7981e7b2aea82b9a8a84764a0e68f16911f3f0529a15deac7c9a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15a50989906b8d7d3a1b2b5c4f6517d06b7ef61d85d1fa83d1bb90c2d900e4d5391def15df0fa12df73752173b889cf92f7b3e65f438d5bb9e6ae4f0bfaa9898372590cc54e761ea15ef466db8f07cb3c95be11992d107de55f4b5f5a94d0a2d56d260b8c763d3441fb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d61fabcc9dcfd8821aaf5b9918b9a401e411e080201d2f0de9d5742ea0637822709db9b5e8b190b00fda1a2088cab335ca20aeff77f81c6bc11d750e53014188815b74aa14bfcbe53680874d01bf2e2b4579b90bf3f51bfe4bd6f2057bfafa07c92067c6995402cb3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16b1977ae8e2f1716e1d4373ea53ada1594204d9852d654611c3d12484918688154e71dc082de595108285066e033df19c2904495e8622cd8244d632be8e8c0022f712179c3bda2250cc247d2f34c16dbf9a58e426f616a9f87a3a7ae1ccd5dd1d813b2422687b245e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3107fa9ef08d28989cf5ed5439673a04a0bf582571ca70716426b72c40d4c0895d8cf634817588a7406ec112652a73e764a509a0144e80b563934d02162d3c2c318b46f1c0e31069d7f8bf91586dc3e027ff404ac6aaf44c4cda546b3c5babac0522c439e8f1d7631;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h937cc4fd9b6bcd76e437c7082b797e959c486059542b271ac5f57aba86cc2baaa5e7d372f4cbc56f922d5db5d50e0eb440d2afd3f5fbdf1c31b1d9c2864edf71b88054ee620ff936fbf356fcf71a25f0f98f7b29e6ccd6f5157bd10b7073f1b80ad2bedd510c07c47c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1073b181439305634cdd321e5e231fb50a05b9ba069fb35f163593f4ea87218a93d21e5f07a76d9739393d54811706c2ea723044377f8c040b6bddc16041ff5f2787bf6b1139a7ca7ca72535b5adc2bf20aa6be26cc09d8c1ce3b84702a7e90d685829ece15033b8379;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19826ac155bb45ab0feefed6689235c7b96992f9523a4dba28d5fe6f593f4c08b0a7648bf248b518a0146f3976aa2061a2caf8579c05d6f1dbd67b6fa90962ca9da3d0108439c0b54a887a26eef310afcbe2de9c0edde38e4b277c009cf8b548f070993c868e4e83a2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3502b8d5bbbea685ed7cfde4f27d5f1f8c37310e8c72cff479350f90baf65b08724fbad14eb363ecd0985917f95c0d62ae2aa134d634b23d7f2d94077643ebd0a442f378b1aba368301eaa4ba0d85f6dce2c0d2ed0aebaff295022c9ef8a4b6d1874f30fbcb3d48157;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116035f8a14f9dd3b9e3e8f8680e134cbfa55f9c8923ab76c925d65b425d9ca2500987d6d667ff30161b883fa34f1429814056eabbf7b523d620cfd8905c64da854da2078179e01a8880818a6a517d67d93e55a0369bc5d4da630da3c19745a0dbf5910dd71c0f8ea82;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd924ab2ab0b916dd09ae0588b9ade57be054b6aab300c511d897e6a914862cde30bc9ff24bba9ac6a17a6be5a446f8f2824c71778bbfc84305692b29b5e5a60cee02d1b214e4150b42604e4625b43c8892983eca49e224bb25198666b0b39d6e46d65a2826bdab8d3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125747988f1b39275eb9dcd6e1607d740cc7963f4616870761854990f24e710d10b77110ca9ff4ae6d2009b19afde0b23dc0dfcac4e2d3cb12f7748cd82a2cd89071961634f676d08a496b94106a8cf0c54859f57c7bb0e7a1fa03a309f3a79d80f41d81e4589fd9686;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h327fdeae343db7eda5f766642d6915266bb0d4ef847eae7b6a2636415830df0d5ed2b67b52180841a9e2b654336621324ee3b929f031c610af290a1ae8a6a4a6b65f34fc56f672be3f7f0ca4cdd689d663ba077b549a84b5cb2d417335ee96125500de702459cdfb38;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82ded6416053177e7e4a23c35c622d95264ffa4fad135fbbf9f5ffcf19390f04d4b43a0c728dc9d28da5f369fe9351892ca24953eaf87a2ffdf334ddfc3b464dad0c67e7295aca5a258780d37b903e488451781664c91a485894be87cd3ead5e3aebde08053b5c9a98;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130fcdc881349dd7c9b04b86c782257fe99e97222ef96e1c25a54faf2e7a565c1c90bb8aefcc535abceb2cb272b0aa40827a60653e008491f50ce4bb0ad4afd446eab02d71cc3b78a72ea1240282210b3b7faa0aba6872ab60de509010b8db78c77e4ae9f53353714e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc6c051704c9806e39e52a582c03242237c4afbb78e2501445adff174dfe00ef4502d3d48bf7b94e49413fe0214f59e7b992d64c23a57e736f8ab43fa4dcf7a5d25a252a89c9097f6abda18c296df0eb7c4999fc7157d2e2905d5680501c54baddf27391b73cdfc50f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aff4c5c01862bd7c380c8c40d69e325506010cf4f38ecb8356f8eb1c9ca0bb8f288a4c87df1ff027d5451129fe1a9fc96e03908f3fd2f4899c458fa7dc6bfd5b8374ce7d937f9987d96317533a2d96c8113a8ee2350b55717c8078d5324c945b726407bcc80f8a1492;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fddd341e3c04870e9e6febfe64e249fdbcb20eae213c6c642894072a4e6b77c92146378923719f7743c605fef8f37b12e956ce7d82a0398a18ddbe3d1377607e08e479f7f05795a8009685e2bc8f4dfd6abd5b81134bca8e1a096d5a16676acdea0c560349b46c1543;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146c840cf614b72df631f8cbba153b60c23efeeb1b99cb8c0ffcbb57d141ff8a5e50e283b0bdd60e6757968f243e6c15c6cd59edbb8b6e136808317389e2ee8f90b378fbb3dd061e7b9fda9b2d88c48b987373f2819bfffe9ab2286034f5861fdb8f84d65c332b538a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf3550cedf452a8272be67ea5697ee815989969cc77f099432ef6cefbf7acb590ab4bbc5f37770a98daff77fc037dd24e87b05e5abaa78efdf3317823ffd6763ad371b0a3a584cc5b248781c3ebaaec21385fe7061d4dc8462bce259e5b5c1e74a3ebb6b3ff69f14300;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd612a7bd2d85f8dd77c94e0bb7a8ee18a4ff50b765e70f74ca236bc071841c7e1e16214266c1161f9f3eef669112c8d3c598497ab6f6223321e7ae728526ec235b35ca5fc9d70c427c2308372d20c4af5fbfca08848af67822d1716fc7ce53b963e05e411d428e817;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f11506587cde51b04af227be4e6c061c30808213be70aaad0493be6a0f6dc7092e844f4ef0e63d54a9b49f6100decc34782b84414082b2e1a9873150d349e679f21df6e1b85398402d81395830bfc0df6cf226c2b8dd372069922d797511ad4cf921cf7a4e9063639;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h166d94ad73d56c0b9b12100eba93bf0348749d304a6d3707af66e52674314dde390f6fcb4e5715cdde2a96e2100490df70b618b065e4c606a870ceed376219f6998e3c3fc5317989198b8c81afcc8cf4c608e89501f4fda89233566548ffe6bd536f9d9bb240a9172be;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27d1abeb28105e496471b160f7baa1d6aba597b80c91a6d8c94d98d7ed376ada4576db76b1fb9abc4db97ec2bce9ae09d539487e800c285acd0c1d9db0d8d9fea59f70b2f4cf55fd8bed08f0d7ba335b0c6a7ca0f76eaacd542dbf619d0df74f849f4a2a8ac3f2915f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9964db4d7fa1c34d892cdc7e2eda7e41c517dfb075cdfd60ec04bd26232f752f75317311c3997760572d15a888c35d1f2473ce0a369b7af1afa58df7ba17da113aefbe25fa252d5147f9f31936fa4b2c7d6ee5bf8aa61a25de922595fa9d9e9d7181650fea318a4a92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1888091730e80861152bf3f56c975de464b80e1b32215e8c4d8e1b52bd3368721a7b10c939cdea060d208539db18800a5f72ab34c5f7904f1723f9f741311767699ecfa4ebb779b04c2751b466d9d9465353a9681f834a8d87c3dc0b4a2a77275243e1f45192578c3c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ff2a795aa47c9fa9aa6a542a041ab662d14ee09a60e805c862f7a54d484b984ab8755748175dae4806209b071f330fdc1565b575c8caf29522428473580b37c5942dba4acecb8aafa9e3c4940e6a087b69ddbb6bd0c5239ab9b63d73a7bbf5a3565fbe67bdb221c89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15755c272c0c1920166bfc6b65c4c0f82a574c688c043e1aa5589b024e097bab479ac624c3edf91f154d9c887f8468ef8dedcfcae4651cee68faeb556cb326bc396f748cfe63b207f012031275cb9acf2b5300d7bb529a3e7234b1b54e99823a62f8bc2b306d1c966cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56c6c9a2d4f73aa0dbe4ba940eca24e76018725caea33b96c7290924e43890f4750f8b8758be12826572e1819b95e6e288302657289624de835b7435c8aa8a2eae7b161ae992237d9a93f08361cb102edc1d4c0ecedb2ba679870ecacc7a49d0a66d453f78855dfacb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1324ce70c67cf2ff93596363312accdff46db6c71ea760b4242397760aaf04996f99fc69eb8f2583e948f1a6cc82c730b713f2e68ab800ca00b99463a4bccadada6df1899da7aaca0df0b2143a341dc1d752addefe8c67191fad83d22ab92ebc001e6ca7b7fc2e6c311;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hff9b35f2c7422c4f54bc2f977b999e1a1c68b1feffafb7d403544cb1e442c0fa97bb46cc87b2fea784894a861b46e256af01a3682e2b4937ba64a3ff252ab51c63dbf9b26b404d36fc0b463fb3f1e3c80eb8d0f561c9b8d85f8bb728561af09a83aa27f9b55ed0a62b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b7c4bb28ac11a042ad3213a81a3027239b1772edcd541409387dc20547148829419327b1e1d751b4066af5d64bfa8b00310282fd878fba46a897f20898bbc964ca76ff455e140b1f7aa8032f98d48027ae4870c6944c1039cf0ce60fba87fb28db5474af913221a2a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d391184e013eddc0e7e9468901876da68a30b8ced5fd3fa1b1de2cb5ecde69887b45b5b2c8641cbb16bc05c50563caf9ca56633c2635db58bacdb128b4728ea511b02fe9fe2c4129c3502c5f20507d8d68410b439eda13b6fc4a17c2ecb6fecc1699b1723bc376938;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da307a9e27adcb4a65a38f9b34f3711bdb47f0e9d95f12c7d0c52a9991830303b51c86d85759535448b2bed994c129a1537fcfd4e33f4fe2dbb3eebb6f303ee72f960126e53f412048904e2b4bdc8ec3ba353e7ad20826dc042df8f1c0fb0a0be635e951156620c9fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a809bd3ac7a266a6df1d496a3369236dcda627ecea04f9d0f4a6f81460c9058da9655de94a2fd160a56e8d57fe666d4b39cc7621deeb725d6fa3b15bc124a79234d4cc0d95df519182633b1e2bafcaa81e7232432da4aed7a8cfb21fd8194ccaef9005618dc0369ca3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h513a40d101e7e4c723a82a5e3e432071f23b241e6662250f138b29b4f2c10dbed6dec337c42dca87f89c76d60211d0613bc34afbe1dfda1b8b13c38911bc0d913b0a0e54b81fb0f0517f5db32e34a8507bc168d44ab44e25f7435bc186d71517b359845c2c1f28359c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h164966191346dabbfbf2f108a0f8037bc0f3a1fb00ff0214f6f4b9dda0689692321e45ad8d50c87df2fb3c7e5318229415e87ef93fe9906aa8e732b7d608553be5bf80f8544c8d8bbe5e1116328d1596f17ab05ff6d2aa681a1585ece957c2c9d975e884f00801e62b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15448d33ae7c79985616fad433e20fab8638b2156830d0e7c906e7c3c7a67436d27b986b4a60e6d79d88770c7049a478440b226a764d71d0672ded751f7a44ba71e61ebf2e78609e4f574224ea36cc24cf34f55dd1d6d46feadce540fce41ef77c8f470ebc3d84c9068;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h663badc354c5d3e3bf864031c35a7b42cc84e8a0e051de7aab8affc5244e44b8144ed73ff56e15615eae2addd8e33b1974f9306120302d8423db5b3a8165ddbca6822a5f62484fcfe24f445e0a9dfde97c9c2e4b645f206ba1d807570b682dedae4b5dd8ecfdac4f2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce7bb664059706579c24f136cbdd054c3d5c9fbd2c7ddb651a0a0f7bb3733f6d170a6807e40a774307790b5f780b5635b8e62435cfcf1f7e29b46d2f7e54680fbeb83d7963f8156a3ad573b465d7582dfac2d134b128921d055fca3fe640e853c4754875044e4d3958;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1085cffbb49d0313d2fe1979b3f2c79b981be38d67c8c59b41195d03e6ce29e5c16a66fe279c9ee21165daee59085d160e49226300a04790ab909dbc98fdb6464a1cf6b96c3952e8f9cd2d8d0ebfacb7fb0d8d8406ba4eabc7b0b7ab0170206a5de0956c37a5ec19df4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd02871be0c8d6ccef412d68b747ba7cc19723cec85845209d198f8850e50a49b77898464d01d2b06695e630d75919f4599787f965c8156eb8d8408687222ab490e08b22e53a644588df598043e4fee625e0655914b29895e5caae0f70ba90e81b6496ef5707196d077;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16301c6277ddfe64b615b2e5eea3d65bf067c4e3a409f3cfe6045a967515a94b43b47a5e9fa7281cb7def8f69ec6fb38e6624189873a3eb5d261c473b893c98f75eb08436aef54bfcab40ec78aaac12fec10c2f458928f78a83205be86f36c639ee9359ad5d98bcb533;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1baa6f536bee2b7d4b114704f77a7ae0e1306ae8724e885cb272b04c8dd4c8ab9ac74779d1bd90e07a422b790705d533e5341b341b4d08890ac482dde6b627728bb63786b7b1ddd173f65e3de687ed4dea49732670d90f53adef391fec69ef73b2ddb6b6da87d068811;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163de422fbe871a6f366d73cd098a519940752a91b7dc339d8a0f45acaf46fbfcfc1df3ac33a731882dd8fa1ee796a10de6c85b6dbb41b4c87b003e8b42031837aabf99d12de05ccbfda746877665a8559293568417be7cd44f2eb65b802cdddb3a76410a709d2880ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1baf5b149e3316ea6e5735a31a7b210e383f55fe6019c2682ec868de15d6586dc2d18f315fd03e9d66f86140551c94e2954f86992e07cda97b326f0d7eddce48866a99ec02090aa1ffbea4f546a578bfe255092b102a9c10be13676b21b5a2cba7c7445352b165accd4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f76d9a5981c4ee1c38cd7dba1bc93b2e7ee140febb2299326dc32cf2923cd31f9fe2770b48fdfdf2748d4f69d9948f603e6c3396f499ce965b3cebd3454c0d3302f153bbc1cec22391e1e6fdfcf3523ec834adfba088a3327683462aee39488ad23932d9c446c9fa14;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h162fb519bf8845a828d44c435a4b7118cae2ab3af6e3cfb452813fef3c5f0408a4761f81a7b2e0d30c78bac9d80478c6545a09d1a7d815993fda288924993cc92ba346f79bbfb3d3c5baf041d6eead5c4ac0c62a3ddc838b833eb810e65b3f8fad920840d37fd1204cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he64e3064e8bfa1ee7c9495f20cf8165e34b0640cbd765d85226c35a93697ac13ba4337bc66e0aa8d6db5cec51d64dd722b0e00d99ff4c3d30c3e3036c0b2004cb645c63f7b3f6b624b8ef465ef59520db39fcb2095169147588a1ada1a79714134a7c1877e135138a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19960f97925a184ad7e47c9ccb1f129292e36e57ca7271a1bf6512d9752e502feeec8d4510b765532d49eed5ce6ef12c6f5c2797b46d96fde365b8abd91be6096e2d05baa969207a570dd9ca4e281f6355957da76b9e42bd4dcf72b0542eacdfb9615737f61e46e6f27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h23d6123ef0a208b55cbf7ac95173e20aa7024e77b6c516b232f5ee81c4195b0adc486afab47415c8c7d96006b49dd9327c96f75b743dc88606061df71d971311a5be952831da083ec42cce55e1d251768b5b164a04351b889241c8888fa304c22d22bcc0af2434f8a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123f071ded277dfa3b5206cc5d4bc1fa2e4fc4c09b5d6153d0bb3abab364dc2923781f985aafe240e29102da453180861763a663af54e801d33fd057ae47b301b66a76ba29d9c5aa4d7b7c3ba738faa923f75b91105d36f46beaf53ea8d83660194e35a8927a43463fc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1360fc148c76832e013baf3a79507302eef6f1c31d7940942ec0bdcab89a6db0e2d238ef2e58da29c3a3cf6a4bb8dd80a9ade70c9fecb0f64ba6e1b4999a09c61b178c067853e469687f85be9b9b3f2ad12a9feb4cbb44cd165f58d70e50a7411bfae193a4e76e04fb5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13604e0e1e0b58850ae4d91228b2e0447de472e6af2960bdf4ce9a9dbfeea03a7cedae84cee2eebbf3f208ed062fa656953f9693361a38eb28dd3ccb61844162f554ea45191f82b669150d81b306668b3cb55b9bc395e9313e6be8a9350ebc47c8772094380037e8c99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha61a00ed2f26987ff1d019155775b9effabb088500109d1379dcab8e7e31c1c234955683cebfce77dde246494a64fe10e537e58e27b3cf565f7777dd8003968e0f2f2700049ee3ba9bce1448f3366463037dfdf288ac80cfe116bb922a066e68a92d46281a78ad92aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1607486dbf254f7bacd15c5f1017853f52eb9eaf04d0c22a6c82bc0f964fe7fb56319030184a7fefa60557e436c6d05fcd6e14c3e52332f23b4ea640e1f44b8f8d1de066ef0b5f245242d1be4488c0095e63ae959cd8f3dc96ed33c7b459c9ce9f150e0773bc5604263;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8fe7b87178e406fe011fe26403f467e1bc73bc06e1bd49c673d95c7357480fa089557fc39792ef0c5a4eb0299b62902607825189b8c9782d95d595c17b0c35b5cc87c22be4abb108c6fbfbe2d7e8874d39c05022b644430f37bd4df49c69d42f1ed908e1d6d75b01a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165188f9db1991174f19b15e29f03b091c57182da58865801526af50f8dc5cbe1b0fd55b664faa5605da676e49a2ec9a22b7118f95bdae4aa359fa63dd0c372746b577a7079675042c1bf42df2cc9a7f5e6e84f235ebeff953c5ccc5148a6d8c4ed9809f7c27dd7437a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbff9c98b944e5cb0346754972f58bdd48584940dd071abd9e57cb179f1f711305f75507d837debe0b44fab02179cf024fbe25cb221ae73039afff3bbdb5b131d36bde7eecca1d337fc476c1f3c606898b5fac9675443d7dc1f02d52e3f78761d4ea38d8174a54d3261;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da1dab42be42e59e29cdaeb536c4865003770ec5245e8b8ff37926e2511c18579d9f1f511118deeb154beb60e461e77803c08a162bbf8bd92f533f48f3e3e454747d9762e1a9405e771f69ccefbfd4ee152e1e4f4dd57892301d2b3fa8f418154b81968efde562a1d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4be33af02dc0341de224ec71e8081376a12241e2f48e8e473b90d1cfbf11eb6a341b01dd45dc89b40c6099700aaa3467b5bcaf5d8cb8715677527053793bfddf687bfbc23475ee9abd33b94718971b0c7946544c26bd87ea42d08c273026e2bc1f94569dc72ddb9f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha1fa056f9718f2433eea8db8891fdd193219c5d107317a164fbecb00c5b29f52c59365e3c9cda161516736b128d85ac1a9967ea0cd709bc7c59bd8fd6af749f576307c30a34139cc7d52b66384c9fe73848ff69c658fdb38cffeec43c9567995d4fe34371bf7cd9d68;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2545ac8fd5ad428535abbb84b1e1d7878b19ad217b4d62479c43b9ec1183ff759a859522c6d25643620dda6f8a9275b426bb632811687e74c32f0e36e639ccfa7de4062fdf515edefde96ce7551a595a410fb18d0e486b9add36e29949ecbc65d40cc768a8428c1449;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h48d386599e51c4c2abbdc031ad8dcd81eb0b624c8bc503a663d915baadd9649ca7c39c2498939ff3f1e0950fc8c7dabcd3a5f43cec2706a4d9a2a50f20cf483c93e4ae2069e198b1a64b1c7a30a79c03a9a44d2c5efc5658fb1630f42f1123adcdaa51978296e983a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc4f2469ddc0ccf36d5e1929f759cf9b7e5c1aa1c6498ea11d0c72b6dc7fe02fafe7731804c294c95fca10db0393d98b67aab218e79198c769a1624b015d2be2da480b8dd9410e3216875398dcf381ab122c876b154ada58bfa503342f60f93ead002646af6e71a76cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6364932713f630bd388c5a8d2f260da1f40232e0bcb34b10f99c810624900115d26a958ae2db88747c466a925e5326b04f40ba9a3b9097ef704ef9d9d769fa72f40f85c129f648108128f9884fe8a126eec2cf3e47062e3ed610f8a144a63cfb52ec82c3a44daaba24;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81c51ad39bb52fb601c96cea21da11ad121991c03e6e706567615c333f1a5a6ee3ec8df78a1e566eea75e382a17e690f54961595c8b1bb7d9a620686c9bd6e995dab0fa41d955626bd1d6e9d211eca95845409b5f3b1f1c75df81f89974e1cac6e10bccebace6da39a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d8ee4b2b64536d28e12f0593258961edfb30ccabf9c807a5e95e66faba7b4bbb7ca3d04b049a89d9ce378afbf70a5eecc29b3f012b8d0f7d13cc9f019e8f5c6e51f80ae269c395fd5cca9e1c1d2ee61524dc3747819d2d0fcace9135bc01429fcf43a5b92a3d14d4e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5d2536eeafe04c1d6e462aeb8fa85a408f4d26318cce7e26f47565f7d4577d55b6e131e12c5402a89bb8d49737770a04a63bdf6ba31f8107c72bc016937b7e959fdd944c611aba69e1991fea461426ae70d6090a46dc8fd2db352593516d4ca169359acb09c3d5d7b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h554ad998db3bf613513e09e8e99e3a65bbbf532a15ce87e32c5a44146a6a8473661369bc27d1a1012a4e1390572a73b619f5d0ef837cf88927b2973356ca5e552281672e68fd0a5e2248f9da98fcd6b5f4419e1971830ae50a992dfbe2d090cb87b8ced3f030159841;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd9befb87043cbd587037b185d6eb17ed14884f23dcad4f8901a361f05454bb036472c5be5cc6bc53868ef2550b70c9f4873cab4f4c81a621dc5a03868bc26890c1615b357cbaef5183a802a5e86b60c135a5c7756637f153a2289ff0a0eb39ac66a511d5d9f021d49a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h189238d1652ba2eb8cf7e33a374164fe03dec0d70f2f0a16b15e756c0837904d89031fd170e47d8fbfebc8a2f70ed0ea484d0438de43f98b0860c55a6a3907a352d3707a1fadee117264c8ce0b227a33a78aa29dd2c216e19a71dd16c289a2383ff79abf0f115f90f39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d48c788321ad80f642591bbae13c35067307b0bbee57b4b1d29e401c5b17bae613b1da28e29a6749f798837f63b80f4435b53ad818eb746a20a592934db4c85e1200b8fe3456ff7c826b3af6871a27521d17862aab816be7eb7525cb30b29642c0de4dea3dda72e13;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17df77ff7cb4053f2d5c167dd9a8cc5a8203e07fe79cb6cb8f603b6ab4dc407fa510e7ea0877ca56642f7838e967be8aab8f3cb2175754359f5decc3a8b242eef5a4c5c9c8f1d50f9bc457f230d01cf184e610366a5ce4e9b7e623258cf7a59b9fc8dcfd1baa5f628b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7385e70059fb66e09d58ae74ec6fbf77e5504d8b7a50594bc42efe06466349c72f34ef4eadcaa08de93fb592d3059f9b982a4541be7129f8cc1fbf096a14826685ce0576308214cecc1fc2d651019e3c8ba34b75747f1ab41610b0420953e98c0b9312398e45931746;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28f5bcc889f7361282079a00b98afc587e9369bdf727407d810487f17dde067426a371b0fc8c52eb67cd6bdce8e0c889d460f95d172c00bd9d7c849c3335aa29afaf36ac70aeeec74f2f3b7c05c4e1334ae725bb77acf86f985ab43fadd312cd32a3eba12fcaebbd98;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18c68e5f2c31ceafd6efb340ead66ffd04c46706d1ba3911b92f9d54db3b69321b56b90b8cf1b5039bb9bd36380282145f6dcf3792bf616bab64a5ba606b93fd855b82a63a62774dbf7f779a213ff08cb8ce694cfa29ef31bd9fad1f7185d3cc0f21684f481285ac0b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16409ec7f3d6becaaeb2f19766867d8df35a36cb6ae31fb9f7ad263bac63f69fa5c80dc1653a455127428f2c5d8552b5a2ad3b37b1c352e8f95bde337627100dee1e87b4d4d9fb2364f39644ebae63e96fa4ca4fcfbb4c9bf11bb9ac5fce0622c5e089fcf4d0be8b3c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h196d4c74e80a9f5dff2024c813abc57de5feefd2f81a07d812850ae8fbc10b0c38b2a1c787b2cc356cc823673790918de6ec86717da23e0102a571d3704e2775d2b752eb6c6b962c2c3930de3fdf7f402723d58e9ad139c0e5198ec3ad9fe919a01f6cbc6cf1fb51aa8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e54412b9d54c4887a3bbf04db20409e51f20e7ad3080d630fd32b02e74b8509e8b6d13595a6e741714417440fbcf2241dd8b8c88b808b8f2f470975dea318697e8ebeaaf92365d34ad486f5874de3a79abbcc4bfb5eaf75d27d1c70a4fcd1253eba8c7f62c5dfa2a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd69bb4895d097a1ea259af906097c5a538432191c6917b34200517d85e380976f09b0da5c90b6742f8bb10857679f4463158cf61679faa787aff2403118c0410997e9389c65da9349b585cb79ebec8e3c380d571311a5947eb127e8afde0b04d694cacf94a0cb2f9d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f13058f273b37a47691238deb06527d7b1c838d595cc20d151955a73972d015a11f5a2b373fbf44088b1c682b6487db8c50ebc34df13a13d9078216ebbff190891681332ecc480eeee058f84d53aa434fe3b245a191b12ac3d54701ce7f82101b74abed74b618802b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61a1e94ef3fd452f5d8888d0ca93c5569bf15ba55cf57435eab2139e040958fb9d827e45e940da5bdce939970e84b50a5a127cfabe2a21259dc619051abeac0bf1bae0452ee7b3e614e63aab945449dbe6a80bc99f5ebf16e737d15105b5799716dc8b95da770b21e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf905e2d2bec181045fb44e3f24f58a217ae42a01ad7eacc6576813b857fdc35705e23c9c487a915028f60dac41ad89c9966430edcca1f0d1b276917e9df30e10011050939bc9a496f1ffdc3ebdc22ad62b74d6fec84ef5d4df2daced286ebf92092f5406b757c816a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdab18e378dc4dc607106597cc34bcf25375795d8103a8a45eaa5dc25c21505866bb607026ab6f761dd212af915dfd7a011dc8fc57b7d0bbfeb4c06aa0e5a1947811b50f64716fc41291aa7c3115b0201a6b7fc5e6dbb3d7a02b90a8270afb8487f2140868254189b4a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a8128b808b3038b2ab354c2212f27d60b6462b7a2e9d71199b6ee30f72589247e70e8652b4d87117f8e6c44c1f439736a5d64effac65221bfcb6815a1c7f45a6d4ea9cd2e4d06af31d1673f3b5aa3001afecc9f670948ca9ae1a0adf3dcc5bcaf50f1004be0146e56;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hef96848e7a2e596b4780052d791c70daf8af5d593d4b65ccb2cf599885bb19823de0fc8c27a18fc96f94bd8fbfa1f84c4c6e0feea0b37ac2b591d70a85634f204b58b49d5caced11cd4c94e2a4dbd9a54d6ef766f3a51bef1b7131c5b00f573b4abf3adc5d6fc2f89e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5e0168779e6eae4902dd4be5cfe1e37f22cc486f3806dcc68683c6dc07d501f1eab0fc6792d177310e79b8d1be249d38fe1a00baac55d0b3f21c3c80bb2b743b00733b1feecc898922b98e5e59822d75c6305c05e29340de76616866881b2c02af956c9639f68e3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h198b23013a526748031fc5c940f264706ba1301f5403e59b20a62186d29ed853c9cd60b529058ff469fb5b9fd640bbd090c92512c936382cad9ec4bf987e929aa924b54cbdd8b7c9c169b5abc53564da364164b9c403ea2b91f489bc8a7707a0819d2c09d397462df99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f1e927e48c62b6883079d1410bd9310ee182fc0b4cb265a3caa3116beafaea6f6270aa0f39bc0a8747b595733f53c9721c0de7024e805ecbfa9adf0b2f5aea0fecbf1db1aaf63fd661b76475980b193ae76e83e298a4daa5b44dd1ba51a3420bcd2066bfb0878465c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h156614a8672df267f646192932c9419842a695ecfc1318727b80593b3bcaeb8230e52979fff81e8dfd6b76d3a546cccfdd3a187cae20d52fe7af1745f7a0ec29929121af550ffa4eb5e0111c3ff2defdacb64e882307e1c0449d3c4c46e879f332bbe8d5ce2cbf8e1c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14207384bf78b2b3dcb543710a1526b6098017474f8428cf6680072462b8b4ac42e8ad89a2a59c1421c5bf76d7ecb6decc10611c6793bfd43c70ed46c29165e9f3b2463510b55cb323cae7bd7443dd3142c82abd9f93185734810ee5a65c0920070e6a84fcfc2fd5954;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123df37b51f166d994f54cdbd4ca95c1fc58a05fd106744f32316098ac9f3d3736817fffc8c8ed7fe7b0f4b259453a152ddd2696116de844573516ddb6ddea978026e6b2ffb0d9f555d7e0dbefaf84cd13d5cf163bb81b085bde9773e5ae576f798450423b6ec1109f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b98ceecd91e5e154b1896bb4e234b2d15bad647229df04b2a6326f5939fe68ad8a4ef4c9236c15ad3f084d6c3331b1bcabf1db48cee0ecdf24f491f6d03cf4dde488d6ee8934447545e72c1980cc550d3303ea0102c6cb71149c79ed77899f5fe6c6c8b3ea3a4ed19;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h120f4af1657c89419e8cb52bf9421600fb65abd21d3be15071c20dc4d731aa64a449dcb8253dcedf06fe91096686c05510e53556daa44af9e84c80107a8871f7a8afd56b953915f956c59ffa9a42db5c59bbbec49b770e7de8908a3249329e90ffbb337c76ccbd12a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e649bc0202b30c1211efcdbf9b8a2d8a1bc5d3f19ee3f0929a47af2a51e03227621b1552681613fa4b750fc949b860233b79e8c5f6247aee70e4eff265f29c58a6a8124a7923e31bb10814e88c8f198d3302ec36c08b32a4f17416aa5451cb3190a8a8db5ee251402;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb70dc23480fe164e0fcf7af65bc7e7e67f924ff9ab798e7a8727e5d931e01a900435ecd40aeb597266b5ae93697344866738f1df41cfeb513dd9cd2e08ca7e1c671978a0926eaea9d9bfc7392f15e52355ad9c5ea9e3b95299e5c835dc40f785b718d830068770730b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167e8e51379e71b025d6d85f5fc36841a0cfe30ae357ccfc6a547d688083babe45a3cd04b383c55d3849e4ab7db7edf287a371c35fb48daae6ae2193e89fbbdd5d255e5a976727f039ba28afc9f8d2e19725b3306d77b0a4bb47621181906fde9382df0934ccc07c7be;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2248f3c4cb2d7e07202b80f88bb23ac4630db6e5e5100b9200dc68bffe8005a4c69dab0e91bbfc2be0301b8efa8d12a6114ea7f918bcfde4a92ce1873ce30a07234147644a88436d2518e2d77bfad7b45b777da5178fde7c7eb0abeb38e05dec363f7485048e7fca73;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132c8574dfc518dd3f6fcaa99cf7ffacb5d7e186fd944a6eeba95bbce902d6c5a994df91d27d23b8ec51467a2a317afb5f2c6b741504eaca7de5d3ac9c9aab0a6415bec11a6d4deb56b597be9b378cec7e4ac2228aadd1c5952d84309ebe400b2b7cff2058673061c1e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d2be03e1907b254a2f3538d64fcedc25c0b1260c60094e4fbe9aa168b3d308e64b6a93ab7fbbd21f645d25ca829cffe5a8f2b2966a65e18c2a21bd77e1477953040a3673fa9321d5b8110d8ce1d3cc4220dd8c94073a0bc9d9b2a2c1322c35e770bef126fd28e223c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1013991601e253f4826275a8383055f3095db2be103fb9ed735354a71efd264b1d4489a0cda86ad22a53ae6b6202a9d821441fac39c6f7059eab590691a28e87ef54bfa347aeca9ee240621ed9956abda6bbb7496ab371bdb813b9cf88be0490be4db8f9542a9c56549;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8d7739a57c07f79b83dddf695f5a5c10452a6d8bedb35fa4c319d30d639facb09c4b155cd96d260ed2846bee1446539734eb69c617f0d917a1ad98f32c1bda8c6462be96ebd020e0b2e6982fbc7a411d763f75cd9d11c9c68c45928cf3f344ad51d6653f73e593335;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2bc7000674503f1506ba1761235fb883b586e746a54210952c509ed8b6c7c4a961a547d51c8b500756d9f3514ea0f33ecbda7d1d7dffb381e1cae1c9fd3be0abba6a6f54deeb43754d45ecba34313bdd603725733293a6362f9602f1f3007f2ca6db3af42e83c38112;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16f53660561fecf11e5af4ee684ebb61f49c34f2c8a5a3b4118e62f0952d5aa3226f72e4a032737d350c9feda6c6a1d8d27e3365bd5f30bbe6dd3a4bbba5e06541954dfb6df3e8edf820b8d15fd17ec7294fbc4d4097161e3f61b78549f7efa5930c1e5edb9388b17ce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a13d790a410271666b6fd33f53bac24d8a1f8397efbef254a7ca1c8380a6691e7d773118ad615644d2ff1e33a77d1003f83c71b9f105fa0c2001b66e78d86decae9b1ddae66233eb145911ddf568f09750a15bd7ed0c1bf7efc36b546b72de797c561a74a3fb5f92c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf200f7b16f370da3879e9c490875b540db2db52710cf9f44da5e429458e4070153a5244071c53ae5512332a9ea69df6cdbe7b7943f71a663faf7adb99e1ec3ef996109f80fbc30f924eba94c493d5c9a38918d8cf60f306b13528869ee005927e39cfa6d553c398e10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17367fe70ab8db4738b8f4bc1119c90b9fbdd0bb31deb0c4eb4bb564a24d1f4b8853a3c3248178d88b84c6ae8490e5bc4175fcf48506c9e20e73dd81057c5004743133aa1041543a8b28a3a660ffecd5ccbc12c998e1d09b997780da4c05331f1957b1f22380541687f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ee1dcf515896f66826a59e5ff260dda8fdcccb0cb3f2e2a2b750fe1fe08f8e7071c0f9c2c4e0776f46153a00722b36c7d67202142a0c093e681d7f030d1e8ac4a95b9303f0e7041c60c95527402a20544bdb4d4996feaffa3e65845834ac2a9b3cf48aa6b76794056;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118b6666cd236b7dad614f50e99a4846177131f92c03ca35532cbd66eb8678cc5f37557dd93df34f88a5ec965cf5d51bd8a2496322aea8d5fd1caa56732cdd0b5a633c24bd6aa10fc37a9de3e43270c61e5e75f898c64ee3cd9d2a0de44bf7208d3daf6193db1ce339b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bdffb40668d2138ba2e14ca1bfe9742067fc9e4cf80bfa9a2c81c159185d138ba3bff5513b1b8e512fcb23fe0f40a943ffdbb1a62fd0e73de1871248ca39c5552127c10c039e915fa690ba71c7f7bebdc730936f949e427c37bba85de43a33bd4b39748011f8061c34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42bfef44ad8507a6a0f12abf0c04105dc0c8fed4909ed7708a2db2d85cd3a35a8b0a22a16e3d36b4cf8339b32794fba62229bf7af6ac669603a8dfac11ffa0e43c97fe7d6c88a5dd54b60c20bc31f6994b36f7e2010207adf1f51ae9cb676f9068cecf4ca502cd9ea3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4a1884f64c443191f9100439dacd3a288ac850021fc8f2f4ce4cd44c1ba5361f53bbad0230ab173392feb8f7a6f6f614aa0d917f65f3f837be5e16d48003de91a9816f516e8593583c8b78f9302acdfbe8b5aa0e3c1c02b1272fea3e2799dff230f879d27117fd4c04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5cf78ddd0f3724811e3c53b2c03ebfb474e5ca37df5c140842ae659b0f8431d8dd01e3d7035cab8e74c500b19c8a547a4aeeaba76feb329f33642d700dd3d98c7a3ff26428cbd74f0730274f78108cc565d20b704742f6e80f7fa531a0af96db738d5c9dd70e34450a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85e7268ac6364c8372232206ee016049b2f37bdd03c780cc8f9cf74a330c968e7a1fdfc45d1327beb613e5adf8f094c69e8f4d71f17ec0d7507645e9ec6854f1e2e78ad22fac43f6dfaa99f2f1148f10b373610d319bab5a43d586d599ace75c42ad97c395b4c1ad85;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17de4163bac8c3f7e498469bd1bc5e8ef1fe81f9fbd4e7e861485545e81202d9aec618635770922c8813eec1feaf39896fedbbdb95e51eb344ef6f268a713b4c0aed4fdaf47ae630d6e1351f1666cadaa45a38c4dfcd146f972f2386387f092fa36814fdf39217a575a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a923b0fdd69705d6a1343bc96a3fd02554424e4930f0fe7c51eb848df09a81df19988ecf5516f5c5890ca994b3e726668e1252fc38bc57ee13979719399c3290ef8c21707517fbba5e120dbd1481c76f4cc20284c284822594d6454dbb7b48620c1d39019f734262c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h109f2293eb02fdc86734ee0cc00eb9d7509ab9b7f7faf07912df845cc2cb9a47c05cd2820e21f81cb09d306e994137638f53ac9029083dd46af6151b46348b602f479e2c9e0bd28827f519390a3348d48def7b384a6d801edb576de9ce0c56616c8ac7ec6df61d4f0f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8cea72738e8c8e4432f2704166b76ec473bca40d2a24152de5660146cff018132fa43950704b687114a3eddeae1b3353e1eb424e2747cfb0d816d790ef0e3792c2e531cf7af7d03b4b8f0a2eec2a0765a04a82b586e94271a0638e3dba670823f4b3e919268af923b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc05a207e5594e974d3b90b4f60eea755fb58ba93a23bc328733f05bc21736d45927c904a0b023d48867fa285d4755c353d345fafb22b3cde52e94949f7cf72c04e5f1f3a99a6a637c0ffd0dab6179b81ab333e3c0b7c85f4d16f6eaf512dbb3b084e3e9d5416c47ce5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f187298ec73251c9e080c0091e8aebd82613c277dcb8e07aed989ca7e71e15ba753e979b4acae38fd0853282674cd2fdae3f34c77c318012421a0a0402964a762e6445c3d676f7633cb8719ab30c8f4caf6be12d72f93161805b8e23643267ffb0681813b58e7d847;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb1ea8b45ccc90eb7f15d436d25316273c73a721f85a5e7b45f936763d8e8f72b63c3a4b2ad4decdc765c479d3478a8bfe97773b9daedbc51552a70fdb6d924cae61c713794c48e0eb3cbc93d473b184e5aeab4013ae72561f42fe6ff799acbf21c07acb2eda429df3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174e0b5a5f41236e7cc2dc739c4a924173e9454dfc1a658a7d03964cab0e78638885e7acc8407a7a6190e62aaa75895e0353b74be8e25ecdd141911804b8d5dced6658c6afa36730630c1f5f43bb39ef5a17042c33500ee6963c013183c13004e96f1d25ed5c7f871f8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1257322e5696081d501beed0fcb277aaa461eb07620b7306f7957f2d5ef0de7046df671ca75e85a0c423e384d3384913606640a81ddc34a1aeb420a5cdefa59e3495b8e2703b4cb3df017888684decf9289a75604a76e6714b9453f8cca75096a26f68aabe505daee26;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd07c9cb229e1c485ab230892f706ede6132a9696416756fe34e54c1e359f4e0a45c6a554909ddf7cf01030101224f79035cd2a60a109c8e818b1f05e879756ab106b702a857866d7011d070392d823ef96a8ac9b00b3f813ee359dc5685df4b1eedc58c59f0145f698;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb4285cc6efe44f28f0b5fd77a1d1a97f411df92da6f6323f038becbb6cddec54e2d190f0d76ed5921350066ff91bca124e8806921b32f7b2c16e1b0539f5df2ec7aa966e979552fd9407c036b8d0d46a1fc08453c0d6e77c82af29275b877438e72fe4a65a6cdb7b49;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e14f1c4c4a9530e2e47e30cd72c82608e4727581ed71d7dacf37b34c2f432b16b41186cd0b434dc6a58e0c6f14f6309c1c37f0b5de90a333cd3fb322f41d6c64917b6944c1838acf98008f7dcd276f711e6c2342629c96d4f7cd150a32029f2ea20c1a81fb8f367e1b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17db42bef2354a37b45c48e61d3ac03d1c907d0c61a6e5d6f937e6973c7b8853214c1f075bc10bd71da9ac9e11854446be5543422a5d31b854921ae67d8aec044696fd816297a4444a8abf99ae06465c0ff88cacf1376154fc6be9ca06cc5f054c31140792a48d4cd7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17166d5c1a2ceac5f8f1f8dd1450257fd90d691429114257e6361474e1d69bcc0c2486e4b347cf442c35a7f3e01e9651dc329d0779136f9b6f7be9554a65d69ec6467f1685e80107130c74c51e0ec611b0fa2ff9cc1df7e1826c00c1b806f5e7698f54bb941331870c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a298475d975317d0ae3ddb9dc624d017df6b50352bf10293e792f26badd0df71629ec71ac15068600e8908f2104e43bcb4f8be7d9f7046c26185a75f624a6aefec5a7177d971a962313d98d18719f70bb77c4e4a605b58873c34db23b364a8060142adb42f8d6d4a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6b6d8e1189a4696115c5fa8c5b36a510fc5e49de909341cb2b10e9b6fa24dc1f5096aea119535e2f5fc6a8ebd1126409b24ec7ac94da8d49629458c3f42c4910be2c14e8eb063f68b71b24dbdc4814b381ce60db1dc8f8e2dcc67bab6db5f015c40f754185d5d0262;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dabfa1a0bc2a233e3f15780dabfc84a0c5c9e10c34562dbf087158ea8a017059e79acee371d3fc21002e75c1a0624520476b8b590b7358011bfffc1e8100ec17c0d08e6e1421dd7f9a68be511e8d01fffd26c3ec5e0c7b055bd9dc587a6619cda6bbcdb8fe1023e3e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38a40aa0d0417e5c3b7da7e7125db38e74fd88d6de2845e3f2820c798b226aa892ac0ded9fe4440d49db682f05a729c13113bc08da80edc3ec725912ebda5a7f704702dee824344e807541192632d73cedc0cce2874a63c3eebbbffbc6febef868f2196dd74e7e329c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18457db09584bcf39264cb10c643e5f2dcedd839aa6a4b6fe5dd8bc388689256d9a25cdaf62058acf947b844cb31bd5401b9bccaf852f532c919ef21eeaae429cb6c82ed9f8e28ceed84346b4c940057a0e588030ea020f5a32b5c57e427a742c26f089287076a9951e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1345943632073159279c7055829110c25ba675d07273cdbf5c48d413a24c71002ef46a48ce82a9bc81680947aed970889f1bf6cac2d609e6bf2d4b4fc5eda3bca3097f846bd05946bb657df550b6e96d7835b91b9681f32ccbe5afbc3f803ee58fe87225edbe1e7f541;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b912f7768e616056c6bdbde2891c3a7d44f7fd8a3f70bcdf5a08a27feb45e2981f031cb1c4628747e49bf27c9d5a450e44b1272be47fe173cd8cf4c2716ec4cc26e75f4b9824c8bcfa51941c1be6994f0d0e717121c909406eafa7c200e8c0b26011170db966ca274;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85f0c90c5540330c38056af873693cd574a5e06f9e477520d35e6e54946f2e66a17a1253d7df81e49c33651e111c7e5deb5569b12721b90060d908c75b947c5eb3b1ecc5b923a877984e065e3ecd3326b82ab08882d2b305d26ae62aa87be20a885097213988864cd5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1c67c5c9dd1688fc1d83f5fadd414923d9f9f8d7ec9a5f2709d4c1f607eb4b8eb12ba43dddd034fff3787600ecabf7eeec758c783a27c34203a64908eede87d0593dae1896ccc1c7b8c2279945a8b1c63c419525b9d546d703de33a1f6e365e1f122b2a3a3222a345;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19f1a84ea4883f265032649ef95986d59a2b72ba08ad98e20c48bb0e9ee04da874c22a152b560ddcf1173211fb091b56d2655c5660ed104e9e8017fcd0f50b745f8a0cb392dfbd2e24cf524e55f629a2fb1735c5012e7c16d284695ce5eb19d64d82fff7b8e1bb9d843;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca9b50294315c2f55c5df54cb39e63fd7028281705f9a5ae54a61f99fd14b606b8d3edf4b9a1bd3583bf060bfa8513c0dd990a739008f9d456b217cea30c047e88dfe100a9e3f338acd2d15ea57b82b630a7da92fbf6bd364d9d2d23d603dc9d683ea1b7aebeaecb05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h117c2effc877115c31e94838c81454f4f30687c9e41f764af9755fe25b85554a50d7e53ccd997c3c9b560638bee32915f5e3d5ea18832464deb125546743b8b50da284ea00275a33bc374be5eb58c62fcb04aa5f7fee5066a20e76494bd4b979b6952d925fb0bf24188;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2dded74b517389741534a92fa92cbd563ffdd0a35832aa915d1075952750ad28b65b1118fa57ad7d28ac6ea7bbf61406fccc6bf37061ab6eeb406432e8e82d41113f61e061c1e0db90b7b4d774d6f229dd2053cf2d23726aa2d5deecd651043ee070309db8720d36b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e768ebd3fc22839b6bd81a1d68c65fce4226d2f298934f60b8e99f9b22cccff8aff5a80184e5f7cbe264e57caef061c6a6c5c3e38f2c7638d20daa9058b50fd382a0a71f2ac7ac0a38c221ef5fb64ee5ef151c1a1a9e81a0362db777fc75108e47e6bdb7a595e1b1e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eb96e054340132e60db103846a1b5060b2d8be1a895dc1c425712689f6df1cae486c2f6e6c05d75ea6f4923bdeba647ee4180dea7fcf52f4c606a3c3f20fd04d95e5297566879ebe68e308ac0d5c7668b7141388575f2c6de1233a34be9034038f3c244afffb6fc00b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h893bc9adb1b26cec21c715e09c853a5bd1332d2ac067b9a70951762003a22d7f3346073d23d6ff4715a6dc07eb7eaf969b77245f1a22d9d3722a9cb965670e7aef732cf4d76c13e5bd5a771ef762b067f6a92648789471044e6cf6654137b804bf93f0b6d7666e97a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab8d6fa3b86ebb49423b21a12612de4408d785f0faed31bd54de17da3dd77ec78dde6393a7112bc86698bd63d45e2a7a7f9d931a56bf4869ed3af52431f9d4052024fdc4afdb146c5a3e25801d6bdf7ed1a598e81d88bd31962963fcc4f26adbff7f0881c315d8c80b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179eb515e815c3bf3c05a550e40f5dbddc0c2efdc23a0421ea63f61d87b1bc82384eefcf1cdfb5ee7e449cc35b4006a5f678f316b4a1dce96a0080e90529c495445c21943d7c205affadab2c4f51ef9024e4daed79d6e8d416b04bb14b6cf9d3e238687deb9ec0ea5cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78c7678eef6893d48af5e038aec1d3186bb7e1e6e583eb679eda43e441d7adcd25ff4b8648d008211c4412c6c21e6c02dada6363553aee6d1032602caa37abb86b2fbb146f53637f602080ee5bebf6de0e81a66016029fc296070db1e59775413aa8ed41469f9b234d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ce1a050877b9ae396c887ad66ef5bb84c971747cf83f5b0c1186064fccd9f5453bbb5c586a6f52d98294bc43158e21b1cb9e3288f843e85cc22795ee8fb1a9ff19596e18704ec33bf2ee04dd9d1fa89b0893660584f989ef130b3e95e3e7f735374f780afe5e44e28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2d30185dc97f4d86781d34d8a70e932a76f74302151b12242de6900747517dd0f7cfcb08f1a76c3f68dfe68ab3e1aadd94fe07ef981dd5e72c0e2f5a78311afbf2fb8f40478a2e3ed3e7c28d5db462e5a52243372fe7a9a23c6222814b8955ef473758fea3d6ca210;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17866af2342f374421a4a5f49bad62d6548279ecb323f3c775aa0bdae40e20d9d835c14474a4902a5dcd5716a0c50385dd09e55291c81bfabb6ebb94426bd5b8400e8a47ef5a1b3c14459f1a539b7c7ece2a0a3fbf56d487f5bad1e1e687426df6b1069e1caf46ffc9d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47f7c8f260a7951872fffeb73edef214cb97a3d9741f40769e8007ac1e5fb4f4b3f67e49adb7f6c22f8d88f5a2d81bc7364ad64ce7a0839ea2bde72e4ff687313356353720c434ac7c5ce5b66cd5784eb70cf0ecc659d9d839d1a9312d457c3e3ce7497f9c886bb1e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he109a8f089f86da9fd293024446881f1be5cd15acb4b75f7c2b1a5f82107445493cddefcde83173144ede5a49384d8d16bce892ede92bf375552808433bc53ea7e83e1139019f63e8880ef370111de49962e6fa66df0245056dc18ad9a993f6068ddb1a70aae1c455d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d4af6f62055da090f119bbc2485012af4e5e0be9c3d29230fa5eda8a408249242daf6ab826e76d1deb0024da36dc8a8fbee2874f3b44772976afeca9782b4ec649a34d80f4f658dc6a25a8f99a64d948522d469d27d9c1c3fcbf2edd602d73a02a55f8cb92c8b9325;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h136dd0072dc9e002a58adf49a6924fb1443868f68b1c4b6c4bb26476db7b0580dc891af4108ea86c6f0e71b3548cb7f7fd1a8eb1746cc76db2546b73c2e53b3261700fec2563e790dc4c3fdbae9cc3ed789654c19ef9670ff2de21b5d722dd2aa1db7b69353a3d29c8f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14f4d773450d3f09a95fd446fee9dcba043cfa09a0cfaebc5a6cd3b0c081dde44ac5d784a41033748b578bb440e1f1d3f2065307d093e8ec319f8e71dc972dfdbfe01540270f250b8293b9645229023731db002936e37f4512bbae8851001c09060d27c25bd773bcda2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161a285418eb1f02cbcc31c48e4902da37024b98ccd9db1a7cd8d4d444070c401162a4d0a78a9a85a4accd749d6e3a98d2d615d5f192ca4f848a93816d6a7b600c0f1a3640af9b5adca832272bef0e77b024fdcf2fd52cec7cf958ae9c83ee2553519ade07dfda09201;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19cb4efd5d77fb0be44142f8c5a3f2a921638d105b9f66fc778ff75b49662f042c0085a934b1fc7fd75fc77cf25ee6bcc9d19d1dcba1134883a5473fcb152f80b315454370d75701aba5d13e131480841e23dbe550cc5f1793080047acd9fdf68a2bd84af678a28d8b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8ae1e18180787ceea53bee7b8d0c88804bbab231200c4c22eee40fbf27b170aab397b76a228909d26504ca58c40ae0d18fc7b68be252affc5b342ac79793d036d5c13963695c0c98f0887662cd1c1935116647c733ed8a3ac45c8ffae97f6cb61af56a1b39c3a786fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h911a9afc554e686c7f64b65571e0e5fc0ea4f32a3335b7eb15b6a3a76ae10dc0bc3ca534d627ab69f6ec80ee772cd8c38b85c2189f401e256b608dbecac2cbf160351391388e12770b25f03463f80c329f976e43d36d01047ed0f1a6ad8fb10ae8356820875b96d15e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf3e18ae4b4110a9da3ce8c48522331da7e3a089f9446a894d0f50fed09c48b9c5293bca31e62f0152710fc556e15c5a9d70e424087a1dc3ce1aacce668c608b3a8099426f7312652de55bf785e8e7c21b4a5683064c890c09ce6d66be29ba2b2ec0b7ecb67d390cfd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed3825e9a66646fe228b13d5f12b2eb75fa1107d48f12d92720eeceaf1b3c7af9fe724f214db457a39d0261019cd453ea437d3533d2bfa262fefd68c8c566f6511a8c6ea05d5c68a79ec9ea259f1a81a4796e211e9a82754eaae3712b0f20818693bb6ea491f94565b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152479eb77968a82514107d49d5a79fc99a2538013a8a38bf40d520a170f14e94602aaceb83a1c3c921fefefebd500b0356e2fb6a9bb517cc263463a731cd17ece7da5a15da22c443fb9d679a99e4f4a245f255f28a2e185481e9e1a1eb2f5507af7ea7eac738a0acff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c623dcd84a7a269502400d98ab703174059c8070699532c105e30653e4eb2406c7a6a1c90bd614752d47fe6e15fca85566f878b8c9eaab020a39b5bb3e011860c6897b4ec120297b6a39c80d134ec21d50335d661668c15060bc640180f256374660201b616b9f8205;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h157fde928c689d343db388e5741fa75ac97ded1d06338a2c340ece1c76767026d67ab19cebc3d49b322b436b707539f8c3827efd142a6da28f279a0fc82350dae98b201d97b16139c870064891e447baf6519033b02d6e4c41aec5503eca5a7a9ea415a09f82b789036;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169ec619813d03ee8df7da01fa95c64ea74a65001b74df9b5529a4d43d1c22494697f748e2bc0ef3bd33380074eb03c85587debcf3f3ec073fab9d225ae843cb3f375ffaf85e57a11f769919ec4f9c0222eb1bb353720f3a57621abe942c106fd7662e6827f4836a063;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123392132d58a3e073e0e087cea8514e1aecbd2df59ce7b7ab385cb965eb3ddbd48e9ff244cf53d850ca069bf57dea9403fcc02fe677a59a65b27d100a853556370462b56648a3d6d42d34678fecadff7ce60dfd17e1775d912686d59d71e3a0c2e5e40af3b7996b5fb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fff898997b42ab17fd6a40987b474a3dcb257c8347685bd8234ec856ae403371470eabff2ba034ed760bfab7c55d9dfa88282005041d9c9f05a73d69b6c29791e4b0b12b1a60246c493a8eec2fa6012d2d299bb30d933f66723a708f64ebe762e370143e936191ac34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b513711a53f64cf3067328958fa182a1998e895ae4f3d4e4c6bf126e5e8d9a4c875dea40f002edb83ab860f5b7b144bcd43f8338f55cf16df69b55387fbf8690a9faf5bec5a654c2cddcd9081142a9a025073828f9f883aa6d8a7d58eb131ed4b82943205fd66509c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a088ce6e6865cfc84494945c293f7913cc744d9a60aca4a63660579782cf1e3935bae7df6f75ad3d32dee1290e4067c25ffd65f84d2ad3286e628181217db7dd947eb626446f5e4693b79bb4ab39bcc51deca801d67ce63f04890e67eb3e4a346530dc9aa33330309d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha00384dad12aaed0ace36bc7228a57e895237e635ebbe5b20043ed921e33c5a3a3091c1d2481e27ae24fdd51bad296847a8338de7fdf7c1239a5f1f9659f7befee78c6d57f86c856a08b7560ba4f6e800e8ddedf26cf3169b0b68474d8a1d367008cc82178837e228b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d684297b7f6947cfff34bbd71bcdf4f26443635751dc48643a1a15836ba6f5fe0280dd71108750d35f69db4a803a3d5e0f76fad87821fc2130b32ae1c8e74cd16b9591d653ebf596e0d09c5d5f0b3f13ad67ebe75d5202edcd881421eda28e5bb020fbb875541a719a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1239ebdefab5b09950eaa4d6fd467ca4e7f4225506f17aebf4f69b631a745fb740ec5c30596ce1e12f30367ae595c9bb6e3734340cbc27ae9949e7f09f838e1158371c360682d28219aa8ae1f9f856e84ec49fcb2e71cf00b96ca66a23dc3c45afe1791844f867ff4f8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe7c21b476a0c609abd8a2323c6d466af4d4a5dcb3754cb659f98e8262061790ff5c8f3986cc5a24430ae37c97324d1e2ad2a382950fa55a051a84e005a71e224322f33fcca3cb3ff1af2166d88f44132c15530115dffa3b7eb16f7bbf90aaa38aae2f539289bcb86e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbfa43d56e424ee452c917069990307c5c10d4411cb3304ccda643affc3727737598f0fde73c7e92e9dd4f0def0de9f93c167cda1d193cd4530aa948b380af183817fc881f67a0173db6f017c1f3341d616b4e8f5b1d2bf20a959ee806fbd8aac6991d700b142ac4111;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14324420a8998693c7f219ba1e57ccae55bd731639058a7d92028464047846654d409687ebd3d9548781dcaeaa98512ccae3ca111c35be641728603cc1891bbe9593b4e3b4514e449e30b13b92530bf00db93c47882c523c516939cb0ba94f4bb299c46c6459a239acc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b154bd17b6672d7d497948ae269fc6ce0a73ff2013ee66b3d0b3240eb1d87b53b3a4ff7595ad320e66a9aeff89ac5552549c2a048ecabbeb8033977319f2fc0878c6fac6a37ba6868a5806abaa4351c17cab40d2a2c7c2800f6c81994061013d878e43a05dc3a3ad18;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126e49fa1952528f116fcc788e2e9955c757d4cb4d0e833bf16208b478d9420f1558697a2c97434a92bd7e9618af5872cd4bc63bc5f8049e0448af0c1316f11979ce8de4bd76f05a4a7b9f06bc5fdafb1691eba3ed24fe3d5225ae4fe2d0103a17575edb1ae871a87d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f9e600f02226157bf905504da9c144ac2761f2e7d508e9f0b0e51458639e0a293cf48df4905e2a38d5c3390c5e7d52e19ce87f99f2bbb5b833eb1900d6c0d694205278b87bd919d79127bcd12ea2d284254c06f8683423ad8c2f68c636c820a4777bdd64bc3da9cb2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5280180d34845d9971f76b157a689c4c0fa978b8f4cdb01fd42ec288fd88586ce3981068a6a8fb11fd45241ae8c4818d9e22fa4dd16912ded8f19a3016d30f9af303560a5134d274bdcf33869f7a2d13cfe2bfec4389b06def0e54ba54a2999fcb2a210b32007e4c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1905cdf22c78f16a4819add001f2dab9317db4e6a290608b4b3b2a8f6af33281026e65033335fce2e082df76bc814158268faae5e374b4df0ff8be202adc38af92fd989efdc78cfcf106106ddc83823e028bb92380c9a7f9b0d9884bd3a19ef66cf5c796eac0bec3b13;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d58caa3a25f14c65d583ace71214d673a8430efcbd587bec58faa10776016e3d839306e8f79276eb60f0b65071eb17c0d4d0893d4219b9b9be08a42c6ef65ab6fbf53e5ebed8d1a08fa76486d8f1c825b84f95d124cb2bda0e6f0483271f63cced3c0771cfd85d1c24;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hddeff6f05d2dba4c459d64af930d118279c6d8716f8af2c2a23c04c0ccffc2cc8a781d7188308c92a3bcf30069cfe8fce862646a1fa0f86b68dee8d6dfb7ae19e90629ef296fdb8e6d9032e2a16667e19ecdad03960b6915e25b74a183b74e247d04499c8b533a0599;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3c654db6cc48d889f4b3d8f66327a12206c1bcb3f0d464b61057eeb9949d9a3c45a7937f68b927ac48baeff76daca61d2cf74eed5e45fddad53d01d922d9d14f46ec5a9ea4c7299d197fdeb5137d23cd62a04096301f32148afad88036e617b4311db508128891c86;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0b874e0b9821f8da9fc85f87b644142d56ac598a1ffaad43992c1ec69bdd03e252184b265191bb24c37a7c47add2c190ced232820b682a022193356262fc3d44e4363a70907a690896963b9fbfd57db2289491a1c52ba7a3741744689cea4dd58424563bd503288b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7211782d2c2c4abdbd895dd13dd9e06c6d337be2d60fc85bf27ec92afa23eeea40827e1b5c535157b7c8d385742ac3be53be189f090219bf55ac2abb3599e381cc4b553db6f76a84206a3ff132ea6423d121eb688c9107249e80f8e9df690be8dbe2a52c40e2a8d990;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb58fd28b18c41cc135e212fc50562696dacbfee241c7d0c9e937b450d388083587ac012dcc9aeff0b42dbadd8293413fd03e72bc50a8688d22973ebc0cd46f6eed56bb3b604e549a64919551fc42069515e0100688da293255f6389c1c018a50fa309140bb3584f2d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f087fbfc1197a71c304082fd57a89d0e23f4d4ff0ab2e2d916219f5814027708bd1b07409625a2ad173b2f688f205b6c6f3533a74f7bcbaeb7c7302826bcfe4d15a26b6c9b7c0d2ae83cee82738fe52074368b893cefe0620f012bc24ae2f9e6ff5e55c272f860b9a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e2b7433028337be2bcab403a0ea5861ad76292d812c350e5c36e22c3b3b365b0dde05d788dc2755b977b50be04c28108019fb431ea0837a1d40d163089a3ebbb86ee06a8e6ff66972ce58c5acb05342a091d1e4cf042e8819c08c19e59b4347997667c414864ff331a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h42c5ad2937c52a6422c2c68e4e29f52681c3a97d86e92d705fb47288787e4b6bf4d984e0a3a1e9edd9b78ba132b36f8a3d9c14bbd4d09d2bc1b849026f00391de69c81341942b6f257b7577df6ee1b6f38061c553a117394d249458c45032940470ae12797e0956b26;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147a13037f0e992eb1fea6818ca962a708cc18743515e68922c3ebf86b1f636081bba203bd810c5cd8a2e8f5cb6ce7155f8bf34202f2a9db6f16f50023b18ef608132143da7d63778bd29b983aa96bee4b94ce516f8b942cf04ebb621b97f807b70fada0919ade6384e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5dcb679429d9843508e43f21178f7ca9a1fa7b7e72d14212863db597baf78c9e832af8c0df5da5adcb7f9b9c0c57440d011fb22de5c07794dd77eeeaaea783d996d3e0cb932e9318247a6415d3b5e3667cd9e0dd0aa5b04198cc5a66751e2cbe1609d91959d07b9481;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4a21d64a1837f4d25209353312abd4f0ac26c79b59f8b61d3b1a3a6a5f9d267738e22b302b9535fbec5bc3fdd0b95009ceed77853b5302f138f7eb743c75707b919474a79903e3392761d18edf15773988506f67242e1145a39543a73dc851b5547f25e756a72de13;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd76a7825ca6d57dce259a363449a3a0708acbb1877699e93e703c657ac3240fe4c2cb328c79b464315d31c17d59ffa959b5bb7c995496ea07313ed4587ed4f8c4227f25f6b5c22bc00c78cce2e154b6c9bdf3cf18aa8467a699b86ac36d0ac6aa80b7b5999699b7a6e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1626a69887e2cc967c1d633c928a92e0aafa4aac40d87f5d569b7fbd15ff85be5161c1b0c42dda33b8420132f2e3f4d52d0f0f031469fcc3608bd5526995be87b37220ce6dcf8467f3f4562cf96e9c2f66a829b25d9eeb613aadc666aeb16a5911458e5b6c5d141cbec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d65163777e11b3d755cce567f2277c3c62be1b3b6eb8bfc4c3ed3252d2c7e62e1d70ecc234c01fb6d2ffb76d46c7c866d2d82d47fdc413a676754ed9f02714faf873dbac5345a2693a1e21b90863ee369e2943725d542e9800785cbfa208fa68ca14a48c11e7524c1f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d0f89da50ff88d6adc9762fe18bfea1e9dfd88eb75d03c12e7cff7090c7a918bdd2fe6259acf9bf4048f2f96a32b4a0e61f758fd0288c10f948b8efdcf3c124b86c32288b47f453d39216ded8233092b2414fb129a2d14f109a44c6d23c7e8a558b91a7e567ba3688;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed166e59c0c76ad32e3a1cd52a11f6d3891080b6ad606a24afad7310ac379a09d029e8863d7ee2e9c9874d591995006d97d3182a4738946bc174e7eab2d0fa64dc0fbc87aff58d445f2234c6afa5a178b7328700860534fff09b17bc1edbb037b841535a62aea6790c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eb6c5617fc086f59ee497947c95745a92836d9f4cb34a664466fc820c2fcd33b6d3ec7179717b4b2d65253cd1f4c3754256b60cebeafeabf4f5172ef572f0b7793bacae7ea3ba8a852e576759da7261a7f709b32da793c2b3c43af986d4b1e5ca23b940ec3f397aab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121d81d1aaf1fdab82df3aec719b011d5f9c65ccce475c121d0504ec374d70aaaca53794b895f211e33453cb375766a76a041600c50c655aa2752799b56df51fec065d9a64c99e676979f70b5c9c0c2cb1153389a52f31d350ab6dd49b77ab997ac4bb0dc09cab401a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he9524c8ce2caa19efb283d688906c1e93133654ee09bad07d384ed4293ba911b01b64d080ec9738c950f7a9aa809a1e4963e87da1d3370b6b6f3d39920c0e6d334b7615b1e9b687b40d3b171d48574788166a2188f11dfd3df786767940aab9432c5af854809839122;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e676cd684a1f147833469f246a015d5cbe59680a5857ec045e02f89803f6756c4b714b386f35172cf59db0eea012dd0642733cb4f10e56bb5a2e382e87fe6a1373258a39728b4c221bbf41eab0db9711dd269730490eb39f920d8249232360e669e64b5c99c7fceace;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7246b32591beb6f083f9bc32e9970841b30915eddd1d2a50b2a1408d8f0d4c5cf214c32c0eabd3efd144d37f4ab8a4aa7a81170dba90e30fe73d1cd55e2642f196cfb0153e9adf37ccafdc8d09e60054fbe5a7a8387ad825f8e8912206c50cee8c3d6e428995339d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f89c72d1189e9316236a5b36327f6eb22280fa46182c790e8723794d9378188b5a4e8ae5d1bc2c2541e5c3b7112fad145dd62d3173c6d2704410fd41e073c42381fbcc02b59874a82d10213589127e5f35d49009f7afdeb98639b6a75daa2545dad5cd7e72f33fb45;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b102e0be0142283a2c5c7c46a7eb9006efaf778f4d3639ec9c6e007aa3329afd6d2270ea98b90f0a857401005de2f16813c21f57d3f446443c1dc62c2e4dfeee651918e25f36ee328ed646b005512c25653af8393419716a1b7dc1ff4e5f7e30de1ecf2f5e5cfe6a06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e3fcda24a83e152a5a3e5fe57d2c6c75a2fd4af7d828ca9dc891fd0ccb52322a4a02dbac7291102e3c82085554f0f36d486f088e570bcbb7e5b1477d4e71a1b0c371a8ac085d3ee6c066477c3cc374a728c7f1989f2aba771f6a7922429b7a851895b8eb76b166652;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb0d84d239f62bb576f758f566a1034dfdac44b9dcc1ba02a2b27671eb8254ecd80687b8f44f7fa9c58e9332b98b1f2478b0ee46f96cf414895272a6b5d8e4690244fb1e24fe91d47e56ca570ce02c16048d5331c9d3b636154e1ddde520334c0c1ac746d2213fee65a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8de33580bb312a02128900ee750c3a5502bdd824705972a7d245296f38716585be4e559ac316ce5bb74bdbf9275fff134a3ae4a7f3a14f3d6428a1541b4eb1f68ba83d8715bef302470f5347177f99eda77183087535e601d3b46cd274d68a14718cc55d973718b3bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67c0a0797e7b6be4f36f7e6ce9a85f144cbc15fd0683effe013ef650231fe0d849e6f69d28bf2821149439ff421ff8243c71a47fbe0ba863a2fe944d91fd567f7702e9b843fc18d61a06b75237e0249cd3a7c6eaa66a035c82da7f9e1b774c0e8e8366952bb6e2d49c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9c8f27c5f5f280c7a03ffcde6593d54000b3fd50755146c64b390c89beb891dcfdda5984b0a7639ee988162132d233bfee27a58bff9b52a7744a5143238a0699fd6dad76d1c77741e3799761979c3b25e3303c9d3a325a21b5e6f783d47b41eb72d5f9f19c1bca17d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc57bafa47469a11a34fe9c50f8ecc02d59a9a541b26e96292441c97010ef19938ef5c3fa081a9100139ae4ce107c1bd1c1ad9d57cdd477a63f95fd258e3f1c1c815c02b9b3dab1894b00cc16261411e33f94c0143fef04d393c535356567de40c7e7c04a446f4aadf4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5967987d453e6dbe8c3eddcaa0ad95114d0d113c5c3c15de0c2d1816c14ea7bb75b28eab9f7644ff36d71d4029321472cffd6033fb58dbd60f75610670bed91677c89413523750cf27341463fe72a251fe604fc98c4876f3cf047b2f73661c93d51f1e1a947ca7a033;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d6633d19c3fa5fc3bee2b836f343a348b1e711b6e292717453263b25d433e255d55ffdb85d5ab8f6f128723f2f14b9cf8de46fc59fff870187475deadf8376190ac3ad2e3169abb957d66c4d427a48b39ac7245e432a03f8400ec9db3d03e1274d31fa25101ae50d4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h223cd449dd99f1eb6619e1f322e82472b79a0e8cab56aeb1fb5358b288b55e8a1f5e5c8c7427766352a6f102ba7cddd5fb04866336a95cf7442fc697ee7aeb747c9eb6af1dec1cc88eb74960332fc90da8c54406386624b86c6138b391b1b04fde65471c3809ab369e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e63e8e68778174e13c8306db670904401f83c198d10ca2b488b74cadcc945ab46a7c2fd8b90213ac20f747c5abf410fbe3b3aa4bc6030808ce2f7a07b1e80691c73b2c9be1a78720be5d76c192df51ee6ccaeedcce1be0895172523017e311495d95bbaab21686e8d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8b8d2accea034f6ff67006b42ebc41c2641f3c81f3c985ee2c2a2d36ce725dfcece73891e70f887c70afc5b04417b293eeec07bdfc488b31b1f54b12f353ad9e4e38a4ded0a91a74ea145d01f3623bc44052dcaa10884eb4f55ef80af627ed1f35107dac03545f930;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h285256823ccaf0465ea37bdb0635f1f043f384a2e743b0ce463e52253fb1b05e0f20a53f8e98455160041bc3f4743fe840c6c2d14dad34fc862d7d501f1d4a0bf045bc9f9b31d0c21fa47afb745ab49f0d1ce15ab7de8888c64dcf80897aea4a029ebb2e0c9ee28f1a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc2aa65c706f325c71585ee073a7a21698f4a6b5cf3160462d3b81e8b753a8fe931c2bc1d85cffebb4ecf58c04ce015df91176d80699b22fb4d46c5ff2337c49bb364e23ce91f24e3f866ba87d87f6b2a9859bb0a19226f3ec11711ad7e59e88bbf61168f1187882d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bd0690ec2c453c95e34ac842a4fcf69d63b21b5d009802a5cce05b86fb288d269f0efa4b23d5148e5b433309f1455cf7cbcba3c2a1ac0cef25acfaab38b6a405ccf73014597436efa309690db48b04279539323acbcd555f6c3bb600904e54b4a36d9040a34ac40ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e1994cfb66194b76f9160161da8f643816550bce99b2219e18bf9e3a7fdb21c986f46be44882950d432cf0d98d3eaf5fa95e6275f6ec4c182387d2e00c5989eb9a4c7227d24e28a5b928c616055fae7da366862fc40409c5cf624ed610694d281fe7306fe1a316181f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130eb05909f4b47e0a869c106e714b9a7b301cbc62ec0c750f15e535e448d6d0bac83d8ebef26948d79c6fbf7bc027b0324e1131f67cec430c2e2446b49c2ae1371aa57654c8f11fb76e218ccedfa1531eee6feb4e49b4ab30ddd079c9e75c34302fceb9aa3b4541451;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134b9f875c913e8c08001a20cba0bf4cfffda5288b5d86c13ea5986eb4427e7f9236a80821ddcfb370578ce991d293b4c1a077dfe6cbd90d5c467d928f61deb5ae24c7b46ced94cda87a0c72b7a6b994cc16bd2b4cf46505d6fcce6c363304aeba80a4e434d3c274936;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1242a50a97c79843fd429781eab13eb7ee12d4e253d4dae63f4ea1689629cf22f398041eaa6da59abc7a7ae6efe5302a35498d4f953025c780bd6fa176327582ab19d1ec45477f853a2d66def3ac9562ef176aba4869317f350d43d466a7b00cb4830eef6bcab915526;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122c0a4e760bf3d0dfcbc5d02e21167982cc4f9568cbcb6fa8d71caa4dff22a8d6428d676439649e91bbddbe52acd8f31bc23f7ff2519769cd0dc96bfcd678a35e4b582e94c7c4a413ac8c9c375dc3049405718d5e14877bec12f54fa525ba2a6676a3431fb37960a0e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8f8d69844a032c30743ba4f157216e3c44621c521e982bac3fd92286e4fe94f73c2831eedb21fc8748eb0363f3d0929d05112e3163bff17e23f51d85d4bb92e9fee3cbce771c48b37e1eef6251dc67140da35e0b8895d2ce7a8fa6b8e96eb9599f307ddb58b8f078f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb111607c86146e2be770fe971108bf17df80f0900038cf97070a75cf1e6858dafad42eee63bd04a335785b4a4bd150408b8948c2a6ece2cf0baf997afae9c083602f0d3415a9c58540f29c16e4ccded557c9e75b6292cf1a6ce0c639ff62106fb199cc510cbb15213d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1293bcf77c5463c66baf11421b61a324c24b99cb073a694aa8e45fb84cf19a7a5a35a1696be00e1d33381a2a35c5ae58a678ab44c5e9f092a4809ff4a3f04d5f15b5fbe12a52e0f758d09b0bc9b4f3c970abc051d313ca9b0d3d5734e51aa12d081e8d4c42d6893a6cc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he7147d7e0394c429b551d06d509a0888f41c1ff1cb8d7ac7c7a1844eb5c61ffa9a3d5673eca59454f9ab36e4af0fdac88672f6aec8d32459d21902f78c0e8d9999e2ff5b3a6e80b3692c3fe1feea7bac7142e1ff6d266df8590b9bb5b69791994074346d7af7278380;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ee941a38d3a19664125bb3cff12d81a9f89e2c79a2d24abe6df860921a553a08dc71cd60ffc26016f662d5810204bfff3f57cd440f07e4ba6cb05995edb7431ac85e83143a928cd1fed3bf0540c88c1b84a87d04aecdcd16d2c98fe47ec6532371bd6b2d6a52b5be4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c7d319367b96e853b743ab88bbbe73548e002029cd6ed31b36fc92fd0992f0894dc96e40268aabe3289f7e8c48b9dd3dd7b4d1909875ca8a3c475ad1a97da4ca042c301233fea8afbfab51d02dc648758193e5f884cb8a69745337fa7143f7506a0207efaa9d48320;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15be90fb0c9c1d37be85949666ee5554b72b67eca1756d7e3a3cf8b7f20d621bcc41c63329f0b0135fc9fd61cae2071645e0361b08add4e9e46cb5977cc43d3e7339d46777978af85841d861a7132c8a998c2f3bca7688b8778164d337684025bab6d9d150e3382a7ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130cdc8811935ed257b8d31f1d1db8f8df466ef39e20579ecc625d2e353e9c5b7fa7586d307963a9dd1d76f0f5607f24ee987c7dd848364d7a866969d3eaf687a6d733390540ac270394fe7783933777bbdee9a841729191b865b8090ce3c69b4ece576b716a899ba61;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131a40d7b398c642088e7723e808f3b2c98e53a4225ca9939c6159d5d782df907d03c99e8a518fc85ea691179858a2611f568ab3feb19abd25fc57a4ab9f386b06fd7c2ac22158500cea3aad05032b56ee740fb1d2b0c305a95687f5afc1c135b695a943fb55266a04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79c427c532c16fb63064e634eb97ab67dd194ce8ef4fc7f2c416744bc836f1c5e263427083a43c38ef506f41dcfc5ce19fac9db35b5819746c206d6815e37c03d2b6aab55dacd952cd06a1165ecbe5052fd4684da51c0a4f3e2cdb93f9935273960ffaa46b4c5fd7cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h223fffc5a09d122b96dbad50eca490318c1de0924fd1aadf9fcf808daa2a92de16357b1349f01adced5292960ad97a825c2fd98634dc87d17874d843df1bbb80776a5d69e1281ffc5679179f186e0d590e8c48f0ffcd90e30dac0b6cfe555833e65633f84f2c8b82db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfe7046f570486ee18ea5643c3cc09ffc2db261362a40fd32a32b18de29d134b134444b287b96f5f88c356433b00f77b974aa4eefa885b40d5ef7afb618ebe89a57100ffc26c4b46de95de17457d95a3a6050afbf7b435a161143b5f195f76f7f2185e2042c29bbdf8c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c595303e2772ce772a9d4e16452fdafc3b696c68d43a1bc316b509d6d20683e9955d75de976bf813a5528762eae546af5db40e1ca6bd3a19f494ba29766e719a3d966c776168638624ab7c6a67ea455c0ab5b934420875828b89ac2a6570499da1fd03e140eda50ad6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f215b77d66d9c0c95a51872c8068ba473cbe554802c943448c42a69e87930e2eaa94bf01e30083ed75b9feff0be9ca0e068897be281e2d70dbc773b44fb763b8ba9cc58191f84d81867dc617a627f2716edb602b977927b8db0db9d7bfec2fdbab1fa740151c123bae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6bf711fafd3e99807ad14c820fc4c316f305adc254503efa4c344aece2d2c12ce73e65c46cc686a0748dc171779939cbb82fff2b227fd4972cdd99b4b7a802cf72e42abd6af85495efdff89adabe87767436b38174c3004ae9c73f75cf4c7a3168af3eedfb26f1cb9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h144b6e4799a37740103bb924a705b72b88d1f4c04506161fe17e60a885d974bfb9ba358ec600e0ab86c566caae9a13e181d1640d674f20004166cbed2d837eb570773889390d3b2418cb3ed960c9178e458ff85643d140caba4243a8e7f1e3758a28d894f758cd35a1c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc8b872beaa9b165efa0c647f50b9d5f1868848a4d5866a495d9bcc4909279143eab712178a775fe161c86bb22f33bd396ad46ba7c1717bab71ffe41ca640a4c1f1ecc89230d5172255924d66ad4c3fe45ce2610fb992f9b6cf96d7f664973a3580b4a390a999b3f22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1da3ed003e9512e26cd8a3ec42e097eff072d095b618602de86518e88902c084df26653e852a98f9b3052e2e0808c55b97855764750183f89fe6c9a92ac869e854abba4e60a7c46ca341aab0f6be0db9c621cc0f4ea65dbfc51cf2096dff3212c94b66c9e134539ea52;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1b1704bb2629a3c0ab4d354de4d3b61c9fb6d96cdf3df0d45817f178e1bca57ac69158f188bc017bc59d54a96d8269029f9d2630845de9d63aa5a1545b9bf50a0531ce22ddfd37194fb9a4e419dbd50f818ce6c5a329b41aca9cfcf0ed904dadcc64662136fc68a75;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131a0bb2ef134d7a85e0d90e743b26cfd381fffbf96c5eb20bf0789c20df07e2e2c2451ebb78afa2f7d24ead84b9559a2cdbe8f4bb45ee71700f10436029ce02ad16501b81749927f6be22a5936b6f84ad29451121e28494de27c6d24552f29b50d2aaed6ee9b56a7c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce9364d951432f2bc8e8d3c6edd63035cacd6eb245e920b46e04732f34a30c0ce917759c5314fd8479625e806e24aadc6be61478315d8ae6d623750d750d3cf3483396f7609d799209ed5ded2597bd4c02d26e20d942e4009c55fca6e39794297f91a43d375789c1d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a52f222cac288564ad0f2c9095f35e932c3852b3e9469718ae30048aaa80789b826bb2eda198e447f397c7e4a7607b9177d6d767f2a5a3fd5de2a10aa9b9ac7f27530705c7defb06ecb8e11b2a8979728ebfc14b29ea9fe21c65ecf2641a1c95c54142e97a380df7a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1753219f6b3d6572291154adc2d66af6ccc3c745eaf2c36c715de06e3fad8d661061c6950a096a2bcba747790f9c2eeaa11d59f1e7d731d975e24c8fc0547c2a96cc769b0ace9f36c7e203f8c0d7cc8c9f2ee5a2347d7a466af80b73d617b8d57db3bcb9ad4a8b33c48;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1136e7002c48cba8eef7375112b0aa2646e7ff5a076ff06e95ae31a34bdd6eec13084dcddcc7840c5c84c761362e71c8ba5174554a9b638e915d010f1f390366f11f9423e51c4ef61798876d4638a193a15140b85ef66f5bfebc6229732a0bfbbc081d04ad9627a6649;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f45b9d87e7d125d09adacfda5ceb3c2cbf244aa552b1bc4d1596325b1f748ae1ba9eff64c60cec36a01b1dcf16d37909e97122aff8cbe592c3713be694409bd7adcd62316fce1b6dcd4e1c77c8c97da9433aead405396eb7e82f41b40f1390387949141556e32212c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82a2d8f43899d68e32385cf3ff32b704128e1e59b5d5a8436f33d51c37bef3b38acd10ab6f5a28778c7c9f5a2a5b1d2023fa6cd9b7713ddae44dad1a034a6a8f4a2bff5896b2296dcce535e227fe11a2735f10a1af2ecc9047a63ee25de1deb098cb7efd9f1beb97fc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e386d2454f6686e63bb1877dfb6a619fccafa6ff37c710de256d233a07002c62fef43c401e5eacc9774e0835415cc80ea2e99acaffd76675017de47c7106bc78ee445736d5ce69af1dc7777d07726321eef9b2d6fa26ef7530bcea5057802d2284c01be0760b9bd30b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b2f63f39d3ee957b5e0fccc576986373a01c8911df43516fab2436f1130b82e562a9cae31635cfa08aa09d2a85b2b5784e4e1fa4e437daf009be3f88afda0dd79eb3424f10e0efae99f652fb68df11918105b7db5f86591f4ba2f77c9a012e50f6b75063771489c6a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14767238ced019976b9fda09f74fb29d7f673afb80d2dbf8b858d37eae5d83bbf92c3a3224be071440d4853bc8eb43259cba728c5fceee423fa1726a4cea0b569d5a4287c74a5768418624a4807ed0db60e59421af1b6a65941676eeee6fdcc315c3ad292e38c73a251;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf1b9ce3a11a5aa8dd1f8ada3ae5020f0830fdbc3692b54f453f253068dc378d625f5d61ad6c9309f87395af266251429b534ce6c6294a7adea62af1145398c2ab8af4074791ab4ba0925f51ece035911eda92431beca2a4aa44cb32a59a0231d75e666ebfd094d38d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h114469f9b9cbfb4f9022f051a2f5f460c9fae3f3671c75ba646467db483140227b636da4e01ca0eacf004fd5c62af1802db88572ec0fb047436fe745871042a7fd727bd48f96087fdd57a83ae71d4d38ad854ada2c731273687aa5986f121229c9536b6507a2b08c148;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h87d7a40fb7c3e0d922fd2ed50c5d8e225b733e792ecd83e76dcbe642f0d2c145ffd1a3ad5935d555e9945782be76210a3b648df06d78bb49f21c5f2ed7e35650530eb266be3cd9e2cf8aa37e5ff06d221cd8d400e9b7855f2ede0d2f08621017b660a0597d3abd3436;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc61943df78d3017f9a9a0735da459046521dd4f11b2079a068b5d7e95516e23d6d94861de4d059205ee34864445e520f21e6c1af43053c692e09516c8b1318638d92e4e8a28c741ff9fe74b9371cc88e96d450b180d81f26f7aaf92057ce7aac2a28353f531cbc03d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a10901d92c557e1b8e53b83276c6490ae19f96771cb2491e69daffe30ac1908d4ef8e0051964b2892dd6d88ff703c5cce4f16d3f0c8625ed67bbbec308dd71c4a470c0c71016bc97af65f93c75521238cb8da46f715f79e7dc4cba7f8a62484ddf5257ed1cfa0058e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16f381b0044a181edd29b860adb7e9803bbd6f26600e36048d2c6cac8b09ecc13d072bf145cc16586cf7a2a534e8ee5679fc9e130c1f163c53f9cef45f116cb08ac2b3fae23231ca822815947073fca22bac4ac29ae4fc77c68655c5dd1d1e8a2f4a0237103ea0f88b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6686e3148a1636026541a25921f8e5bd90ca6807d27701b151dc680d410699f112ce5aec1822bdd6fe918d864ed0ba8a5a64fde1eb967901efa5422bd990e634be453fff4904c23313edc195cd2b0c095f15f3707332d37e7df7763669ee3b1531764af10db4b28b77;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c9eef4e838da8cc9d715ed16fee36da65ee82ed1390115220ec7891b461a8b87159a52522840e69679ca13440fa812664a1c191f6f3141e102ddf34597c983582351685ce01dd88af9138e0d254fc5709cbb7039cdf31c9682b7e69e3fc8d282b0b04163b4bf1efb06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b035083bc55dee56225584e205f20e3dd1a84b77a49bd445225b44488800cd4a3c622eacd064bedc0a873610c8b4b9414aca279206a926aad0f08d189b30c07478abf5a355af159fdfeaaa09db030e26197364d3aca7156dff113d4850b00377e4015b831631f684bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11de6c3b44c92b85a8479f8946bcb4ba6ddaba8d0453608a1d24fbc5cc09b3353297baed1f42528b278a44d051077db7eab5b3cb6fb18e1f95e8a1f1e83b315849f5fe73fa9a5f4f40b22b667fad5b4f6a66f2a9229136f0ac6e1f7d7f02c254774f0db1359d38c1693;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d09c632e1173e0864129ec1f7d95a03a9343e834b41a6fe5a136469d3036ad12f01ee525f9c3b7b4c512411f2b718f9df86c3cc609a8294694bcb05e204d15c462a00c15272f7e19ecf625278ae84e487013139e56f682d7c62805fc704415042163949b45243ab8a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4c5c8ab09c0aa7ac5b8def65737306ec85ba92c64b1458c555fc2c16443256d03c4e3bfdc8eca50783e5e211418957561c8be7292b11ac607371a7f07f2d7278598ca2ea6d2bba68cc7f78f7ac236a12c2c2757db9cce9af775e81ed8df93b60a6889ba1fb99a83e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h438d9bbc955a2813fd4597bf85b08f879f8d5fa1dce07aebc6eeaffd1e43f5cfd6708fee7ebd4131d948387f25faee0563a4038c76b62113eafc94e376d78fbf40f28484b8cd4ed563b4cf3d9cac089fe1fb7fc00ed4b3c20cc540929a7ee92833ec563a62cc7a231;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed59fbd3066e77900770061a2ff74752d2226ec7f8ee2dcfc8a4119befc77777d9723a20b15e674a12c928a842016afd8c56173108704b5f38d9bff1c00821c0ab7837dc7de692dcb25b85e28792ab4a665bca92ab53899517b7348154d62116894390703f021eb04d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfeefdf913e99ddaaa13e1289e34c3c46c347d4978feb4b57e1594cc0a09d48095dd7f3f93a2813910b60f9d9e5fe025922ebd889924dfe1229f8bb6fd088b32ab4e1015a9c22086aa045d9633ada8c48699ebe9ed5e6522d3d42114f0a1c58f378ac216b9817bd5c21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11a7e26c08765072fdb48c70a7dab487ecceef85d1b9af8468ed9aa202bc95cf9f267d84cfbcca8dad05cac6c61ee76a1b30f74af8c10cc6e5de44ca03fab01c400b534d53e45a6f940244b66bd846eb2090fb47a0cdea10f285707e4a42a86635eb24488cdb89b3217;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2e1d957f6d987c1f2e691a6e9645ae2859ada253e3229cb59bd87a0e9a38129ea786059a1e7c979f20ecb1cdad4c5331bd268b0b289d744b5f15ea93e3cd98329f9a1086635cfe162858604690a7d7e999bc3e1d5db95f3ce9131063146a8bae8216f2081ef7dac57;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa33198cc57c3b400bcbd64c987e308514f0b44569a11ff1fe42475a76eb355a96183d098144cbffa6186837daa324320127d30aaf6aa186fe33ec2e7982f16584ce0584d75577a3288aa2c55c9f77003ede740a161b35eaa9d9ed8e0109c15ca9e24955906ee67efa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed4bc3c41fe361b7d50e7c29563f0fe9170d3a2333b223019819071a362c696c1c86c0848615bc25f1c7bc6d808ce7d169dde42c1cbbabbd05db24eb27827aef2b70f2232d5b59fd9697ffd20d4518bea09c49bcbd61fb99ac5b904c26a3f00fd37f2f7b4def8adab1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e4add48d7066540b7823b4c5ee5943e663f92998672368801aa635b21961a7a3b040052cb514de9e5e59011c5516b1071e64c97435b130116bb9bcb98970d9cc1ade9028fa487f5ad544d52412125dfeef0fe004b4b18e0ad198e50d52ccaf6c2ea9d7d0f817b4378;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffb6c3b923df688df5cf7385df5c66f622cec0db3b8091ff5dc4cb8aa93634e14f7a61e563382f1de02ccb6c8c50aeaab5010c70a324f6f476c5dcb151c4b3bea544245233ec165bf2d2c31922fa6237a43dc205948e02bfa95f763175bbb69c31462c940dfddfd645;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d32600d41cb5e2ab0ce7db5d76c56711c333167fc1fd09524bbddc91e37900c536ebcbd99e618502cfb1de66883b1711ac21adf03b7560200bd07263f2c5ed879a929a1445fb438b6ae319d236bae56708ece5cc70160b93644a628b77a3e7459d8ef7545700371099;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61bdb73660df8c57f206ced810dd07d0a89975f1276e910566bf530b9c12c30653d605cfec714922ebbedfd1759e8d25c762054a8a1eaca08a05cc3e48f4c89bf7521b9c38d9fe8d772999d2e45ad39ac25efd2c6675a44d5f27ecef94737a56a09004e0b497ab6fac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a993f958ea72a715f21eaddc47311b170e12ac66b5e3c7015bf7cf49c8b9325a7735a8ca9ea88b140663bab7a74d669a3068d0ad7ee4933901c99995891c5537db345a1fdf53f5e873818b8e7a71d21bf5369c68cb2d0f8b41245ac4dee2a4e52120a61c085c627a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fafa92556cfba9f361851dbfe677ae308d4454da6315452eb9145cb02cc849a76bb04612bfd13dd1278ba7f433ee46553e4c46ed6ecd5950c20d4962b72ce157bf3780982ac97224efe25632c6cc6605fb7318af4cfbc3a76fbb30636c721eb624ca6b067c1b7f3f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18404f7837209cb00e460b2ca24a98d94dc1f3f5f0702271cf82da6f515a303ca4d5f76e6000a35b153f9101f83c75f848f26e2614ada7d86150cc3535dc28ed5761c156d81d02c5664960c2279a80c7778ee7d87afceba50a1f55b14aa6be75463f42e99b1603a72c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f2bcdfea31e086a5470ee844f4586317bac00670dd47709d0d546a7567cdf7d0088db018ba91d3534510d3dbd8d05bd66d2ad91eaacd6c026ea9ab13598340d5b08438d08788727d6c893dc76205a779040041a32c3a08d89960aeeb26aa66a1b1bbce73497fac41e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfcd28ec6f1ab0e23d9e6e64290a934708f05405fc2727b65c74d95edf3245da168c667080316f00796b7f9b566a5bc7e7f9c05137a9d31e77eba56345d40f86bb4e6e3139a55e82bc168e416bd6d88a1fc8805c975be1b4f42f603da699183ec20e3ff2727155ac79f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12aaed53288787b1f983ecd692e24b5ccb75bf9e6cef9f7d19b68597602701e88041e3c47c231382e3dd3a8f9a1cfd03fbbd98e379b5d59f84e6e54a8af50e9b345fe10db987b583aa8f0b3998f7ce31670212811d0c0c7e980dae37d9f3c26f2d85427dfdba6f96d46;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4430f245dcbc95c54270c84c2becd6ed8de7157707259b10ddb1e2548471bf3f89aa9874448614b31ecdac4113b0a880586d71830add5b949c7fd8659661d495a391fbbf3b7629c0c0264bf872b0abb0d614d4ba2dbf469b5f40572eefeea9de0051621f428cd02ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd0406390f104d6dc400bf6b015999d1a84d20b503fa4725baa41efd787e0e915aceda40428d750acf9a37c2563bb8d0cff6a939218d642fb02bb2d8903c9b41d4ead69aabe2037c10c9b55422f4346f3e23570426e8a7d2216d74f4bb999bc5f8f0c9e575686adc6e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca59a8700d8de422c7aeab23cb074d246b7956473345542a75ab49aefa93712425c008059960d59961a687bfc3f7fb1ae0f96941016ed584dae25ddc7073a9452767a4a19180fac6f895255238721adc0d72000aace8e41bfa40f6798861d285dd487458f116d0c121;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77a500c421d74fc4dfa95b65283b4cd7d7413cd9b67115e2b8f1336bfc55ae2a1cfa7b2140f3f46569dc46cffd675c54b1cd09f5694746d2a93098da34a499c7424d453484b3a4dbb35b89517200041299682da9bc13797ea1366aded79cd04faf9c1f7cb02f5e8d81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h314f639dfff4838ad0ca788e37ff4132e5c0fbb6946b354906122859d15ec5f400eb9efaf65845a55e0d686ccab5014c471616576b4d5490cf5722988aeefb80bbef6bebe89ac58db84e1e6b94e547f72f36fd80bfef079529e664d992f2a6b98c1a3030b7d05711c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d29e1c6e0c33fa0b08ce0503a7d26ae733b91241e032616956e92ab2857ab6b816c25a9f39a304fcd184a1cb199c878c0cc2cf9aa0c00efae275ffe9077b5398f96f04b590f158802f70057a9dda8b50eff596c0bb5f3372944ee626285df91f6500bb512e8ab496ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1254b9ea5721c92e6f6a7b8e42746b40937e2037ee01cc8aca5f63dd5bb3667fd01bb5b0838664b31130da961170b187abd9add26ae76b0056961dda83a430256701a763d689dbfed30ad90c7d6126cd15eeda3819e112d77243ecd4e03b8e3e321bbd8c9f5d9a62f78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c53e774fbfae18a6d92093c90de37b93fd28efb61e62e60b8dfc797786dd887be6879621ed1a3fe049579d2c5d9e11f84bfd5db8cf143d56ce294672fcc413885b0f96d82b94439bd6f5d525b02991c23653c2d680ddf41ee45d306a7e5fcf8ba3576520a27b33409;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc841dfb839fb7a129f55c2cb1c568d4023454511aa24830b7da874f48ea8461a606dcdc85fdffdfdd06b5f9938fc03465282df71a6609058478f1f9921a140c57fec750443a005c012c842a94029946070c349ed9b1871ec02fd1ec930d660b2771996f9a67f68d24f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h393ce9248ad83f81fdad5f3f36d0dbddeb15d6599310ca96d50502903d52aaaeeabdf67435505486432df21d90540acc0af5f7dd4be232e180e60f1040328126d0983fbd7329891f3255b5c9927f91223c0cbe11929bb76ca9ed5b26df84a151c9286fe5df4d9001a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff18a3592818752eb1666a270473bc818e0a2b3e6f8f61e0485d254cd46d7ec9a585ea11d37b2646ac278a6c993c3b3041a4ea45ebd3503412e809970964da76ffdc85e4bbb101ff12ace77352449f6216cd3745f3b27bb6b10df75a5b72e6247eb398dce1d9bf8fd6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62c213d85a008d17fc8e633d78f513107aac1a7463986efaebadb2143deebf8dabbd28649cacc7190e6e030ebf2c90eebdf4bf33fb30170cf81764e2e778807308c1210ea9c6679ae377c39b465b4ca93c61d2bea84bbd55c85760c53badc6baf1b078d78f214a7818;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f3939cee528fc48f595f8e285614329ab6d9144255349bf5c33804b5bdc9b9826d775c95f9abd23cc0087d9de34da0320d5645ff3799159de8299f84a8b7a64cd215a7b7aec87a3c3ce81d8f37710fd6463a7e9866ebaf6c5918e1734b4e961a38b439880c1970f5f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f7f3414dff4a173c6262cb4d403ecc66e2ee22c110b0f72fdfde21a7c41268e33b08207032399d916de6988f6a29577edec9147a44058d8969f2be2befc96d85db63dbc4f6688e6e6e49846b89bb458b01cf5083ef0a89b1eee8acaf444bf807d3891eeae80193750;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ed1d0ddd4ba99348232cba935ceca61eff3775a451c33a3cc735915c3660f077695d72afaf323cf3fadbdff3810f1e9da27701882fbc3d757213b6108085d75ac92bf8562cef4b4a15b3b3b5f1845ad68668ad2c9a2c20ad2dacc0dd85a4272415f01a66f90ed9c19;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8fc70a21a0b88a18ae05ba8730616a9cdf4693e9622e148fe9c55d453a339fd9d82c75edfd3e33346949a4f140823d7d2daee51003b01db43518dc4cc544f0cd429a4fd555d2de9a6a7dbdde1c31e0c7582f92dd0eccf5540aca7a565a73d8121c68eb7f3520082a6e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1757a48e7bc844b3c6d5aaa22cbab47d9dbfd50fd24aa2b9e25404534c67ff9168d0b00b8721040dd53afbdfaf57be4d0799ff32701715feb255e6734dc86f0e699cc8b00a0da728a3593fb2f1677ab5cfaffcac68e7424f1c75c79460cfef9a77a02380ec012cf4bda;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbb58196f5870ad413c79d5ff27a095677e76ad9d9a1c6650508eaf98d5e447353d19f59eb838ad789135b1948a39297909f1ceb5b1c5a33bd7ecc49a353c33a3236abcc5550288c1a04659e7e059954f0aa0e84ca3b4f5a8a742f251393cee39088712d6e14951172;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdef2210313823c15631993c8a4f6faf07d37bfba79e0b111e82125f6ff750368ec9babdfdcd6ced5d56e1dcedaced4ca4f2e88ee1e1426cbdb2b257adcb28809ee26808779bf712fcbb74a8244eb5ddfdc5b8011e62c0b85439bea07be9782a0073e9de8a40e6c32bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c71da12c7173ada3eeab5b51529dd6362bae05a93e236cdf170513e5bcb807762dc0da738850180e8f746961ba04779a94380b309a80b40220e13b270885b251631f7923b89391953129bc0242436f4741764e622a7c6364d5c0314d9a2f7bb26659a08580d8432b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1934afeb5b0f15036872f0f11a74693df08a26eeedcf5eaaa30268855ddc8aca8cd129875dc05bf4d52fcb76e78738f84f727a575fc377d3d2f07ab98086944f5ae40e88da283bba8654f8a963a1efea7c9489753a7d0b9dec5b19824f5b8e7dfb21b17e33c494c930e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0e68a5625d3ea3a23bf685267fefadf440f038125a5536cc76850646cff03848f5b71af4e49a289b29eb2f55f69db8b46c6c6fefa6dc64e84e715b47c961a47a891c095f5664a22496561e42beb81e6923bfef2e7c70f19728a04e62447536d17d9388b7ce73cf4f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b7d05740d80801c6be4a82aeb53961d433639a3795d742db97fa037f619fd1b3d0d8c7305e5bad41235ac05e8f0c1f278b743a0df3b37648995d2a4619f20321dca2b17aa4fe8875d52803b36c9b780ce7104afb395e58d98e66484c867f9162fcba838431625fecf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h733cb14fcdd68e75b734f629b6549831d6dc7240ba16c71af45d5c6b459cb246b89bc30eedddcb865e0807737e51c4a012d24d8b916ba7613207b1847608a66fc891bdd9771242529215dd1c5417a290cfa0de6579df02e9635e3516674fd3e6461aded4e888ef301c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62e3a9ade04de51868a132e6fc947f2df850eebd767aa7f782d4f4c04a3b404a47884193cde538e090ccf9156cfdd0441c482c1c81806e4ef3bd29ec2c3f1f9e6715477b999a34d3b349997b1685e79f28873f2dfa95156a3763ac341bd1f3cda3f35ab6b4c7c0743c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h194f9d1ee6197275dff6f3a0868f07260ae08176b28a96d1403ae8eb8397face051a7c251e9e0fd77d19ccc5f2ba8c1b89c9e90b3837d9772fec24bf84dc5a149851dd85ecf7c743bdb7b02f990b0b2eb217514b524bd62c49321ec2a1fafa29b2515a623c7a516da71;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9e0e8ef402e2ed8ae8ad9e00f030bba52243e5fa200f7f6cb8d42de8cba2d77c358adc0fbba5a88b4576db50c4c366abbda827a09dffda89958e25aa54f262d546452b9da76db6bd064a01e39bba53cbd82cd56c8f4e059137049d17adab878d9bcb4643f72d00172;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15378bc38434ee2a176a87a11460a0a3a495e503cb772d3456ca303e5bd4ea5c31e7ca5b0d5aad5a2ca32b92520d20a7ad7348a005489332c53a9004821f0bbe3e7a147eb526588dae14f7832d5ed6463c2ef3c1404899919c45f571a7a36e2450f051d433ba0d77a76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13243138b384ee954bda14b1c509f6db44eb92d9804bd932cc9051c9089abdcf7ac883b44ba266b874352a66b8f1df5ec47447b22945f94bf611a26ef684fb40e1cb430833bfbe7d2271d7a01f5bb52e13da11f821a9e09e9af20e82e41a0027d1ab6e0e823f7aa4713;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e179b0a8c5b975c2d5c96739f8edf9c5dd96d4cc2282947b16b82f056333b62ecb2636dfef1851e85149ecf9cf448eabcd3240987c51db94cef1124e7b8d6478b9c6655c0d6db54caaaef8665e7e0e971ce339e37d31a81c1161b8a59c9fe77b202696ad28dc1693d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2db2359891490fbfc6b8eec6edfd9bb41a02bfb89a94733b5876db1863a50eaee6ed7693f21d107126d2f0d1f25cf447b449a5f54469023e6116c28d6756d0bdc890f83dd3f7c2375838f88da704629b1fbbb2e262401a13c5c7dcac82e844d580cbdd0b13900b242b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e8210c059e0d02cb774fb695ebf0d389ac0143d941c789cc1b5b189c6d30ffbf6fec823525a6be294ce66b8c087f7d267cc50f0acdb156120f9000a234ac0962e105fd8e06168acaa3e592026df3271e57a35f6f0a30340223060bded18388300a81952801faac3ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19dd7d3a321b6eedea3dfcbed1a569bc4e977d567b4226b0eb06acb1ff37fb7386d5ea9cf808fcc920b1ccf297e8c910883f5f9ccc2079c4190f1348985e12aae4a23d570ac28ecd5cede7f169509f4a9140a186109e5af578ae80305727347f4646b7b35a159209389;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdefb771dca251ca297b40ad111cc008897e0eeb37b4d82a6ea89bb45c6e4ff83cb45effec5c56cac04740cdcecf01d03815457a55119010733c87dfefd0e539a8178da466ccbbe5fd7cad72c030d61f1e31f761656dc72d40614e728df73cb788de1ea5b31ae033b23;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5827c0e46453816b7f9718a2096dedbcab16d6a17dc2fbf5510c5cc1c007ef88ff8324632cbd4dbc32f11c8dfd0502a157399c0640a43b6489021f2096547d71a46402df57b41451110daf1b8df1637b14bf24685d8ea9ee4679bac3e662f0e67352f1dd86fb39ebe6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bf8fce8c2b970f8231578a02c8bfc68fa1b163bd91380432b1770df0a6dbcdd19cbd1fe85c55c286918c899797ae3f9e32e06df41bcf9bd4e7e16edd2fb770eab45fd39b5bc6fce7b1781d0f63bfefe5513883df81601ad796eb2cbba241f5071fd7ff3ff3799872dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1690e4077c59dfdb8235ec4d4c677c6197274ee89fd311f50033e9dcc5efe547649e98c7e0bc50e66c1852b669e34f577b5be3e2a2a7d325179b4ad8ba410803b2b6ef3d2aca2dd061c1a7554b4835f19bf62dc453095a48a42bb16470ef65d819845aee03208bfcf1e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d067d19fd10715589e6cbad77ae33007fcdd4e2acb37dfb576310e49459f61d8bae34ded9e833c90a2372c2b18a529eff3667538cb8f011461058cd6f9871d55994f5f3fbd0dd4f76895cfdee3330bc4d4043c57bab6a04321b071da520ee00a7a801fe81cd7efa698;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8d8fa31ed4a445b9d89a7010c1fcb0deb46ea56086249692596734285f585ad0f9d05c51817824530cd1e2b00c1728b89cd0d74322141a45c9df35638a07b84f6f9001a14a23947bcdae16bada3a3e372e3c3fc05947839cffc588e17533b996421b27eba8cde2f91;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h56e3b1d15792e4f572ced6d62af94f13e73d53f011400d33cfbf59f93cbf2d1b9b9244969a8fa67617c5bc72f1fbfc41b89ae7044fb8a18dff0e7257f56337cfae639b4bb446d092e94a617ce7b7b6632ba8a66e7ec304acd05520cede3f542cc05d4ed139e2f34797;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b90e4cd4710c0b25b781e8871a33ab7062e59aaef11259ce0b8d62d6528a234fb6a05e46db3ff5bc8c51ddc21efd2e06f286738e0f445269e9fbfc8edd1e0ca548c6b2ccc7579706527a727637d853a68f30084e9259c235e9b1424e2a73f729c39424689c112a913;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b61dd5abe9fafdd3fa222e9d92282b0b9f308c4c1d822acd408be447a07030bd7d95c9591056dc513e72cbbc7f12b68995c3b77bdb7528f6bb99e584e81f5e8515663a961d537f5eac13a25bb3ebaea69c7f10de71204a0a0faa7fed1f27c5f1e48a267bca968e7424;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1365ccded463249995169ebc2d588060fe3f3381788dbc4757ab2dbb1abe3aefaa314f06ccc1b076e7dafd71d2098f5d216d4ebdba1709491d82eff1dde246844004c0c847989c4ebf437b164de23074a73860c29de47f527304ad70db239f62411e1cd8712008406d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14e530e46d88c804f8102e1c64394366cb56a426c2dec511dec34a4a4a30f1fdbe6459d2f1fc6e19a4012cc25a574ff0468ca4e6afabb50aff171b0dab9dd8328318daf87fb76a03b7e43de9447a9237fea11a8761fbf234004c7d7c2b78d561794777c3dabdc966adb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16df6d875e8ab7f19d4fbc2f93f12e29e4ef911ee723e929f9663329f581dac41981ca665115de8bfc9bb38d8aca09072fc90ff7a5763d2df31bd620c083a0b01a00681d7219b2a80fb14a28b1044aa51f12dfb8708abc7d7ace10a682fb9917d20d5b2a05f7c241c14;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f1d50a5867940429522b8b856da07b235f72d7e06fefb23c65ab4503259b4c82bd4921e6cf2606920dfd1f040d64b9ef80a4c2f8972ee5f09b3f8ab7cb961fd2d9bde19930f8c4311d45297f94f71d20788c1983bae5018fee488954f4fe4ee4140bbc6efd242e3c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he990c4de700cba62bd1d9b7b567996a4db2041a54e7d121a0dddbe9e25c9f943eb49bc6abd002f5cf3776e121a6ecc2e81258206cd6c1325880276a2a15f74d8cab91cb8109c1f71d6dc1530b2dcd76185d55398e0d17346a306e51b91ab53e09e2a62280c7a63e13a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he959158b06a04c94679f953113e6a3de967788bb946b6575b8ccaa6144e1d4b30e2ae43aceeea21c642b51e68da1dddf1000c36cf192d725ed47525e2a4b82e2ead24fb6093898a0ccda9e94af1d6281ebcad97a8895aec245abab092c588d395bb5827dd710c12597;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba111289778cb4345d9dca021452c57f39926e1356590da9b48ec908d1d53849cc634e25a63b8ad1179f2c284a1237847edfac6e06ac7d40abe4af471121dd4c3bf3a5c3d0ff1e52b90396a84d04f456a65e602aae7af0a42d4f2eb1e0373edd270fc1e9ef23252ccf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc1311c4fd9eb96afce358d99e6d6361c540a61135445d880d5150f6c83e48853b43b7c624a15d589433c3e7ca85994cc17cfb50c943f75532a2a2d6fd8819c5d0231c6caff036f5796d9765c288702585fbe99724c2a0b26b538974d9148f8bdbd2687a514f64a6921;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d99004e27e7301e2c02114d32b11956e86549092930875672842b2097231d602283dc4ffe1eaabaf63fdd9b6437dc279d54381662c0aab7ade1d1f9b1b9931c186d97e0a9087770bc0edb84cfca7c2729173da52e0a71749385b2d09d8d0832802499602848c48767e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a0cff25c64d54b36ce982588d0b7fd2694d052ae60b90cb618188b590df028d85d94b8c0db8799105359e0b3bdf259faf3f693fdcb722618c1f2e908d16d4a432438dbbc0ed40929e1d5badbd0d9e6a5925a23c93569696846c0480d25f7b29b98988ebe8083681f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc71bbf3e3094b503a33d7e1de6fc6801389aa62b7f57d49778a7389f12844ac851da232241f0de418aa9a565114a903858c620885cddbd1e272c2451a44e083109a07026b27c7c0da1f0cdb787cc89d2329fd661c3897ea77371bb65eebc67039588f7c63fe8ea36f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6a2c95e95d352aa1861b56b0cc442a174d0d974d3309310044ce317ede4e3fa768296a10fbec1159a677f8d20211f54e686c61108e475f574574125e54641e7d78a5751f5c9ea7623da6926f2cb8cb59fd4149b75d9de2c77e6c0fb29ab16ee5e62cb266d62fbd51c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16aa3dac3ea4457aa1c217172e779d93be3bad8630028d50c08904eb0cd276e35db09c5876131160c76bb18827a00b529b15c9aead913902b160006812e6250f80459fe6d6a3e97aa82dc8624129c3ea2e4a2a7349b65d836b1b3525c3bff08c48fb7938a121cc9ad6f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197074227407fadc0d71ffbd3cff7ca9fc88e8304ef996f7e536291ee3cfeae233c0e0e53b18be0f0d2c4109bf734867c9a692b10a69a1a6336d5489fe170915b3253e3c53a96a9ad1c98be16c30b5e07a4d25ead0f7ff8d1b75d4385f3b1db167cdfe57061298f22c5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf0c449d6db6e5150e8aae4391799e363796129b2e3c76526e0a1566f3d2684a2f5ed567f29bba77ba9491634c3301c98b59a0fb5ebccb7a4a588c771a8fe63cc4863f28b4cbfa3b9d54e291c9f93df5557d47a3a13804a31b0a462d9d9e933bc540343eb9fde530233;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h83c8200216ae866289eeb3ef24fa10b385c441563b665efbb87376f0b6998a87ab0fa022f330ed6b208f17134dc664e28ddf3949a429556ca29915540be4c7689d9ff2870851027f73c152b47c3d727df6776eaaad81a19d9f0b0c26196bcb08164ae959aa29c76f81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113b3b026e782114de2020256eeda123077c0d98a84dd72d8d215cd630c7a42c25e71584adbdd1c5a26d80a4e9fbef6bbc84d001a4aa2650b2451b81670de5531d0eb713d359801899b207b29831552fc6cded226b98e3a1be9ec4f0d34a3d2db824dcd6a0103aebc1d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h422dfe3be2af4ef6f98ec9b682110fdc60b2df7738baf5fbe03ae0a12a474e1c6785af01ffd35247890df26962f47b4592eda3f51d660ccf1f45e0675b57d5831177f42479289dc8ab97b3fa88dcc9eb13746d9546767c6d988f21bb3b9d099751db65575ea1f159e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he66bfc3b0d0005346b016966dc16086992bddc6221f08165796d2e55d033b6fae84ae73db2279101d89d1d58b89e7413816cc6cae4bdd61b02ace397fd1a4363711960c33ab8a6caa594422b08c43aec7f02fc24e34ab895d7ff3be3a0829e3a1261fcdc4cd2fef67b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb8dd99badc1066fdf712e5c78747a9060c3d5f48623a8ad983b72192376a5a3e66b1759907e6e0421ba5f6f4fc8b43c1ebf343891625ad1eb854b6c13ee522598c83da584cccc45eefa0110e9f55b1d4057fa929b2913b548fdf2302e63965745053b9ac206e153f39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef62585226c9c6d1285b0fd87799c5344fc5a500a37da320301ac1760840d14cd2e17db433f796365563c260cdc66a3ed243be2c0155c31e6dabb8454386ffcc702777a6ba70bc7d0a31943432e05f228d214103a36daf4b4048efa8aa232eeec02b50b3fd73289797;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6a9ae490796a2fbc21ecdfeabbcd6853653351abc49c0b30e32d21b96f889934a9e24527afe03737f3371d7a28dc67a79759b36ea6bc3621a0bc43e80d6e0646bc882521d04ea2c9de37175b60a269fab2f999b69f018f688dfdf822e104f384aea14a958a9c4d586;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hac9aba1b51b2530fc386660e14c7559d76ca5451a5ba0a0b4ba3beb685ef184d617872e8c1618f64ea91f2e51b8f6f909d8ebfc12bdd6b3c11932fa16bf27602cdaa49ebfc853e914047ca97d8477a0ea171e96bf604496edb80a6e389fe2b0ec09f8150fc07209d8a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h935b9281adf3896912d8573a9f935d08843c77ca3af5cfd4550cbc300e9b5e89e6028b2806334056a14c07eff31ce9280a7ccb1ead7cbb9a8dd08cbffacc93844f829d9aeec408620bf89adbe2ac3ddad049fe515ae6afd654ce40c3382f5ec510bd61c2f9e028d99c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7dce6cedc31c6913a00b2008e044ff7cc9936e2bbd03a6e06ccf7c91b18f300c480993f53fbc9904a9790a9109b2ca5d161387a9fc25c7faef7b3172e4007bd435ddeea16c8a8107e2ec607c4b29df0ff43da75c1faf10b17aa895100b601046a0b6a6a518486f1ab6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c17f4c929fe0a8fd682ef231a4475425390c523fd912f1d87aa563b00d044e58a2c49929970acde70353085cf749266df7aa4f30b962110f34c4a16ba0c2ba74556f8fc78bf8348729693ff5b2897815bb9036355d3c7a22060038826563ea4bcd10813f3e019a50cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f09de2ec7529e562750db7852b1561d4fc700fdc29822357b493d223603e94ffb3dc25a4494fefc5cf03a351d88d1d28e6fe1f104176e14dc487f69ffc85d3f86176169ac23edf1841c093b04e23896e16f0595dce708787d86699725024a8c5a544aad9951e572fb3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54ce0d5e3f6b24725c552fef61ee296a05c5545ee3610105a82a9e22336772a07f7d809dd153816af2d5be93987363e4a76fdfb450b8f064491d73952500f1f247b5528f1f1799d7791cf386884d330bd9cc6096abb3e1b1386c2959406a03a1fb5ec8fb6c6e1b5c70;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19a9134fd0ac20e1afba88d8a07591278172c180e756ef7e47d0ad97847660eb7c39e023bcb22ddb6249d4c07e368832eca7b1c135428d657ca258e40d1dfdfb7c6b02036c90fcf8b0c5622a0bccb79ae120e0aec58fbdeaa3cd8ec428911ee37dd631464409f9c93e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13a03239f5b0cf454d99c75815298e5e66113d42e3bb9ff79e7eb2f6de4646ffb62628c4bfcd95606e124f26e70cfcb0a6421115417af9a15038fd4c4a0d42ca241d4074a80f8cd9eb2bc62f7eef07dcbea3c7bf5f000010bba746c8d9290ac04e56f73eab3880be016;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b9995f102b9aa432df3219794f8a4ae7d0ee249709cda6011c1dd498d99f2c90e396dc9cfe080889ec42b8bb4a8a44414ad22a4411895093f660c46e0f686bacebec887b1c26832da404afe3023caaedc5e5ef9ef59bd85b5df615871c1e48b4d656b5d0e5d8a2f463;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113bcf34154fe8e33cb88e7a9af1f2bbc154db5cd3288bffea31bf43fc82ae45f8a798e167b58336e21bc52b5b4112b536b53de0e7657950d5ab20191fb02ca67d7849453ab8fe6cb8e92afb535e73cf0555303ed692aafe9339c3b9d7739f379921bc0abda8ac2e026;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eb4e57fbacb43671e2facfc7098f36f4817c9e18788a978fcbc2ec427ac61277099b3a9c6f7ef5065b758c9cc9ad4d1efe5ff44cbc54cb48f24a199f282f2ba10d30f2c9c74c5efade5a78ad51fc8fee315af9b333ea5a5fbfaffee76b8bc2fef3ec9a2ab65c8f9cc1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd94527224c512b94da994f823a2620be5dee6bc0d01a58d8d705d3868bddd280943826136c5f7b26be01a5edceb5b431f7a0b6e145c63b3a9e20c337135fa544cafc97d68687e9088f996ef331d696fb0bd757d5a0431ac435e30ca97a4cea9fcd5882a8c1eba44bfa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165d515a79ba791e3dee7076cacc3b531db61a9a3f7c7f79daf32f2f05dcee3ea62ceadc37429fa558e132f5d716993fefe7eec5045e2bf3b2be1123d3332d05ac1ed29fb2b5de02d833b18f0ea1c3d2e35c4ed73fa48dccdba545537cf0de058e89c87df490b477d46;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cc2826857539d90ac522e14e343e43c3e9cf8ac9793a370ac10454b346cc17a3d5b14bd2adf0c7944a0cdb5360f21d1ab1a4e6358a181569fa33c8a0af0b68ec344123715d533c17f1571794378b958778c9b2df32f88d0a04a89e28dafab00492bc75659030e6697a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e71d655566d8a255ae4c1c18d3d84f82bc53a6a6dbef03cd82fc710f936864ff6ff03d07f335988dc4d53ac6ba5c30c87006aa256ed0543e39909cb0f40a03229eb550cc8e6de956ff8561dfd7a911b30413642d6d420073499fbbccec187b29852571a4f66bbb9279;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ee32c7b2a46a5dc0e941e77fa0bc0199808c1227c10e397c669860c7a6c3878704a61c6640cef8320c58f9400baaa3dc8f4d9b6afd86289818aed85f400d76fd169a5395fcf2cbd7bf468d552e2c4fa5148332749310aea058cfa5170a3f16c13d94e81ed2d660651;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd586bc9fca9ec8d063ecb6dc65db51864e95f619b41823fed69949a156dfaa16c0e1a81199de53d42986a13cccb46e2442b4b931ba55834eee64de525f8a4ae943d0d7071dd6cabd3381d53d289a93cef3058351f404b0a4ea7a0d920a0d4e2cc49ed03a8bc0589d8f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a61dafd9b2bdd59735e66999a582d77edee3a9e26c8b1f27494c40c59ba3799120c08297c8ff8759b442a3166c2e8cf2e3f89dbf7e638d55d7bb6a4c3e7f8bcf1046c23316f47865ee160a885eb63e8a5fe6c6728f29c8af4341e0348d2f60903a3d0f5f8a0db2f62d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b012d324b136ab4008951f57487672ba9f7153c2c704fff2d6207a43b6e44ce57371b3f0462b7898b5b6c855885eb9c4df9652561a1c19a4da7ad68a91b4229fcee60cef0e6b160ab0fa7d24f5ac3976fc97070abe8bbb20026a29ab727cd41e49b737db2a6f891a29;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hec696c863e1935495b76ae4031534533195b9b915081b32a48fe754e44c3fc730f683d3b201fa855f13e3de32a40a6b1d2751aeed5368b115c87f1288afd8cda2c516f1aa2a793323e30fb63682d1d80ca806206ed60f4b0a5ff91715bafb428a2bfe8ca136dd0e7c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1457a3b95afba8de2c8df458fec56a3be075a84c134599bc356ba3cc40cea80b65c4d3bdffa83b2ee2fd997eab2139bd03cb7fac5da85ad361a34f151a36233842fe63902699075e9f76f9228c48c8478cc866ae0aab9f37ff55e041f8fbf940850f932ed172a5ad9fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10076930e905b809913704afc0301f3e8b16a38810a4cb3127a00f02f3ef1a8a44f2228c5006d6a7aa978b652e1b9e41e4dfc4c86e9590a529327bc95f6fb2eb7495e644e80f648849406b82b9c7608dba110743c48b1918f015e1502f8ada383421256f8c50e49ed3a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12053d11ddd2c90ea6211464f7ac2c96fd15856dad4d46e1ee034bd0e961618c6a128fb7ab931504c2c9e5a5e16cd5652388eb2fb28781cf298bdf42cd8d2c3002e8a6d120629d2fa61ee164a22f0fb71eb1420db17fb48cd79b3a085fe8f69465d1e1bc252081a49d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191536f055cd6c3ebea1e23be8e188dee2799055e1161bdd280a0fb38d55e1ddbb804749d7bfa98074e503b118e4c89b6225c632c36d4df656c65f656ce45fac1396e78f62ddeb5f1b7ef587754c1cbb91ba088d3ee2c68d941028544bfaf2da72cf22524f998cae720;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb120be7e7be4bb17914cb1bef94765d373270610cd857d29245a585996313bc58faa23dc86e63a0fbdd4c6edab35458b5a22e1154011925f7fa22085663033e7dd7a8e2f97ecc9a6d6761564939e921d6ea1a931677c35d7443e04cc04726f998a05443e98f9a7face;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba8b0d361f28246756db037001c6072b818c598a1a6c43d3f3a3714ed3f7f06b9488781003c2651579c8f86c0048cc0d6fee71d07634f7e6a4b349458cd3fe4568501cacce182fb946ffc2d308573648ae781672371195818da6b8e6c7e3a3ca530adbb444a94b41ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e863d89413a1aea5553d4c3ad6dcfb7dab689c638f3b45ba51714fe504842f5a34c26d6f641387b24fb279addc02d1ea400dbbe27d124ae58f89aece247e100e3c5d25689f25deb741e7342a34e1b6a72085e298d21f20c4c499ac8dc2b5d9a83736151948714646ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha99994ede0a12006f13ce5bfabac58f2052e3378c0869a66a27075aa25b8d126d70da0093f8c467aad88fdb2313b8abcc0a4323a46b713afa70ab0ac0d60fc0486b51ba9742db9074d707f4f667a7e9ba4e79a3003194d444bfeb9cdf6d6b129b6b61df807431bb293;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e882d7deaaeebe935b092d9c3c39641a1c2d0c14417a2439db47c41cbb6198aa2270d37b6a9f8652e6dcd8748a95e4d53fcbcb0bcdf296a6da853a376c6b3b4544670516c2c1fad76a7c52ad52987044e00787d3f75e846c09ced8cbc99b3c569a27e162b747db0ce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15113277621fd0adc6966f38e81007fa56d126ad8bed8d794f9d7cde70f0817f88929a61cadc1c8c02edbfab8b0566218f7f295243f1281afa280ca328a9eba4fb8c48becdb5c58e235525a4a3e13ea3924cb292b695d4f3d58c37640c1d3327b454a7018586d41d74f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hef26d83a8bf1b3599f22577ab465d662bcf797ef829d2b2b1e1544645abe28e1dd8b30018f046d6d87ef5f90eddf2e0daf877b9c8a99ab979384cc612a94bb6ec552a4583179c13ef7a0c3157937df54bea4929381148797e3eaaab65ee1b534e9f69f271a76e2928b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h20dbf428f129e9cb66dc6994ce716b627aa076b5d2ce01444bb5d167eb38418e5664fab186d550e951d5300070222effa31a0483b4ded597e6da4c1f648cddd6733603b4c3d30fcfb67b1649dccad43de555f3d0d3bc7b237945ac2335fa94da3dee64199ae82b4f59;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3e3f7f34ad7b6e3b4f9fb29b5a7c4a9383a9a4dab19b9f33cf00b31938d3c34532ce8c940c6034469bd8854ff3751bc369d23325535891f470bb5019ad5616cbdb87fec084c6f5c7f7d12429ec0d5b51fc92571a821f945b39fcf001a5f97227e0e9c19dd40c96eb2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad9a14d87571e8d2f0a34d7207cc135c32687ea840611099fc8f81b0d04323f036c65782ce060977441828ef6f44fc83a5fa187a12840d968ddb23f4cb705df8af690927c87b512bf45e0f169b462c819aad7e8391815807590a2ae93b745877a8a123e137d3bc75f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1523c58b3e83d336e756b19abf166ee593fc3dcc90438589ddeae8dcadeae007174e4a377ba27f4d8302238dc3e51560429b74dca42b5f8ca0a7470e6740f76d7852baf9f139154cb44bacd1a56c68b226427a8a6835587ee387e7ccd10d2431ccd05efdad152e3797a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1480757249e771f4cb482fb43c7d80ab0bbb8030478ea081c0201a210dd240d15f3d836a1034d8bf04bbdecf363ddf406953f01df64644a3e212bfe4cd61f6ef45b7b4423512c28d74df7dd2338c5bf104e20a1302ef50167f0236a8ca845b18b82c163a2b455ac3d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a83eae2830105830d4a6710b4b7c375e9a50111a3f1a8948381838f4e9e87f87680c3c2bebf061df4be1e1ddb818cf83903a2d66139d913a8be8551fcbf2a298b9af698195a625a7fd7391699791e32c3677d1630ac95abab099438d01c3b5328350e346d2c7af735d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bd4c23a3ab85e24ff259746031d6d28ef4477f02c5771d2c4a5d9cba50e10e3c07ae782571dd4882ba4bb70cda0b083f15dd2ee527af5f5b3629ce128ba9660b32517e45dfc98e4f46ee9130b193ecb1bc02a9c9d0d65610565615b7f3a5404cc4fd652a4a49b8c7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2ef461e44e607e7b3ad8f6ef263783c459994fd08722d4b1252b8778230b9efca19e95b3f3fe46457afa04ea277456f8326e2ce6a3dd611179f8b06e51d812de791c08e3628e982084e67b494ef94ba4a6c71f1c24b707a2bc0f718095497d87b2baa76024c6d587e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1df128c86a0e9acb735004c076dc3f436cca9b97c8270197700398193c2afd5bec354a50cdfa95c4fc87f5aa78dd9ce2222924708d067464799f53ddba4ed3fe9f994f5098517565eb417dc9481ccea7049b98a345d29953c2b0b8f07adab04f787ae6f5a6cdb0b69f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aedc46a9a6cc8f74b8ae9c980722ca099aefa1b392507f51b8091d1f69154816299f48717ccd58810c5129ae13def4f0fc457f7ee5734476ee1c1ea0aea1761eef57aabea6aa80daccb3f19734b2b2631ce735434f85c412294eaa1bbc207fd85e6b32337097f46887;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd1e3f8466eabde301b464fd80783d385ff5aaa2c7e227a926a64924b3cbf82b8e5177ed42b6d853c4838ab00a45c0fb338dc7b81da67d84cf41d2fc9c2d34b0b130727c5724c5d38f8989ecc02b572b108ba7126f05d8195e40a7a0846dd37b097a1b9d5309b1ba839;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb39a384711cc3b07c439ca035f30ec4bf4d29dd66b182a71009f7d3898aebf280081a4397e0c40d3ac6df880eb141f4d59e5aecc764327ddb723b822618705d9f1f4381b339b075032786ddb34d7d5211a9d2a6a6350bd3852950cddb2a4a56efcf68983c26c2e09e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8240ac25405922cd283b6d5e6364aa91c0b1a143ecc154a60513029b077918b264bd332a05adfaf269299b0348b72ba3aedb5db541b981fb42f567b1ea2181464c002aa510447d5f291bc1340b4dce3ef3c16bc35a749effc21d6a4f236558f43da154168b7ef4f9da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he9093c0dc62d090996785a5cbd3491bc6d0ae1e6e8ddaf66859f4da9933a98d5a154126bf4be5e07eb30ab83ce8b4a7644b525efb9e8a49d32d2035093b3ad5a5496343902af8d51af9bbc67a7465f48623fe7e3081cd00e2ea13f11127f1fa507fd87de9f3da75a9d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h189e821f4eef70984fc2e89a8a97393e1b1a28ef092a532d216012393197726a0fed7a30e40fada99a7fd09703e4677a93f68c1a766e548564b66b96a338ea6d1b2d7df8a081bbb0b9c133ef32cb7933b3e8801c49ae3f066973d129c719f390e3185b62c6373df5e47;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he36865182f68b8936797915e339ce7c17231b87a0b2765c2267989763ba1f36e3794902fdf88217f94ae9e51328ba11df64ac54f87af5795afe67f8d6456c8b510c8cfa758e8d626bdca223d3f9750b450b4955545db6a79d6fe53fe77f6db18dbf47913716155d672;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hded54c7d4194248246b0f221083b6f5190270d7af3ee37a9aa66977d937fac2d483e5242c5690973613f93865946c4701615936e2ebb2224fffca45d700124ef8db5b70b360d184d81287d0d11f74b1d82f029272feecf3554e29b369463bded5f16034bbf697af4ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e9dcd589f2b3be7ad633b230d60100ed24b8254bfc1054dec61ba409cee3168eb056779d4232731df5fc22bf9b53ea0159d9575eb4884041dae0d19b2d9a8811c7b17915d1816deb94457627d87d36759a85b255b7f21a1adadd8b071e3a0bd652295dfa2950bfd63;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h364f2f02beddefe6c844160f741d00eec0f43bbcb2798414ce3bfef9277b33de86b9635d0d355fae002e6ff8e120bff58d7e7d80fef5b307514e75de3f7d676f0b12beb9e06c8210e366b24ea1045699e7321d71cdf68c0a2b483a9a3a4e3ac1322041564fe4fd5646;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e89288e89d0888507360e73be810f90f99a053518e991aa6f3d6f4dd1ae0ebdb79353e0ad3374b6921a57b0ebf36497fc01dafad7f5f640d10adca6e5173402045816ef966602e51e3bcbd90e97243ece4eae265c693a5b1b773fb5cca9fa7d6f2e508e10179fa080;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd5a0613db222d6f41f9d9e789a1c64762f9af0d04c8d748d496504126cf368dd7f519c4333d64338498be571d6ea43f490509df484e67eb6e9150f97488219cc340221906b752ab47c1f20f520005ff47afbe8fc074cac100e23e3f728b18cb0e7b0a3227c6e9f72b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f99f67a533ff8a798d6e520103f9e20b7390c0f91a9cda588d12c540d9487c676f56b5fe29576626430d431caec532a62c09d663f433a6ea703d148f7fda2007a2beef82c378f67f621ae198d56114d309b612058e4f258066372e08c29cade8bc89f5dd97f1f97413;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b59abbe4b862446ce3c421b7cb7890baef1767409ce45ad165827007f765bf17d403b3903616de6447ec809c343ebbb2254f5f0317e11e2fded828e76966e1b66ca6e912ce321b7a20076eb5ab3f4424343aafd9e8852d8b392db98f641d5952d645a0b4a01d794ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had8a6b5063a75bc520cef3cc5492cad06067ffecc166d5ba966b35b8f558789c962b065b549a1d9482dc4bd15c9db59389e076be137cf88d22288e347900970e8dbae0e9fcf288cd60bb791b19b66cfec423a0671a1d7afd318dce22e0d56b4d5664abd4ac6ef4618f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12455b7bd1d1a578c9ca75a89f51f615930933d8b5f1be7b63ebf9a2f2c5a53c3218259ed55503f949e6b324bb33672d371c0f1ea14d1212ea52a67ee41c2030f5d6ca1e9666012afd1a137d8e281c45577e7c80d36b7c7bf2ab25430cb479d6624da1fafcc57fcc5a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd29a8ade962bba6d1f6af4538d6f02e57db6a2bbc6f4df62369520d4e6b0e93efeeb8b1f003b930b6664e4e7ab48fdab6f27af4d2e4509635fff810e7daa2b66149166ec8872efba65c03b65debbbdedd0ef350fc36808436b4cd0fb721cb3e224ca912092cfe9784;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8ae686a8c61572ab611d1a06bd54c048989f5c295b1ca52b0150fac7100bc16ec102e4cabc7c29175f0a39c14c60deaa9d3735d45b7fabdabca778637a8afd20de3607ac98447d6cf4383d0f3ac3fa037a9237714a3b0d437c60977229b2c0c7a63c4bd0c7e542c8e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc40e68ece60742beb116fca5f0a1f25b5c374bcb9841335cb9af724b2cdc0345154422123fb7cb9afd5f9d8f49fa3f19ea417a703345fd000ababe032cc6ee90da607a2a7c2ad8411e4278be024b6127d9b69a93324fcde4b678110fd66e4b89e34d582f1ac5aff21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h92d3c3a24a5e6631708a5b08d483672df0beac913a975f15854f90507a6049389b949ba6db54aaf7180f6f1a67129e7b5a4cb98582876e4b565f4831387501d8f72ce128ea152aa5e2c7f8b9aa6c04af876099badb88fa10e649499b8f4deb0896e4527643f64df5f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1223443f26eae9ca785d262531c64f312fc6a09abb15e56c140bcb8594df2b7d53be7bdb667c524f2e15df6dd7e11802d2843aab8c30432ca6888642a8f9580927ac54b8e3d139a32c0a74dd96dc8058afef96a28de6c00c61607e19d5125fe62979a3e4adc7a85b96c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h38539ae136156fc0c47f50966c8515dbac96a895dabebdd34a90151fe4256e84e24ab748f41ec993438647c367c70540c1618906f8fdb5ddfaa13a3c36b9920db8d5cd75e6b4f460947caf92f269d6e204687249bfe475d8d74192ddc083ebcd9d4657e8c8f4e5afb5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ab60fc84894beccf7597674f072df0e2216f504b15bb42c7a072b05dbac5d33e44eeae47fb3e59622adffd7f9cd0a9359cb5e97673b1b5c4152b46556adeaf94fd2f1a2812aa637644254f41f0b758048c2c88448adbfcce8945ce284e75ca86da3c55cb5bb1a3a12;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf50f71dbd61749332c9c1a0af307d57515a090814597dbeaff46f1cfbe467f4b6709bf76bed00271fde9e4f030449182c2790b3922ee18ae086b1d021cc0f9211570e116f2a2fad83ecd19543577cf875a9994f4a0ccc648bcb3be69837c863dc1d3c6b26a3b6d02b2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hca369ff5d4ec010ac5a3de3b9f17fe4843f6e46351aa76749b5f58bc98efe4fef4c5cd28f39d09f7af7c0dfa4e7e886d5bbc78a43cdb2bd98cf5c387a8cf673ace76f6eca0241ca80efcd0e40d7f1e4aae7acd0c0727d96362e06996e2cfcccd62cc911cc1541799e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17611cdc51e561425c3532465f30a958316de13dcd83575309f5a6dd5b2607e2780b9eae1c9dace4f15a9be01e2fdc8de1790f8740ad2039bd636798bdaf31327aa9c5bb909ff6a5c2227f07b5c99184e8188729be840ddd6ce278f062bae6fab50ba2e9551d108db40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15c69f5db26e2a251214f8de43be307994b794fd264e05882d112c499bb33b14694608cb5643cc0ebce928bc8e1e070e437d190c860c43f18c030bbe7ac97cfa351936366f42dd40e826b28d3a6ed6b5d06b500ca52b46baa055d030cbed5421127937c53b31401ddc7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10e3d912bceae25d95c42bb418b6d10dae7529cace849cdb0a87d61cfde5caf60b1a9198defada5c791b129070017b4a5173851b57a774ff765ac7b98535a54c70eb70767a0b5d5ab953343256447f35e2f6529711c3d639c8235f9e902a2fd24a94b1caf543a143b0d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12704b63151e95fa1eed63fd0aa237ba78ea434b53d3d2358c499c4c4375f9c224a98dcc07637b8bb833fa759614fb8259c69e84b684d9af98935c03a1ee93b2a681bca8bbbdaf153e70a023a93be1620f27bbe744528010c7a3cbbea4bc5da8875785341c5c255745;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b241eb8b26de79c61f5932a08cd058a17c6e7c44e40fe7d35f58af0dce822dc1e00f3209fca3dbe4403d2190a2d51953d30223ca9d06793a5fe145f3fc7036a31876355056096959558fa22e838ad5197fec19edac9b6437e57525d05c7b93e3b957dc8cb4574f43b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ecb5e0a391b4ccf19ea3d0602bfc9a7fc7e14c684940f7c35a2910a877d12d21bafde5c9ad67556f2add0ccc089a36d488e998ea9334d865573ec8a44bac9398b068571d36858469c0e1cd20c0228f4673c59a69d93881ec434b126e28c090efe0cb33f5f9a33f8ffb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108ff9f8b6ec85590ee4fc0879d12fba5b77e15d0727f69a8b894cd36d0fdf13df64686256df110b7e54f275e562d54d3254f82ebbc8353ca32bd682d5083f7470425df3ac5d0b1fce09403f00a1245c9a33b87d357ad3c68e298b01657febfc9aba86fee5fd8730145;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58ad8ae958e898ddd86b0c1e9946a9b91534a9f9efd46965299eac9fa3bc11c8bd49a83acb822b737675ec8aa2be11a5acfc6cb57b52fe1dcaa1cd7681ef9a236f3b5c9ee4c000c6c32cc198dc0fe0437d12c2b6dabcb8bccf703f8a6a74ec78c497b8287164b03a1f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc4e2faf0eb0eb64820706a38945b830b28aa4995cc9ee6d2baaddcb47f51754654ff13b533acd8377fca1fe696b9f4db9a244c701ae9a9b30de75aeb0d122361be871739f4124df65afcabca48ffaabb9398902640ba8a6e7c428ccdf7ac9dc9a561b7fb309eac16e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122b641fdc065256e14f72b6b57d1f91f7855d3e3f76d90684a8551e8795f5f3b9be371e8ca76699d896e95cc4c918a848473337fc06619996386854ff9a40ac3569dad74faa50403b21198bd2b0ad242983696b8ef52822159bd5cbcff69fe8166068077367fa7d3b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5b09feb556c9653d8a63e04b61991c9c565d1ea939ce9774d865085cc365abb2c156f56953ae5e65ef9988af086c635de816ccaaf0ff636b2f117fbf0735a21d4fe654364127d752ccae80026af09272af745888ba5c13c3d13741286580e7ed503edecf88d85c0f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e0ee272a3188adfef0ccfdceb113c025a379a0534fd534702abc7831f5051f81447de51e1d88ac9a2aba44ccf581ae5da9fc8a0e6aaa8467faf53adf42967ad219c5667a7412b16bd94a35eb34f8ea54de4d668f486257a2168874607a4bd7430dbfd64c0fab975f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb84ab10b98cde57565221b48d4844419cdb773d9b22426458489d475ad2dd1a323a586b802f05c071bb605b75a81897d7882363fe355f95e58bc2fc8c432620fd5745e0e8ba870d95f16824e8400d3f9eac73efbeb4002d292458dcfeba1c63c71ab451709292f27c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fb21ddf8e0155c9a920563c628585825e85a73b7c3d09a91864005beadbaa9afd35161bf5a6f78e4d76b21f03333d66fc2604f5ed1154d08b453d9a8026d182f7806e390a38912bb9a64c06d205232d33ddb0fb023491abfef83f5672f68355e2db5cdb0bba0617b6a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb90cdc849600a3f3f828e33f07e8ed6cac6b92a4ed9c6828d54b9b127acff835bf56d49e10c17d7b7add773283f9bfbe6f2ddd4aaaa4ae68fea8dee188db971c9417128f328920e1e17d764617a3993c701ad0697d3ec682ed4614bca24930d82a1d49c69f7213cec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e59a971be11eb4c1e43fd2019d8881a706a5565af467e3e6977c9df2801494985942bbef1ccca4a69b0c65cd73b069b8ee3864fe26a9406524efeee815cf9534f64e53530beef6e43be41d03e5ea998f000578e12c65482f682aacc7244ebf5dfdd321e6084d9710b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb9b981be66cf20ff7271cbaaf5073ff74d9bf32a4be91434902d3c4cb9cd85972fc9d9d052280d08c5b953fb41b70a795f07501364ad5cbb4eb36a470ae6f423c139a3bd2647ff498f38990940139b6674249913d17caaf237c3878cb899e772fb27a4f5a46eecf43;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h762113f1f5fabcec35789ea1577deb5c6e87fb6ac3ba2a3171939038bfe096828007c1773f2471699779304e58d1d4e57d6c8f44fd66c297c3be4bdbdeee00717c68f3a9de46ffe538ff946c274e3a8bcaf64a86a115c9a23a37023e2598a3c219a67ce47f0d9968ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d49ac8f78e1156577b53e6454405a90ebfa52d7d680cdcf8a840d4fcf0a16016b970e9ce20125aef24f0418c39d02f53b3a0c1ee5d33c10f87667823ac974609868549f71645c2dc00c08bc72cb306eef22faf63d74d3684f1331d303ca395bdff3890033c6e21b616;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90598b464b263c0b7bd9317d254c2154d960f0dae0d98d06bc951de9b6457b6d635b34b27db253be640a9e6bf78fd6ea59adcb9e6ff7b3bef388d1cc41e65f402ddea1e67a5efb3b2c6ea199918ff8af64e37d50eda1f722e127fe0d996408366754e03902b3fbd874;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14bfc83ade848ee59458425ffbfc802e80dc96d1153ab728e8e21e6cb777cf206251b2f812efac009ef3781f783941537a4105213ce83096fe839681bbb68bdf9bb69647776b5b34bc51ec5cb9e15cd088a189e681a30715837d8da66cdc56320797c57e644e1483544;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b7812e46f7eb0545510f80d0e6842ee240193765ab0137492062a20ea5e487e86c7c4a66a30419258644c9a02fe598683f6eeba3a2524da68f6e6696b168638be926557945ba8eef195a76de62f9ec49480cb9af2ef4dc4c4bc35926ff5f1beb5515f1b8ff1f3eed2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e23f05af3b7cc26dfc5dcedd266b72331c2709a4c187dba68c0e4a7a2a9944d382f8cfc4d04e1ef761152e72521d766c35fb6bbd58d2576271e238362d79070fd7b90267013c71e5a2ed758de952201910b61e497f90e3a289c65984fddbe347d2888d6655c489702;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd110f6afa6a90468884b48dac5c1fe1ee4bb0b47bcc216e24aabca40011f5fbde6c72eaa1883e26bbec586fc8c42639d8a99cec58a1e622fe5932467d11c037978ee58bd3d38e83b7806ddaf1a3c148fbfc06925561544df28b8324778749a6c39ec537039d4a1c4e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4286f0fe74d93c76c106883d509f1953d606ae2ba3b67a10a261138eb021159a05277c0622ed005605b6ac9c6c66a80d87e350a97b6deab64b0106e92b34c81dd371143bd4407932f343fd1c7e24c2868a17e077bb83e8a775d9f22b29cdbaee33237f5d45ff4ac0f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19661e785679e6a1dd4b4542a178df2a483b05a13be3528e845504e4e4a2623c8df318065ccdd5652743d26f86cdcdbbfc4bea7de5efb492410f075786fa618a79c7bde79afaf50676d84dc35502f8d2cf3204939ee76f11a07c0818d8042a8839660c516130ec574c3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcaf48f2598a00c77de526daa9ed02fa102a374478db9833a1a4b897948859baaa7999d1bfee860854b8f9c7c5cc662e9d88dac4f83f9384113c69b8b386ab7fb5d3cf91e14b73549ac1a7021958ed21c5d3f05ae961319f6404b49581fdab37fc8ad2cf6fbccf0717d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h355cbd7a5123c4769fe8de16f184d60ce3030b20a1e2f3fcce83e13d595ad81886f23629c3ca0d559c3a0527615fd06fc12e6b2d0915cc9a52b1a8c51e8bfa4b56b6aca75444e47ddfe7fc3bfecbfd9b76ecc95982bef0ca0f8350898ccf2efa50c1d16497e487b7e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h400750ce91082379d0935982a5a574128575308db8864be82d1b83583f10e3ca77d8a81300c68c39c2c99ab805cdd74ad1933614c088f0600309b7e170c597c8419a91dd5931d6f37e1a864a2a7b2eb6db2a21cbb5c1656deea1413db8bbd775b3a0e82658a4f9b642;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd13669207bb4d9b55c51ddd36453044606a2f3e9581132d38f78b0a9e42892d4c6453a4e8886b4c49387d4ed15cbb9a2bf3d833e5e6ee3cb30005db844836354cc67c4550c82f70d8c3b268e3268d461819a5deee5202aced96b70cda5adfaca16c48935b8b68fd04e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1103432c4d52f746ddac697c8fabba54a2c0acf3d2325b968e88a60ab645048edebeb8c00b81d17ad996ab822efff4953813662cff697217546c6c987b1b180597791f8cd98a09dce21825fbc4a57eec6435c9373abd2ec21bf2f37011240f8f2af6df3070eb7572755;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d69e6b91030bd7634b37551766eeb1d55a207e909f1d231c061ebc7716f2ecf3c87397ad12254560d464423eaea4dbfe282c7f5fb7fee79fd398e7c436ff42c122b591458c06b0985214f5406c0ea91b8256d9b8f03abf18ad73e73fb33c38f5466f02f7c663a7bf3a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h77a3498105a59124f145a1d97f36e3baebf5ac92c7fd3a93576be25a13b1aae64521cd108e1656ba0f966d0634245ace7cde13b903423f563d270cad4ad562db25d68b74df9cf92fb892470b25113843f75293b1c5ea2eddab36f41ab0f6e1b5d2e6b74c45e1b2fa7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdc03314c736616da54c3df51edb2f0903d61d0820d7c3ad9c59a42a2b045542ec14fcf34fa6172189b084efecf612e3c2e26fc4e34f6f74e69064f65f2c04e3cab9654a1a2f98df71cf1a5dec806759e54f8288a481649dff3b283adab1173b18e79acde388931b99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd97264865da5b6f2d39423d7ec53be698ecc433f485cdb7f931c047355cf1ffde8cbc3ca6a5fc548a9a79296aa4262f154b5f57cb0bc5c27dba51f7e3891ef8b1a1deabf051a031971da972b37e576af35edd72ed5b4277522c2e9e8ee55abf33a92aff77ff1fcd356;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d466af3c7acfdd37a93342da8633459d4a80bb81c2d56814fd4b01c9ab0ef47f6161474d024c4cbaa249d64241703ec30f5b026f38448a195452b211af518cd9b9e8baedbaba3274b7e15140697d83074516479631076f0cfa0f75b4dc3587f5f67c75a957caa1809a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a942e9507c69bdd40a2563cde3e31db3181e304ce29c9f13d01a85e8a16fea649e2ac2d7b6042fac4665d80c00924d234126ed16f89595dd547508f4dffbd40913e407c2fa6bd3a5366fec3f5cb4725725b11169cbed168207136d7cc9ae3d7def80020d015e7dd19;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb1c7b043dd43b1a7b3e02a222946f92f9c04e5edee53093cf49cce3e0afd44a2b1061178c2808b3ae56a15b3f3af2ea2ab0af59fed266c97c09b0c515c80f0b4da600f73529f636ad359e592c6f4c0f830199b887adc1a7449b3090fd81eddf2c64ebaf9890426d43;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf19d068fe8d7ad5e4389d66c03520ab08381f45220a2af2fe370e9c890b3169b8c76e8a315f0e1be2dc56fddf4805c72acccd77ffb3848124935343a18e3da9710f119a2a33e01fc1dfb93b6c8eab216980a73a127019012e23558d8acb6a134fdcbdfcb35c852bcdd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbde7e771f7f7c40aff8367e5794f0e078b353a29a0aa0e0ee2dd7bbe1fca31067699c2981754a6a3dd79ea06e7316950e2baee52164e6f715aef7fb0871e7cda74fa7ea4bbdf53edc9b0b801c79668889d28f61341f94b96d58dc2ec0a2f03f39fb29167e895b3505b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h880df8c9b943c53eb18bf04998b212ed46184174245a32ee1a177c15ebe546dae33d512f68c55458d537db5ba98872b0a6a831349378e7945c2657f3e0f14cf7deb4137a0bd5a212e1ca5da4a4647d2b5da98aa3e3fb9e8e70eb3404576e254910300697c867039ac3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17d9456f6bf03259be3dd9d6d88d694d86d8e44c3c08223e3cddea4b1a1d901c34226eccd29279e76ade40c9bc679cef52b20d0d27df8675717d9c9af73be6bef5c74d8561f4443503c6e596bd09df176dc52fe1da6ddac969242d07302285ded2a9e3ec2ba5443b7b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b1daa16fd2b6a512d15cc5e274d3db8fc6f62c96774159d0bf491fbb71b7414b34b792e37dfc713d6862fdfe10afdeace08951a5983d2d6378cf46d0d61cb4dd3d2318c9c5a433a9ff6d555c7bc0dd993470a714b61ee8214f0fa11da3e1064b14d37320f5c8e3abec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h89bb3aedc26b905b7737eb7578a21b5ec1bf6527a9a09b868e90b48fcec2613f3e71d2dc2d91b39b404466eb74c379d56fd96d42e9aadd2bf04b170b48e6c90c2519af4384965f12256f454fc6f60e9e51ca40702afe37901ce7fead361f3a5af1a23e8a2cb6117072;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75be39b197f02316099f32dd199ce5a233f8e011861b0e53605d4132fc03c65bb4cb032b924fb64ff1af26bd6bad7e8fa626f78f9018a9ab6143c0ede10ec2dcf0b6773a2d7e09bb2b3e4849da2fbd0e2681ef53d7ad8b69c2d08f152728676b8c2007c1ffa71241b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4f05869b6e7f83b45a837e75f47bf7d5d235abcc357274ebbfd03e3450279ad20c4b93b42697a860f90d1610150ec8cf66b4c70797f194906724cc228f9e1232b9f61947e3fae24246a38262041a54943e5bc8c9b4fd0f8ba9cec000633306efff12901a18c9aa079;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1df876c79413f881ffaa048a714b3180237ecef7249291009dafe6be0b60bd199991686b3f382aa70daf2622285dfd85b6b25fa6a3250da316ff2c43e9cd29313e8ca39a934f76069914a796e5eabe73fbd2e8caad37ce18ac9b0c040108bed2a6b19e1d10e26ff6d3d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f19d95f63185be8350c81f152667b7ddbe36b7216446e37d69c23614717271fa83671aac0b760994ec7104864e72efd6ac6b92cace2907f36be0e3a24d17afb18812723cdfd36d484013311089580bdb98ff367aaf238629cc6840bd2b10c72b679183e4d3367c232b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7654287127fd53ed1985e8732fc1f11b2e5fe24eaf3d3d5e9cb36c0f390058603d4d9cf686b2299b0ac942b2bec62f5b8ad77f16b8aa6106d7e0a748491738fb04ffff1439ff0f32dcd94c4ca60a858e9e4aff00cc8fc8a313372645bcc56e368402ce28df50564ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h129b2969e7c9a5d83aef7507e40c136b09a566028c85e0fcea16f472c69119206657cd52ddcdb4e0b4c36bd2210261186ce0e953b511e69394bfcfc6f023bc0569faaf5c0af530dd2284d997a9279431da7ffedc16381ff56bebe1281864419f0a2dd9011b2420dc49;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h113621915d6a3b59a53181fc337b10d07d0b583bded7030ef6ac809aadc3609649f341c87410fe30fd735add365b4eeb3a96cfb82757328a64926d1bbea86bc53f4d9616155c32912c38906c374818b4d6aaec0575debcbcecf3dab35c9328ce6c1d7b483ab5f053312;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha9e5217c0ab93465e382a73a93fd217933618cffdd867e4951f8385c9a95369b91331863db82b5cfc1a14d22bbb7a2dfb6021cc0b9e0d776f2e87eb69c296318d5f8c6afb0ba20ab1a66e74a9be4502019123595e35b2f7774cf68106019e9542d940fe6baf500ff56;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac91c5a2c4477e76d8bc5b00561bbbc2c1ec96e4a206cef61d98860210082c3b0e7282e79c2aabff9a1c05aa4bef398eaa4ebbfd3fa540c98382028dc2eb2a5b86e0e384c27fc1c6781d3d7177150b18338ad138e8c6a3eb15747f00fea09b65c0f5c1ca4202bba6a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb476f4794a1ad2a471db7462ff1be7122f5e20a5246f0cceb39d349084c2adedeb446968570a3ae0cf060ad6cd9f8bd1d56a8475e179d30ed5b011ea0acffc5e13988bc92fe338fc4afc069b3a556f8de6000694446fa36ac732d62c3e0fee0d1fe139a2fe210ebfa3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2df73bc67c5a382204d8935b120671e94a24d9a943cc888376330c45281d994d7564216a94543c9c418604021abeb410c1b71d58dcb554dcd54ad25d91e6212a77d4feb7a453f15662a85be2fbce075ed3b06b33fa0b6ab2e384dee078c66e8bfd13cdbf2361365622;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha78d68330c7cd5bb76570180a86c41321a86f786a40588257749be7de0e6ba554d47b16f9b8516caa27d220711e23d70852499d9e8dd4bcc3aa3256b0680acc13f4d6c84cf0665ae9b79149a26fe9ac9f1ed0bbac633a7126433b227995c37b134487e78cb1abeb5e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h583f43ddd4e38a4caaaa58b50f6dd892440200ae8ef117eea96f098b3588a9fb333966dcf22fac4c91d4f0271dbd447c99cceb1d418ef0fbae655a0f093cf488a84a4e6006562b6f783bf3e675bab24cf055ef8c1bb9358e13cc5942fe44194efcbdefa15014a47c2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c24dbc029aa5bd5fd4813282a1fe15d2886d10f28c66ab4dfe55fd5c4745a391fb71fe1deab76c27b96f5bcb7ad33094df173f9a9a61759435c54286979948205ec575e242d8b51efe23a8365249200e1aa7fbf4f1fe53ea2de5a31a4fc61968f9e089bb5a6c96e3fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e4a83209e3f1b3af0ad6e8d07a68a6a787a5a9ad3e69a18ea2a67142cea5b1f00e83d456856064a2527d32133bac94ba44f139ef5c0750e71fa0d6f8f4bc6f59764075fc78372eaf1759dc868a8ec8fe1fd18eae3d2536003d02dcd6ebb33ec9ce88628fce7cb0d16;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c866d4a81ee27f4a5e30d41f2547b489a82e6549da77421be1afbecf16f70b2065013b4f4ba1f4daee0f0cc77ddebe7514764cea912b1b3938998121b55044fa66025a581f21db5dab101da8722aa5652474a5d41a26135a33c06ece00d86853217b69c0c5ea5ed1a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15654d2c6e653ef32276166819cb31a3c96a691df73eaa5c9927133e2fca7277569d3836e8210e834ee0b1a9847111198eb04ab27c2adc257ba6bcceff0ced18cfa3b75367a5e7985622621c626d53b9518e9d2b1d668642c53c124f1c79d2931e027284fae7606c654;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff011ef9fb4d524d4b5943573a28fdcc2effbdcfadaa3da603628ce09666d50c4525f619ce09fbefd1eca25790ee6395af6926738e13ee30772457ead2efe1ff276d591c8e5813e48e9ae2d094e4d74c118ec52d309c835e9b2ae36ef73d73948f975517b3312cada9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c55ab344ec6c64c0ebefddcb550b416ef91e008d400d9e761bd8714199eba79d0347088fc65165c3ef082b8faa8706f3dc857f3b76d05d191cff4cbc63ca22addd19fea93d100b0854de33f51c4bdefe750842cee252919817e8bdd109c22e13e162963d6e6cd9f297;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e2b6ea9cd91a203d6b21509c4cf747ab74f5cb65711ced89b4a403549b76907eaf269420075c89013648cbfc2299a7da16c4ade5e6ddc408f90498e88aa56ad69242de63f2eeae88d4fc166417cb5013096610379606d90763598e3b5119bb676125474e743483b7d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba405508fd1286707fb8edb17192ec32465d2da6ac840a80ad6e9448043a9a4ddca091d8c0bf317e397713af99db95ef483952800a6f2fa3bfbd231c5f7685d5f60352a4db55593b6d636bf71082624fbb6e79303852e77f8bc55009e367aebca0e45b604eb987e410;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99c162b03dc7c64c94d7bfec19c4369fe0e58254c372d39aa53db9f463e1000e0219b126458a03bffe07de73484f496f5dc50631099f28c193610829642f307503586438fd7cad0e97e8768161ef1b5fca8a17c5351b71b15460549a04087f404823ded9dcd1769713;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11c962d67334648c270f2ade87cee2ce1a218931a219e88391aeff733163b399f5ad507f15161d814abc9228f365251a9fa32cf9d579392067fc271c06f6379be493ceb64747fd3a3db7a9dbca9d9fa0b068f7e7579ff2838e8703f10ca7777628365ba03525ba06a1e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h753d3afd8caff8c07f4c1b71c3e1e3ac72fd26146383362738b5259123605fcec39499695b06ac68f071c8fe8f863b66d6d5075406f43498996572ec740aebd8a1b79f7d7fa2255db28ffd083e04ed026a3ef7c7d4e511fbf4721463a2ba4c972776e29c27890d8ad3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h252fa0dbd410de4e4f5deb5aad3cda40000c8ef9ce747b95d8989af187fe5cf6d5527ff3f71997c3e6758997571ab706bb0ac7070bb8b03ce8eafdfcf472357e9aa6e2943113402ff191d9531d7f6c6627d6a5a3da9b0af164a71110e38578c5cc0c71b5ae38042333;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16600176b5099f39b3c38b27d38dd1894a7a51c7c0c86f07781749a6a8413377f7e4cee0ec885364d9351b070f236682eabdd3231cb43404dfe568f60fb935afb2dedaf01be6865f83269df52c1be4e4694d88e88768c7914be305a310478f9d1e7b58b9b115c74a27;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17340870d951dc61ee32fadf784db5cb0880522b00735db36afd9c47da85b904ce5d5f4d4c834f989937270b5071d8de5e89dfed9ac9d7a1fcb29d5b2d43f5e3cd988695e8fc1801e4a65bf83b2f90e74a5876adefee04d497a7aa098f04d5c28607750aa506719b5c1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h504c9844c23e7e948cc5c42bc2cc2d2e6da6bcca83e5a91bedaf4a616ea457171cbd6e067db29363304c5d7be640f3c7b0d0959b1589c18aa9b5ca2f8315a030d814191d33e70666234b6aaee643fce3f0afaf3eb22e7a071c71dc09e8b977e87e92a633ebbb44b982;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf97cdc300538b9c36cd89cdddcf24a81277e76c3ce2f71cab7597564baa81cc8a1b3c4b7602f7a7f936d38f5ecc73bb4231ae9373eb38e4cc3e5cd710ea00fcbe2cde19d4e3c02325dd98d98a469361c690fb4363baf466be353da48dcbc12fa7dd58a44a6cc7d1b06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h61fbf639e042626b4e69e513cdf32ad3e0b6f5fbae673f650dc8e43387cfdabf57477f9a6be3e1fe752d0f0a889cc9374cb7c04899b57019931bac253a683706c1071b1ccc75dab7e27db5a993fdfc02e42234dc8a7821b13aaac3613cb95da138790ed4fcbb47f244;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ad6508fded9abc4a1f106347869f81738fee8f31b967d413a4a7e7ae9d2c18d2cff6d9c679c791b7024786d802b0375e452c54fd7b3ed80857070d50227db3ab3e7c28c2401a322a2b4d267e53ebd3ef5ad071e546a37a6589b830128b3511febda63e37e5afe3720;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59cf257e0c2593cd95fee67bf117e6ccc11ff71f6256c881362730ce3df66e16c0aef28a6723d5f435986d1da58e2958b039a50f4166a79733e45711b0431cb8f47d7df9fff9a3aa7b97b2fe3cf2a623e21aba3b512d55b1b522904d9564aa8a50b6b31d22c74e68ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ecabc870b18908e81bf3981f6be539a39e9f404ffe99f93a782aa3768b77df096eaf8a364cec7e7b5e79453c99db82e8055f2ac6ea62373b0a4bc56290c51b089a326287311757f1ea0a267fd3ed34ddc52782526098e5a0522330b5943e447c4d3660b08790697d58;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd4ab99b50abec1c6ac3a0b995a3e938dbbf345864d762fdc0364bdd7c2a727d09a3f42203e22a95976af2f6aa3bb6f0ad1ae6d0522616b937fdb56b259653b3ad7041de0d5dc11d2429e6865179f87b702682b3ba4c7323a6a28572a27609cf4b910168ddb8072df0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ca044c46581a529d6722086a5582a841ac34c517b3b0f7a775ee7daa92d21117d79234da4d858d1069c863f7e0f5cdee6db4082afd6bf158f300aaa9ffafd3d556fae7de2f765ac60c1ae85d8da6b669f28e45e479017bef6eee5d63b1252dde4d4d6736ee5f59bb8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3a53526c59287aae66ed5cd38be74ec289fb618121d0bec3d51912023042ab8145a5e9ee85d8f2a83c84a2ff5c2b882dbe0bc76572c24a2f7b730ed4c3a281e94aab52e28a1a429aa663eff6b703ee13862beb1402ec8082523250a21fc7a71e9c38c8a36ac8f6045;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4167abf66cf21e142b57246ba48a19e98cf444715a2607a25145fefb9d3abaf4fae975f6907ea641e49f8f0f9dd37b251178bbfb8f63dce5c9af3da3f0d29883fb411a0ad7ffb0a9f698c1f61349d234ace3129fbbbabbf0cc7bb5ec42dd731532d8a630e3dbff9ed0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1587bf5b03316316d43b987e75b936f67de1b631cda9b82ba4023721dbf39f0295abf4a1b8a000fbc2c752731a91800a78f3353f5dbadd0400c3a684a04136e649364ea279a2f95498f2f5cf7d96577c48bdd583e047ff600dd0061a72c3b2737915b58630c12e15f96;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17208e91171d4667eeb640bff5e97881f56a0a6e8c98a281c23136d924c19bee678daaabc0dc29d857cc24d6ff6f0d84d34db9a2fd69ce4f7208f69feb2c4550813eae216c9c7c442472e2e0e3451ec791e3c333db994ae753cbdb7a2959a8e277f1e48482a72b336d8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2eaf2ff5a9207608291d0bdd5d2a844319fed271fce1eee011416398efc3f992a2806619a93c7b8a145d1975dad74b167fdfc96787ba17a8ae768b753e21b7a1c483146029ea9832040368a654e028c02aec233b220ebf1229e5a10c97559de40aab1e7c03b0bbb0d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haab55fa844ec1680b710dc1f088dfaa68fdcf013aff87ecea759b4bd7319c8d71e5f8f1ef3a2726ca3b7ddad363af9924ade5c67ec9e09e78e1850bcbfa6fbae2d831cc07cff427baf0970941b281aed8b5cbbdcc3d7f3abf1553d45dc2cdad5572b06ba0fc3c89922;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd837d0a19864a600724afd644880a349b2e5175d4f6fc8fe55fba8c535378c11c858d796bf93f19edabafd94c395da299e4fe55b4efff5f730c6efa4c7972269ee075db65d2b16e6794be9f0a983f1bc4102cb67acf995c1816113d0834c6b91e7d8e37a50dcd8ab13;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1458fea0cef3468b4c99c8c3971ea3cb0c4522637781224bb3584fa1af0d726d89a8982bde79ce55ad9a56ef7ccaa07cc6e306d9c5268b49351524c13ffee820634e7b9657ee0357258a886b696acb64b0a224906aaff194e4ce911cd812f147a2a1609ad19faf467;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1728ca73fcb4b71bb7a3cb41e704ee1f35bb1b9fb6d557999f4e2df9ca31b1546bb2beea5e833ddbdee1b68f92942e40c39749a7942f54f661870c803c7d5f6e26a097172f5d8f8786779596ee76419b962b8f5abf00916c6a23f4f0d0b966cbdaa38c510f93720886b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha9c90308767bb6bbe1e96bf302e5add457c547d56c11da261daa874c110978d9679e79064089069b4399b4f0ad15a19c1808060c991d61ffcff0fd721e811f1b97b7025d041e360f49acc95ce75853825022330c2e8536849e5871ce9fd0cc24a9990b816d0a9d599d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9b2a6acbbd3ab4af0559ac70ba13a9bcdbbdf5d3b7c42e03bdc84d2bb01b368fc71a8ec47063ea7d23cdc1ea6945870b47f91bceffefadc1e0f57d3f57f338ecf57c5e8ecff73df17cd26d1db4e53e6a257a5b071f980b27d20971a5edeb036ab6e74b23527e19915;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b8e782c79d0410a3425ac569b5c0b9bb8c268d6e6841c56fa9d3a7827cf295684f9c3f9d5a35b11d814e8f6384d1c7cbd7a53cde81ccac7c92a7a10eff26b5cb9b28d99b8c181e64da3d6ce742f54962b709b9908770cc2a6c4dfb3eb5633f0c3e0b3777364d65c439;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28a52e118a7e080cc4401add558e8ae9c6e0539ec684e810337cc398d0f216fcde561f817186437cd07b9764267b685d611959cbbdda55e2eb4427c7cd8c9f90506bcd24da4dc2b925a1c58e677f4339096457b2c9e65322c44e636bdc9850e03d9f99072c30ea92b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5dbdabf878222126d578d68b9e05123ebbd1fa9c08dc92b2d14b928eb4e2ff58c2f24fc08659337c02a3059c49bc3963cff08cd1ce03449ba9caa9fff96472be0ccf8018a716708c926edefbef3ca57ebec9bcbb08f430d46448ff6f3036dedf0d188c1e0ca7f77733;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d0ef83a9db9d5e75d4d740e965dcd1812d1806af1b846ab2154201a52c2292fb828e34010615a2b48361024a91800170f55a20d08438bef4d1c8b87f5913b0984127267f97f9af8626f565aa1859886157333801c97f3b4b3bc1fc57e723eb8e6c06e4e2a32e0161b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af43ee6adae90338266f736b30e6442daa620b5d6deeb4bb25d1d2999eeb5ae456141627ba83ef7468076c26b675830b6369a1ce8d5d1d8756ccb510346dfac6697906c674dc1329d3b7e6cf53f8c190f86a1eb0dd25370cdbe43ca2fcb8ea09231758d749d6578f62;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h191efb9c905e6d91b29aee7463ff89d6a6faedf54d77ae7f65e27022a1ac5214d95dce3c8d7b4ba8954ec80b5a96759a7d174db87405e058cad4d791342744fd9fd889e1dce265e2924d4845c2efa58edb5ec7e3119c3252cd8ce92b5e8c7d7fd1fcefabd8ab55e92cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b327f1517b3c7eb65ade8e9fa4208f5c856d9cc42c77420e55e1fec806e6e7daf80f37c62a71a1667c610920a03ad616c4ab9b0ebd75e9d2f131d2c9662d7e5799354ebd821c1ecd15126523e42377b8c9c9aee16772742451f197cc903f2351f7f227e030640f66c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h51d172d525761a54a9accfa0f4ed014a95bcd13b261a17192212adefec74e0c12a73a0cf4bb1b16a3fce26eb8728311d9c8c94ad36be4b7ebf66b7359c3393e7c6380b41b04f957fe7ac9ffe1577bb67285f5040081477d2ac137609230e019e3e7293ec4f154a76bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ef875f9240f24187a4a260be25979db126e9cdf293820b84d95158ee3b6adb0e856cf65df48aae8c309dd247ef6f068eb6b60338dd85e75b6dd75a6341e0d02232baa16aee40a66661b2bcd980d62abf83530d3020394c5ce8d55f3def5de0c9436379e44b5b952d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18160ff132ee235690a008e58cfa9c27e30096503f191d4ff63d7880090807846ced029e240868a0d97204f00ffd2a753e3c3bda990c3d4ec813a8ccda41d9710cd1d27078b529f2447d32a2dd9619937520be1eb9e4de411c8ac173a41d13f1f6edf74e4bc54e23981;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h764d39013ba40e5b0bbd0d353e6637df86c7c3315a8bc8cb2a8972263801bd928b4e6eb8a424522b1900aaf63d79f09055a2b75fb9d9ffad6e2db647d43c5c73830e2934882126e9c87cc051f0a454fbaf291255cea9c8cbe241e98d9402e9ce7cb89a15f29be924c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c727dfe788200d629cd874010291af4d46e68c6b158bf1acc05902dbffcbf943bbcc2fbdfa35374a8e5b0df87a16039acb8624a60e4e38a334589447a04eaba70d4f7593f5c437b1106623d4a0625312f2afca8a8c7f88b5547f629eb25d38c14d61bc37a1a49deb03;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c5cf3e4a123e45eb036b4ec61630d40679137bc79952eb25bed3127ddf1b2929b5153d0cbf758fc63fa00d297ae3223a2299b635d53eafc0abdc34d7d5983266693f342ba1473334e32a88ff5698c6043826c6aee299de33e5f33ade9ec8b4a9fbfcb6a9a466d0169;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ddae8a111e8177ff5ff79462925e103c74ac181df956a88dda9c515f5dae38c2f42fb00ede9f29d7fa582a8fd4aa8299b41582993adeffb377e03eb9741b93171198cee225ac40f29cd78a861c45a18d0d6450d1d2009906974996e190943ecad3691a2357c63233e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1791f8adc43512985812de51c2d75f8f24e036bf5e96287883aed275fa5c7a63a430c84d1e27e4b6d2a6c3809776fe61d577e5a08e3f4ded5507a67456f0d9c4f6d6072f47d29032b6826cf6175cf140c247a76c357812e26957ce2e8d6e32f123e5a809c47b77fb7f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0f89151f7b395d08a1a1e123b1a6f17d681bf7162312a4da24654bf0df67509ab01de3622b4b90f1c55ec284abdbc4f22a0e0d6a698dad57f01af86475cafe0d36bacd7220f32db1ccffd4323277bcde4b9e712010617d968a299bce393250cf32ba650ef2f5997da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b8b220bfd1d7d1f9fac459ffc4efeb8d428955a6e380368d311dd0d305fcc0ac09b898771937872596af373065ddbeacf0efb8a2cd643ec4907769259564968a11dc0ad3825016d24fcc24a187cf4759b25f05538f0c7dced4b5fb780185e685bc3f199abf5e15dd5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he863419f3473985b12e3f97d69e3c81549a3ae3daccdd2e80680bf29839a3b1e12106133f77d55cf563cc16f56a621d4dd08afa9dbd24ea859f648bf75b83845aed35ab967e37eeca6e7f5c74e915a4130d98e4b8e7ba07b0aca2d30ae3d9f138644127428a744ba20;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd6cef863bf9e2d5b651a19f75b8746c72c72aec74988aa65ef4275c7c944c77fd3a257056abc02ec450e2975de1825799feae08c4bafed24916884f290ea2144e9116fca3edb84a7daa409dec3d09b0793a9fdad36f3437887fb1a29602ef1ce124739a0746b5f3e2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d5f6cc8aef39fe5e8dad7e216de3dd806a255d6b9e8f7c135f865f02b73e872e15c6bc9a4388ba5096dc974c478e86a727202a39180da842ab306628d8de9dfef785696026f821291bcac62b6f93bf57d511178dacbc06b402d3472c663913096bd60f7e4f025c89fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11402d494726fd419f2149cb0b7697fc67b238ad037c413e531fab1d978bf40bd30620f7637cb8a624725e8f8f8a6ee4d56f7ef2d2a4472b94800f1cab821bfe0f766506aa3b1ba4fcd59613a65237670dd3141cfbf6056a1ce5d100015119b54fc75db6dff0e6ed456;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ee89ab90e44a805da3c17daab204f0f683dfd4c6ba0565437cd60d4ab633e768687cf266e39eb9ea4067bd82948d8126489ffa34be948cb7dad8ddb286957c9da05537d66a7675c45ad93b5a2891071e26a0f909bad75a0f57220642eddc9ef2dc5806b93488d772d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a1d9a01b8530d6d33ea88423f4306161d81c9c206b0e9a30b7a818f52473a91f33c6593b4c14119ec74bfbd94d1afde37d4e8d3f39f05d58171c52912fd3bf6c2f19b4fadddb3ea7b7a11e43599df225f9984a636e8b9c5b944782f0c2aeff30a14de3ab71a222975d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbe57c2fefd8788a10f0238e64eee34fd0eea233ce8af18282967525e8a0297a80f2f0e8680645e4e333c88313df3eaaf0c3a5de4d1f64fef767eb29eeba184aacbb2675aa2ea196ac2264ad75b82cbe131c715adea20bd5590402253ee90acd7336864a412f550a641;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ed9b83ddf5835aca10019677088021ec663f2954c557a0439ea7536a08f1a285c4887a1b21f05a70eeecdc6e1b63bcd92a482f44dee8b929dc189ce55fe300d6f7dcfdb1ec2e3a0462cf275804f8a2c60ac3af1acddbcbe29362563a78d9b8018c7cd83b4ace240ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h20c2457f5841c7d6ea37962c5eb440486b83a7d80602495368997e2a469a26899318222e1ba54951acc2421245831a51df57da60288a1f46ebf55afbefe76bc2880046d450dc38d354a5e59a0886f08764a1402546461a5c36915c46a052dcc2ff853f796d8bcd530b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147ccf4928925d7b92e30de70f8f7ad8d95d4685a6621cdc7067ddf584d5b8000e8e06d8562652a0e8fd67cc1d85a48fed85d5669b71d5ae48d3b7b9f536718a74fd75afc68f67be1ee817a8a78c5ddf4b12ed0733afcd6052b381e3ed58bffb3ee0e580349c4ee1d3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he386d390ba04fab7cda5c232275e037f10ddcf10b117a1ef6022e96424855929e32d6e833dca112658d69e05edf2c5d7bb23587f16b0e6edc6dedacfcef4a6c141f39d8863f6fd562d4261d1070b4a11bf7f336e72d832cba56624b0b5f62a183278a3cbac2fbe366f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64b920f798a21adda7f714f09eb792a12d6578114d6c874c59951745303171b5d4c1316a203588de784f94eac33905017371758a2719a37af31291bc45c638e0c39751f656d06213541da209a3a6abeea184a28629a68627299a0f3b296bfc64abcc0227b09d64e455;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102699e03390b84cfc25305a8412474c7770ab0cd5f864fc7b1418825dbc4852e66b95c9640292f868ff5a90dff9836a970e05ae08224b4a816d9d7fc85c26c8f25ed8c196af2f7e9f8926ebc316b443a2d37fedc13237bcad9978ca62a0f665ae6b80d1515ee02b9ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2342e5a05d1ea07780c2558c8298e9140893a3d5a77b92e0a4593b0986c4c626725ddcc1df36313c8c63fb38690766cd7ecad9b439d92cd969ce29876b990c9adb47d29741086add8b97960f2e5b9524ae5bad755899b27d78d867dac91e06a1059e178a95e5186e79;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19bf54c9d1bf1eb93a1a3b44af1252eed2a01242771c9e09f9d9e87d659b8e96985ccb344da3d6ae8aeccd265820d1ae2ed54ef9d1f0eb7dbe8d546e3bfbf2b2db00c89bb91d9da414403c163fb2df606b376f553b0dc84a17c5a1db9568c8f5bd384a2f6f25051017b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h112f7ecce6e9a17ba854f9784a0d042a7edc324de6eaa9a0cbb2a5346f1bcc123e85f7bc7a0e083bf8f7ba2d81b1e30d4c238bf896b155f34cd93f2b671876b9d69f18e328ccaa93a3bc5fbd967bb5dad7d63858d75286204581b3ff781ee616b5428813d4ff063fb5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca3946070652fb253210a983e89d5fe5d6da75b8087154791e5da69a684b8736ac3a4f8bf73b845da693dcf8a98e38b946ecd5a1b4ec9371b5b3912c4b4a8be2e99948d1be0462d4bc8a10c993318367049b48c931f373a1ef40338b0930deb9fe545671724d7825cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbaee236dae8871dc21681d30ec0bdcfa9ef7a97b6b80030238592dd54b940a7bc0d175c8c89e861af17643931797a61444e6e5bfdc1847a7d990fd48f02c661b3596935033d61172b1eb71ec9e8b7b8c025808b5628883c1d65f7d6858c4af67795286e6cb4d6ca893;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ef83630c72cf8b3ef636ee438503a1eaec901f872ca49282e4cb833b17a39f1ca93fa3416f91b8b41a3a0e71e016dd601c0217075ddb3c87d29915ab70fcb191e3af3d1d078c1c4a3454d9498ea98e891f54b9750bf82bf89cb5069a0cde18944dabe7d2a40591678;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ecd2cc499adce789308fc2cc176177d008bbc8663c877223764f6d839b8403e73762a60df052aef0774e8e6828d025402b8940890952c3beefb4857735395c9be524dac1081b772eca83518239c0ae1cd002ee0b4175bceab20bebdf88e228c97544aac1fa618a0462;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7d9e7c4d4932bd2cfed5bbc8a2ad2b264d6f84dc48e9883a7fd95e1fe5831d5ba77e3a89529633e400b6f391347468ef83871539d381ea185e3ee9b0fff1812c719e0d3e3273f9f217044c964e4e14f4c826bb57263197d69a0c09a361e6d03d47eaaaf53f5210db5a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c6ac206d0a099f8fab9ce8ae46f4266d693ee96054de866bef1a545c88cc6f63b5d632f10a18a8a6145cb11757c0961875c7291e88b4e362116abd431e8056d09c7af19d146d1f887f4e037a538a9ab9577a6732d0de22aef1b0d2758618fc8a4ebc7c6d993661683;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bc3d1ac0ee4fbb0b90032031cec21b900ae6bc6807ac1ed661c9c02e40a2524469e141db29d5589621ae8ccd4705e840fd65faa99aa5c272c5b3c860129c8e29b00d1d39e33c9dd18ea4164e91e96ca012eaf11d918ef4f40083b185d688bca7a3f9c41c413488b54f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19688f9dbc3fb92bb26d590a0cba9c73511a9670ae11433d164435ebdf1cf79ecb740cf89e71e1dc9203b544c048ebe88bfcf4ad5210fafc22367acc393734d89d8ecb1cb71bd4df1a259b59465e1b3b37e7c804511818564eafee2c69b066354aabc123d0214c50187;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e94c1437fb49c0513cfbe6c30bc5282bc9cc5eab0ece79a8a1d634e30aae1a5586180d4c144bd04852df5fe54f1538ee2c4f5d1bba000347f9862b359ea8cc6f32b36ef1c5dfa79e33b58af50ae0ef4f8547c49537f8c4bb828d10bbff883f4f7bd5900d7f4393687;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174c5346d7b2ab94d2d7227569b49c9a8e6573e13405781b6a26a8221f0d16ebb359d81c5d01d008b0f79140caf27079b787214d195dcee0fd59e90493328ec98a83ec2b58a63b84413571115112ef2bb78afaefb634185b777c6645fea7a43f6e649692e1137ac4001;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6777ce5778a5da30bb63d853985550cb7d7b551868163116e07cfae53f5cd813518825816d98fb70ef3336e84886f5dd4497eda7cbfb965f7032f33b362ff0cffc664184cad7108008173e75434ddda5b7ffe6a96f0639820a110cad8542cdd2d13e93ea0af5572162;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1055f91b4f6e90448cf02d2aee76995d522edc04d0f67f9d0fa2018a140333bb6fc4e90867d4afa346b448c2a7f00a59773debdcbe14ba65173ffc4cce81f87a57158a6f68f62a1a1eec47e08367db057c93164af770609c6e4c3cb29d50b9b20a2c8dd2a18339b3b88;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1531019c21a912ed4360d35a9f0fa5ee24bdad25ceda4b7779de66f40447c651826fa8715951b57582fb9e921ef5311c2264a3659fa0ced7ffb5881a81d3e16501624b0419d72c24c488883038feab80b6e8db50ca44febbdf5a0482ecb964f4e872bf5329d0a0cfd55;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d854e1ca40c61a227a2cb09dc015d593dad1bf59f883b745a88be51e7a36abc154fb089cf6873a8a17346691b42800ac01c371492142c2c2a2ed8311d29c69db146e2a055ac3f7a87aee9133620644aa35d16cd785eaceae896345a61717b48d474b5e3d6fafca2f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170534b0559d071ade3a1b0a3ef1dd4b1ba366615502551da00d9d55e083be66f0988c9ec27fd7437a131da60b8ef000626d961fa765f4960a0048c021c3e26a808159e4dc04b210ddb8792778b2641fd0a4b00214295643b4320d820eb17d272b9475321b0dc5e869f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147a7c8d8196312c9dac4c74e7b24488f1ce0b68f322816994824ec8009ea956d86852f739545319886458b9e3390b4a6c2132f9a26fb1447d54251914c74ce779005b70c8a3a6486c6c297ae4abdbe547b35e27b7feae6f9cb498959a8db2a7d53c302ccfd9b4842ad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aed48cf7884d11020fac8c23eeccf5f66d0072b34418bdb5dd690d7f69b90d2442fb9be811c89a4ae1591b168d86cba453358651a71442c15628152f3971193542ee2c59ed251fc116f3d9f265a72b0ef53f8c388859c9215bbe4e6ea6b2323f56e45142466b1b0bf6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192e215842e728540199de030b3b2e820e7016d52dfdc463da0e20d879a6c7e1b04c2d257c1050456839735385ede0beb2004ca57518456bce3df95c8c86d5183f1646ad3ba89e8f79dee3239ae98d6ed0d36da3662a8c2866afac578acb5e6437ca44e19e74440bdac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a4a9efd0574764b5da62b90117c4d2c84c535187188e9e185ec9d65b1627894d395d5216ff70ae17ce4de9e85221db4d70089fd0ad458fa84af8a1a3ccf2f4273446c820412827d7866be956eb04afda190257125583bb9a89bac270d14c3c5682491fe35b1f3f42de;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f90179dab530fda97d9189ccfebd1453543522b6dadc2cb54f7d2bccaff2766446150440b91de03af6624a5b3fa911067c16dda28d6bd81beeaa9cff3ac181aeb5712932dcfb6aa9bf804e49af1daa0c0d265ca396aea139db5b804d9b4788a50e251f1442ebcff25;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1283873735c888ece25b8afae1f007bdc1a28030d346aa30a8f84757c1a80c604d5cee268f9bccff4e68260252b1fb340f23e6accf8e0773419725197a52cb307d7ef142a40b3682a3adec0ba5134c2eaf4c38cfc275c473de6218c960adc0e8e173965322de0d8664c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha71bde729564e581d475009e46d8cf1df5b84c89b47a302efde819bc594e5f45557eeea1ff8d73f54c790bd8f59f3d8489655ad53eb79be01b6cf7c34bfb87c80c4b876150b53ade43724c9c8239e20bbd6038a45adc58177bcc6b6bd6a3f01c7fd57096c38a20e5bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8cf3db2377f46568c231bcd8a51f067906d826ed0f6b672f7ce03d77cf35599e081bfbb1ae08c8ae5e10041c2de4139f78b5dcd3bcedc65cf86a25df06a8a9a1fba7097a20dc7598f05b5a16151d710d20e529e6731a4cf7a08fb07e2f6a675dc661cc66be87681db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1204c84d3dd1962c81b0b2bcc299e1cae0e7a488c61ef65903c9e232b172522bba2041dda8c0bc8db9ebab202188b3d573e8990f284ceadfdb57d0cfd6b3421ef5429073032747f290aa3fd55b13af38f9e0d52bfb3ab6fddc06be537fea039a5e5b34bb6f5521520;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17c84d31a73a4d0769725739139731f9847039ba521888bf8ed8cdd8b11f39378d2a0b2a900582e40a0c65c0770ba6d73baf58cd8d0e5c09044f5689f4a1901d96728328c2c372562100bfcd8dd43826b1e79cbee64dbb724750d204f0b239b9afc8572fd56d5c146cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1546bcb40f1d001f370abcb9c6425097d3a0248ad9ec64ea94d73ed8d9cfef792c12fb773e797621e64db49c83422a3d1a18ed8633a0ffc52ef2f33aedb6e4d159edc4a5814968ce8c28f71a7688f7d4cacceb27ed07248ced087a73326513d0ee120e411f75d7c0e96;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he5f33d292929f35077c23efb8d7c3862fab27f0a18e1634f39ef7ed67ead037832463c89adcc0610789cea3db975cbd5ba303625427fb89c70572d5e65e6b65a1a5b41ca0d8bfa36a3a0e36552bf0e49f440a22706ede7ab7cc9df1feefacad8614de1946590d2da64;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hebf4b2ce2136265131ba484b4d25fcb97ee4a5200b0177b6426945e886d67fde16c04dd2cd50dae08e878a176603046f990d19e1f27766871458757f60b224259247ea46a1b1e2383386f9ff05f5e1f9f9bd343369d80e79b29e90815ad1e77ee6db245074cdf502e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a3f2fa853b7125bb3a74eba47e7eb0791001b15a67c1a7ef2556041a97bb79fc86544c24ab99da4b65bb46374b9961bbcd43ca1161d6a512e35af3759a6573b0e74913b4927306abc3270f860c209ca3e6dd813bba4859a77d798209de9ab1706a0a2de1ae9435b7c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcd4db9a86e47c65d787aefa333bd1da3f19d32607a24b833914aa1250d6ef5d43febae1c6cc31ec0ed15797a3aab42bf34cf911d25b1e70fbfcb889f8f873766ae95a99b3c83545f93d3bcf29d7ea03c3ba6fc105dfbc4848e79206ff12b4d98bdd69503f72ac94597;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6234722af1cfe48d785d817ff8930882c386ae4a05e1d4f2b03d1f52bcfa29c785b075f9c296b94a37416c8321f6d4bded34fe5f00eb7c8053d675c1b744f4ed8ec41b09d1b0a8d09677575045b6509e636b554b422a9594162b75d7d1bc77c7623c68e35e7ee4d495;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c13c29a6aa308f1086874a354c2120623c3fc8a7b7aea168f2e0ed87ca34e41d2e833a2e1caa1189309a8dd7255aeb1ee9111a77300a25e882e90600ef756e6849b87d08eab2c5bd6413f6d71efc4b5d14add79ea7f19c083fc083b8af802a9eab5c904a3d225e28c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he4c72c3c1849872960b642027be99601d20f8147e1c9b6b351d38c2af31b9a9210387e53acc105e0c82dfc67431fb071e8f08a0f68e11841e7fc3875656aa92fc66b4ac8b2284fc6f81e08ca3a408f7ffc836f0b66774c34ad6f6506bfd0750b7c3d3e3315e193df4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h858673019050eba09f1bdbe864b9d980b1dee9bc192e219b4814e6fb1588135f038ecf6c9b257b37d9de9d987d5ae5b716ace0b1a63afab508d4d4c569f2db28468d39e8cd8923fdc9099c8cc67a272561a5ec8834d7400307a3388e9de897b1c0072d9b3a2a04c14e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbfd8e005c6ad273980498e2b7eac677957d8efd0bf008c872e98c86a742cd7fb0fadbac4d821b9324320afcd27fe9800dfd12f23519ea886f019bbdc5dd4ce3db583424ad6125316c7d6089a332c3457bb30fabce68764021cd6ac14f886821708df7f7727b7be2a3d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7074cd76d02e66de2d6df6e741c7b44a31082cb5741d1339eec0bab21878f8ffe556ff5a4aecd73898b863ac019dfa39571660cfb13d62dd6adaa92a4d904b6e0904edf18242690bca4f3b8b701ea4ed85826ba6c6ccbde8a2a4db7e908454b441fe82bfeae02a292;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf370bc823decf48b3ee224895b5dafaec819931beded3059757ea5be913658a70af5ca190364084c81e1ed849721ba3a7b5683ba5cf2ca4a1335ccef7d56a376bd98d964c1d39ad625c63b3e054ac157f34597c650c932d81fd8afed0443f270b71f1851eb91868ab3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9e8ff84dbcbb0cb52c20474d092b956dc307bd0ca9517bef2eacef71c5a1e7ac723837e20145ae1e1644a71ed355388523a3334a08ab91342613c649457f552ac751d10b856556f8cb97a89bef5ccf79fc0024ee7711d5cf526b0b14f6113455407dca1e5ba4fe7103;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148d1882abd4933cf0c7ae05f8097f35f4118b8864abc2411653ec93175386c05f10f27380629f093e59b8777b7a418115a6b7c3e44f648337b1648d47f9a7a43518d71b29c6feda6fe6a105461ef54f443ac8547622f1832d3a2a6cf1326288b48a3cad2d277aafe58;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc54e8e132f1ff0ee2f1cc7010db12b23e4d0f15029510ae42a10e6e6decd1d6b3942bd8ba51505865e329989be45ec07fef2a56681ad133c2c005061f7af686587eeac2de83d1e7460f62b81c4e0f429ff62af968f35c2493ed4c022bd4d8ba83515a3115399c3961;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc4f296fea339743ae128f75e9c452279d239a8d7f7c726bf607530335ef52963958815fd6a1a33f53d87550e08924fc8c061fedf829db6dc2d61485d2ae79af278720d920b0afa12bb5f9feaecc39ad5ec64cfe16a394efbe4dc43ac820c7ed218c9e5acce325a55fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f46bd630ec12e604fd5d3c376ec32d5c65a2b1472c87343496e6c14e68c82f53daae5b4aa74e566d28f7c7442becaffcf1695bed3739a07929b2185c3b27752e093e7d9f29b8778b77e1ddcc6d396bccbe60154aef036895c668273c89398821e350b41e70d7353d03;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h151fd1c8d5d6772e2bfa04eafbebc6e58d0237eaf3a4d4018dfd0ee525b4c7044931a5271dfc0c9645807e4ae121d6f5d60ccda58811a81e0fee4c034fd6c0beaf82ddd66a4c06fb70a0fb14aa7e3a1fb7e1ea30fc44b12a2666344cb6cd1233f3a08188126c6e2d897;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5ce782651da775cbaddde4362d3ea987f6f5d969bf2b41764492b92d7aebf514d7407cd3ebf8b06087c52f7caece3970167f13a01169a19351c1f4d299868426eac1aa335c2fddee6a8e811306c278d56f1c98b5feddee9af761e5e02acbd0615e138ce5e2d52211c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17f4ef2b4a60fcd5193ef27c7ece350dc6c6661ddfa67a586744292af439989cfb4a2f0cf7a739cbefaf651ade7aae2501df72d1bde7792d6d49db0064f4a2cd9648d07ff25b1d4745da5808be9bc35a4a31b9c5915acc37e814d4d0fe1e4687b7a45f13f1ac04aa9ce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65d319a1d63f132f0bfe86336eefceb8c901dc29c829e39f48644bf0c7bd33eb2ac490d1c61257c0fdb7dea5d8dff84c534ab69d2bfdebc745b0a0b8b17f672abd967c85c96a5233968fbff7d14f1125e67cc23c8229790134b2fc9dc0126530ff84e9bac3172a177f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e5605b09f929e63c309b116c8106111edef20b3298a05c8449aaf84016fb08c4c5e4ac4d43f2d57c89e53777da73bfa34924103a7fd9f61ba22d8284666d4973040664caa46e1f4751a5bedceee63d113735791ca43fd2083a1e1e8dff61e85975e2d8fdfe1f49573;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe1ba5009b6bafbfc4eb766eaea33ae2de8ade080f640990d66a77a280fc1d5c14fc0f41d4958829a66b96404172caaf7b135f14fce430e4f2c3c7df0c22b6dae3b1fbde99709c0381318592527268df956dc5f660089894b47d98407649a35dd05b5d1bc9331adcb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce2dd6a692e0236e3f3c09e568dffbd8d885fe11a73ffefce4a3888c327f4fa968d034b8a78ead0405b3859b7f01f46865cdc443bea7b6c5f454483d7aed4ecdd93952a6c3ff3e2df7b63cfe78477335c1a6fa7d4df9aed64de33fab93ac149c85db0f5403277b77d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d0490dc0e3deb8a9e60e45cdcf4d951e29f725167b0080d88298c394e7551fef5656cd191abddf199caf636d06e953df88f1617b592423f4219fecf3b1aad0d07c7298d7451939177851a677daecff92256eddead922850bf116926e8ddc3a09c0cc1afca40d8fece4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha826c240d059b6ca6b6490d07e14bb85b5fb23b091890c1ce28eeb59dd6cc8c345e798493540a6ebe48364204347ffb2ac23b3d41fb9880b4447845b85f81239335c859f36526980d1e0f4a6b1a83b327a7d21484e30a05c9341ec7346f34fc29e556052ea35958016;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h49b90bec3adbf809663d96ae68152e42ade168839d19af0e0120bd3843fb41e262bf0fe4ca565eea42ee34f323c1f29e3798c7f6a804ba2cb93b82a4b56a9448e10a5e4ef674b7984f292f708f9bcbbb806569172c147e3e2a18c5ccc6760f3c45bd105ee273329970;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4aa9003202d883baa36e1f237333acfd51a2828cb24f55f865617a6f4b09623611e554e2ffa2ca8119dd8a594fa453fbc19e51010befd5f693f132a6f06cd22b11cdac5fd0ee89f6e3f3ccbf84ca6bac82467c789c2080978a3a368539c8b4ac4826cf5e379a6b2d14;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4cd96f7f5bb202e2ea4640820894157f029ff1ef13b8793e04dfd9aae12002f2bd2ed351a5e93ed157865637c7b66b9206884fe6ccc5f3e46590e2170c67628dfc0200b530ca3764942e719384b84e546de40c371e9d3d9f2b81a4e37a2c03e2c4d6dbd0462f6eff3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b6b4dfde336a6ae27780a18d58e80361231b4dfc3f3f384d6a38f34c68aa0be765815e9b7da6bf91a4986beb3d1b0dbb520ff83aa48f64da8074e67f53edc832dc2089a8baf913779892898e7213d23848eb33a5a915d2ebc51123bb5dec66b4371799d4f25a47d53a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11d3a0e042bac5ce766a29eeaa91f17eacf77b78efd23b0c09f987b513ad08e8941563e976911d660f210129d81f7f5054a36f1935974349dc6189dd90835d0ca034ce785981146597625d4a17ff0d0a071e6c8c8c65004a42433fcea21f5036201cbc4c251ef844a4c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c2edc5190e12914d856b4b9cdb252c662660f9abc7ab36eab4e5240889921d860a7c33106121aa0e5e33d4377e869ae89165c962ca01e1d3e47eb49c3125a14f47f29f3a6233bac3a435088b63ce5b9b424e05c9e47b40ca02f8ef857c66122b8b61c6030f3de3b107;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h966815e135a9983cd63daefe7ae91e66c0d5721e4d498408a4bc1b299e25fcd488354a0d9654fee829158c71e774569e8c957bb1a68683f15b095df998ebea51699260bb495c4c237a6b723e53bd18e3b11fdcca08f32696471c017630dbfea46f5af49772a233fd37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h184de048f320ef2b0f304da9bc12fe9ac24b366f095d59d8bcd9ada434129d8ef82ddfd547e4e10c8700599fb17da2e897a078b6ea0b9d37a58b705b25688592d9d853e64089cfa801b2dca8150dbcf9a253e34cb1d0cdae7d28bda2aeb8b4913bff854b1450c6e70c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f10090908d521a72afa44d878a26621ff3102d70135b02b14f813a7553cb07a06188e67d51ace2ae7d83571e6a53362e3cc487ed957d2d94033617833b32e6cd6f9eba17ac5d02c57f045d7b06883db86b62c76188664df301cda0747139785d3161bd47216a516e4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f90b650a7b4b64aff86fd901e8a6b43e63625c203625a155e5f0e949a2bf4d2612a70cc40e058290bb7ca7c41c0f518d4bb31c4bdfb6346869ba1ae1a454234bff4c22a15b2b748177a6f9f5090d2745f266d250e70f3a9663b263126014769e138f1afa6007db148;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116e9aa240f0d6526bd863eddeb06fedde4cbbca7ba5b1c9169d28bf98bfe6418bf2b0756ec82c7cec6375cba060c0f4495b805b116d31cc6c71d4c9b571ea9083835ce56df45157163c73ea0b8855dff8c6bf0fe7ce3031ccaa9c0d3e720a359ed8e936137784634fc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f988b11db7ae61149fc5d3c8c1f0a557506dd6ed5e842d00651ebc7fbed766d864e4b23475f9742c9004f249f03d3cd8821c033cde003087e080b019383c5a0893feeffa5b7d59c5e6bdded42749daa02e4dfa85f8cdd2a5f78f5e83ab4925b4ded43337c607a0c598;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cbbdbff4e6532c8283459687b77f12a097c587d73ddcb0872a819a2b21e66d8f3af467817a2d6eebb14177ce1ce7ae1a4917b666ef7e34cb608a51d440ff7743e036ebb7b4dbc658305c427e28f46ec6272be30b459113dff609eccac9be394e62a79fc8facd77d0cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h676ec79cbc0185d13079906624861ea35d7716a16fccca74a127bac01e6c7abe2284c7e6e175d0e9e806d619bf07a75bb8b56710009233f0191f0025975aae83a25a56d99ed1bc95914cb001cd37a5f9b40e48b42d5e09e3ce6ca349993e9a6cd613c2b399106066b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad1110d6361861c46cc25c3da69784687c46a56bcc332c5fb22669121145b13eb2a511d7e5907ed289873d41943ab9511b2aed44a8d87301fc58c2790ec5c05428b0c04c80793ca5e0735e6edc23d506ec7e6c7323983e963803a0f42cb2bef8607240dc07be30fb4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc958b7e91185b7d8a9c20d44f68645f07bb7b80c63a3a10e813c2e81e30482667e082d0e960d76f26829412e2eee14d24d1cab8797e7fff91c94cb6ffd4ba96e0c5bfdcdf9983d0440bcdd814dc24f4ca25ee20b7a1eca113c2f56af1998cd7892c1687b0745beea8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cffaa69c5b2794527f643b186239775000608046087452c20ab0ad60a43e696702069bfbb07dfb5e97839b231cd94d94d7e7ed8145e8d8c3b7d07bff38779ddef15940d9d513bb274fca3c692dd14771b0bcd6bc61e4c12fd7c1dafc76994044b5ef50730ab7e7e0de;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h546e70050f370ae73c455043fbe9f974ffa1bf3e6fc610c9b6aca0fc040fd8101df39f4c411ec51cc95f18a2aec1a07b19f20604e094ebbae0bb22a2c1febd7d83b86631109bb782b6843100a7333223dcfd99102b48ed8c734ccc2fd20f704a1348dfcb0388330b0e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c3c96f21a678c2b3cfbae66a56bda453a8f16b7623b81ec9b8aac1aedbbeb5f6ae879715d3bedfc3b22ad1cf7e3c071725638eb670707f6e6582cf3947917bf52ae30d3404273834dc2b861c17947edabd52922bc9d7c6fc5adcd91db5f5d7297b909e26ff26768b8e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9221500810eb2eb189384128cfb9e09c5d6dbb1f553681076a82718e262df385b234945926b37b0fa72984f27b5bab3f8bb48a05115e406f1949ffe7bd0ffc7bf2f69d5bc2fc4c085565b2d7ded169cd98923022ec09124bc01e4363eacd16ea25c2994685ee9e6dfb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3baabb733526efe3c8abf01d530071bf6c475e714ef5121b72aadcc88b56a53b878460339244a6646cb0035956b128faedf6fe1736e328f2ce52975c595aaa391cf5a8d88044765ea2a7010ef50d8018974960c56a7875edf558eeaaea02d91d7556c2dc732c6a515d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h93e327f3e1a967b73fa67de5e996872e5298fc6dcc2d8933bc4ed95910814e05479e324ab19738ced2770a173373f27692bb0bd01332281b3921e392ead2d443c2d8c764a303a0eb6de52a6e70b80e64028afca63a71e5b43c1bbafaac51127d4916f772a4111e9aef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he6c25135dbf50af7462dc2aeb2ce85cf9f2f013a014fdf0afaa5eefb725df8c73284ee38909e9fc5818ddf6247a5c06d80a56d4bd51e0c7176f746e4d29fc5c08c52e2648b6b3168da0ddc5e1bdacf170b28cbf2dc8acdd20ee3aabe7a0941524608dcc3c4bfe06ccf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22726528494cfdbab03f9cb51ea93890f690e5d048727139a67f8d68e7dc65cbe0ab9b4a6ddcff45f3516c6bbd61c9a7dc355cef99f142917f4a24130ffbc920d7b7753d2a7b82255dc3c4c539f1bd7681fd1b7ac2c7b94f30aec4106c7f83d37892d399ec867e53bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26da5de368ad69634c4179839f7ae6049e2182b212886092e522a5c17532d00545d54b2ef788089154da42c85517331a7ed5a4267b2d94cf99555297a496da79e7bb652cd6bcccc7381c6c28f2f1c3e73e06f467c8cb0959960fabc6b35d7f5dad8ff3c1a5d94d6d29;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8467a56e154fe1ea0df85f71a5b07bb1f5eb6b654cc4e2e6cbee5a5609fb5464ce0ca81c54571fb642b891bee38ec53931498595488f4de0a11722a490d6ca70fea8426380f80fa060b5e842b8e7dc51f154aa5f8de49f5157ed8fad14bdb098fb35ee30f2dc1f09;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbea2e8f86d01cfb7c05842af7cbbb582d69f64b21eb81d4a4903bc19b70e30913c9cc920e9a8a499110062dbd2863757205f9230164b0fe1111c49f9afb121690b251b1e7c8d219fc81ef3e86c887c2d3ff0e2804a99adee43410105317c497f36bc01d91282055c01;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125ab33c8b96f258a3fd157604fdda29fe20ba870bcef91257cdd7eb02f503d33c519953a999d01f46e8236e9124a831170ef9011a3c0636d18a3a11abb1eb2e7ed4fedf2e3965595ce7279ca6402294773096bab7b708d32fe1d8f9f7750cc6fc7300a03846ea0e5e6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179102ca88ac442021856807b71efef9be7bba2664e1cd92447a7ba5f2a1d72b2cf482bae6093c311419ec4fc12f3c3aa990c2189d39b386dd7be20f1e6caf455c8c2cce7d1c69f5a30724ec09cf509abefb5e34c8824cc72c715e9925bdcaaae1aa298a31deea942ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1feb2e160ec11656719a60296e8d268038f652b6b8f9fd006558f591455324dce8642e866304ab398295e924429feb9c6f30c40c3837f9135b28d95272470ec66d0cd79cb501807e9000bd0712002d6581f38969a72d4b0d14b3368491e092f724ec6a762bce37a76b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h115deb8604049a5f4d4e61b90a2172a0fc0b546062b21996be40ea1b8250256d3b2eaef2b578c969e69229f4d348a378d9d8fa806475e6e2e261cbf576315493cffb49d4c6c0a0a0e0cd3818d7b3664169fec9740bf0a3a4f39980f325d9765135aaf87cc4daa3fc9ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h290b018af7ccb4c6f7b12c78fb4404afff14e5ff8cac43531af743655812c7d85118281c0a4752d70bd5c906e5a4f4f6b9f8518b8cfb702b4d873d110e46bcee2f71c7a8de7ba7828d529de95766e5261e1a6a9a50d5b1b311dfc6b154c5a8c56671d54d61add40cb5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hda2a8267728513a7efed38096e3a9b792742642e76c17965fff1010c09fb7207142bb550314ec95ef5444054853c91df1cb712887428b7c7ed5726e1455a7ac04c6fc6369c1c17478bdcfd875b5a9382d9fa18b9ddf564fc14d4cc95d828b5490d4ca67434ff3e5ed6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1abd6a24be13c98fd7c20bc31ebb249d3e0ea6ea4596af4cfb200b8aa67d11135f7bdb46e79e3cd56d775841601301661a71f69ec73be7c937747d9406ce2f7690d079fe6632251e9fd7f83cbbb4e6d8aecf11b103dfd8493806aeeefdcc207775a77a171a96b7557b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167d3d7d2e22923a3957e3c02f3139520cad0d7a5005da605f1200a4cbce7f6e1263d98f8b412fea3dabd222ac046a10acbc3c83ceaa3f8739149360fe404b36ad39fd7b142cd2181a164959caf3f261af8d1e2d606eea5429ac4b30cc27c54aaf5f78c11dd9b67d211;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e0b50b87bd3b06d80a4d9089c54d20b91163360be684cbf4eb8221eba58cc49a1dc71db421936847d0b549b058df649d7eba19219452a7977087dd60d61751327379356d839192ea2f78de811bfc5a87ee4d25914017170d85d7b2981cb5aadd5de916311052be89f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6394ab6edbf4dbf9f27026cfe039d635e08063251a88eb74a9619a34876c4b6e8482a78c34fe4ac046595ed0cde303547b6f5c5bd161bd3a60079c66d538b341ec895a7f5cfc18454c84a09e87b699ad43c30b53169cde86f9b7661cf80aa9c05c36afb350eb34fbef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c440df0be379b1af3be797baadb4e4edec192bb41771960037cac1f10d45d7d1db924b0fc30e8f93b988fc2cf61ed9be40773087496d7f8371aea66956b1421455b396ce5772665f84fcae21ee95f418bba2af24101056332b006eb5e6da6e50708753e28e3b546662;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ebe89ee4f5825263f1ec0d2102496eceebcff79d66261f4eb67f776528c542b0efa562f2c03ebe8e95d42fb4036911a2248e2efa1c5d38e613a9e4182b8473a16cc0659f65eccd19470e9bb322991a3029bff60961de7456d373f52b8c20a4d6ee82c70ebde1385c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb77da0e74959a956f800f60023ad8a6765b9c3e0d4531f07be6e5e5e47001fb69e231b09b4293e76d9fe8c52a8d3e8250c72098e42464abf11f420342c459b7e01351a5a7897a745228cbe0ac5764243ffbabecf10961775dca680f39ec63e3a9f25301457260c1ad0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c8dc3ca350218beebe986e27d3bcbaa558f58d575a24e914f5b0b2e842a31538863b9f9573d956c8bc5e5f5495f2fb46fcfb8458a25828df2c431db683a7c1bc6341c58c4d97635474d1202b8457c0795bda919c3fffe816700268390be377d703d452dd77164eb43;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he20fb9b6659ec464a234b23fd7c5c641e7ba02de0cb12c3593eef6624a2a56edb5fe71d84d76d0a66d66e6520a2295d21099883b90f439b78cfc4505f8f28cda032927f2437ecabadd8b3b1dff7ee82de9daa0b351cda3b703cb04725ede9728c4fe1308eddc0cc352;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d79f51d33d11cb11baf921a62ec850fb4cf08ad1e067ad367d9de878625aeab28668f3f07711caf322ee0bbc7cff9e312014adb40fef06bbe3b6719ac5631f2d166e96d7c73344228dc09b25a69f3b1d202c133259c0be127bf73e3d8bc9ef7636d0672c25bccd6c8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2dfeede969b17228b611417e09b12d2cb0b82da40433618b18b19fcb4aa7a559ec945eea787121a99f9fcbbd2c4fbcd2064111a86dcf9a77385e7bcb33b5fa502726e90e48d9ed81ed55d1017d70ead331656bbebec40ee2f8797b2c03dd3a829117d2ffa5414fb909;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcdf159939f41b1c8474ee7b0acfa039da26446cf31bab205d2e0adbb9cae2deb8135f440d06915e9d9fe16d6ed3736ff32a3ba68be3703caa66a1dd521a577f0c45259e645b31e5cfd7658c316496857b6f61320b8c251280204883149b2c5a362eceb301d0e547cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131af05860a052bbeee107e28ac4974a1b3b70233419be26dfff300885d5ee70dc3a72cbb89eaa45a56f2233e1b7c1eb4ee6f8dcddb8e8d6a0a90040f1c0b46503f67c22a80236e3b5332b62a0fa5a7302ec5542eca9851b09102f6c386a593642249b123aa7d900817;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fdbe8555182898150b08a11becbf9d0de8cda5fe825976548f1f544e326a0cf34b7abc4cb1222cdfc5630d57bc35070cdc5aaa75d07fecec34a7c2cd7b4bfdf18636f7fcb0a4ddae19184e2348ad6b43816306c7a8a9adabc0860b6df46a8e338ddd5a331d608f44f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h816a544911a2ab306c43c0a79ff91a78f678b9cd1ad8364eb4dedc8f8b908b4411593da875072d25caac104ec1c7d2f4c355622d239721d5754d7199a7db6780aa3d14fefecdbb2b373dc006dce2c8c6ec0a5f7adbfc444f2cb1dfc341ed956cb85b8379558166b82d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58fae1ab970688e5640477d6a6d066803342fc7da196187147eed2f2047d9670ccb736367af89539187d2eb58648dae6629bd0b88b9eb94101bb3d02bbbcde8c556092c68923c5f69cab614a8111e9686a75eb1c577d49bced94ebf1ec744bfbf1fda2d402319fc1c8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2ac1b72f91ca0890819206443ac68f0501657821baac65018fa215c5e65e1a5100581ef3638cf18ea94c22e354181f4e5b6e81f95e13c2b3e0c8e8d2319bb4c1b4a4e284a0367695ac447ae4ed0ca471220a5d0512a50d645425c08a65ca249711f267990ec09a2cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h606e349528fa600d7346cd27d9d76a3efc1b26c7c0c2b89e28b9796cf17b37723ae03f215a95bcc449ce553e2614301094f84bcda58642618dbedc6630802ad4a8692c0bce2992c40c4293fb31391ec5a92b42d8bd13ff3a7ce018b91726130324468d9e3dcd169c0a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e3113b979cf97598ffb529699848cbdd9ec62c0a527238a67380b28dfc11c703217d88a1160fb024db8d5d0b33e98f0e3a8d6674a5dd0f3f14a7d9864cb5366201d4ed88ad27a3cdca782580a0656fd01fa53f7aa239b37185fa6c847dd336d25430b71fb0759b545;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf82bfb1f0fd0640ba1a2d4c313b2f586f315ece5e027972752f2f2f8dce3b02a8ba6c481aa0bd60fc2e3c764e51930befbca19fd80888d83e52e3ef5e4b6d26fede77205e4f39ce71389af628d7df94516a0b89976efcd6117ad0fc23916b77509c6617cfc68377e99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f9a627e5a5d5b2ba3465fa43e44a9638d0b621047d2d236a6dda7e276867ba3ff899b6a170834b7ee9b95d806bcde8486571672e7380c0eb65f77f43332c8db87194233c8ac46f432c58b75cd9a903c8bb463458a43bef0103909773157c7901c85df18f5fe66223e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf64d58cf01ed0fcf6e5965a914107791b7a8e63a3bbefddf0b7ccbc0e939aeade037b4bca250ecda7ec389c756a5b9a04235156dbe3d7d16fb453ade0d322af8f00418ab21f1889fab0d7c7fe87fd6eb0335a8af6b691f971e9a2f72e0665c3edee1d5aa39a51a6f34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67446356332dcba8cca3bef9a1f0a13359b1f61cc4b043a7d42648c9e4f6cc0e6bf7a1156f3d676a4040a0896bc0226553b0f5c2f5bda98e3fce298c8ef3a29d88a7891616ea9ad7733273b6f6a6859abde7837c14a581731e8f2fd8d04ef431d25b4f019acc6333bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba7fd4ed4e618b768a4345e639d12999ba8f6dd9c46a56b5a134f50f7d2cfa6fe04af58142bf48f1f91564614e0b1cac898b3c6adc32c89f122176d6da57506d991fcc63bf955f9409760a360dcecf4179f2a3d83011a9dcaa57dc7407fcaee83514fc51be32906fd0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9afa0f8fabd3fd73aa0ab0d8504dd26190d245bcaa29f7ae5832b88a2cf4a45439f165a3ff8579913124440ef261e258d6f0d2c91758953f50459c9c31c5596be2522c60cba369407ab98b1d7df6a09932885c038929312c40346cca7b54ba0ed233d8d355bc69708c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fc4e52349b3eb166b87588cf38c91db7634bd26e05086f9732bd7957d994bba4d3750e3f30bfc4d066c889cfea4d0a52ce2ffa77e24e5fd8a682269375d11743f6577a1bf5a638cff2358d628f324c1a9eefa152a93104da74063b33cbc109ab11b46150cf5bb2917a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ae05352d6b57a58681d3a36a92da7e0fad6ba1c41f9169c3d7e7f9923da56577f4fa2d0a9da7a21045584fd76b0c9ed7342d455e243aedc1050117e5c2094b1c52120204515a1020f1645f1aafc9f4a7efa59fb3ec29ca00ff855f50f861c5a317c26bd3fb566eb17;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74c16562582b55bede2d1c54e95e29933bf8fe0d09c6951cc68cff67d080fba8a6e54bc6b26df77bdf057eaa20668242a80daebfb48ce5a04681951ccc1372afb1895079753a7f4c95f9ba25c4b7b913b85ead4282af0527d299262297b45aee06c101ad797f2de596;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1506d32c4e948ef037658f49c82bda8e54e852da0ec19b11f7269f1bb68ae8fb690dd9001e2158e2606c8a3629835d6a17a50a5cc7f308d2baf161904276ff227b1f93074bb826ad4a4080e92a88b0021abbceb5cf9cf708655f7a9a8c7527196a459a042a30ae0f3e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb8dcb62e3e497aff49db643aceaa4dcd74b8d9a54c7f59f62cbd3fa3d5d3322c2016ecc12804fdaacb1d432e1bae667cbe2aeb381568e8808199e1d806d28625f128df3c1954a8c5892eb9617feb242d71389d839ffa80e6a677636199e18c0cdbdda9b4d192132045;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1df78b72729c0ec90c67d5852c6b53185037fc445675c35b4c0301bfb9354e35820fd16aa3db4f73f04a661aab147c5637cffc6909e5d8d4af8d650c6d16e64a926e39aa68600698e11e7df70139dfb947de458f96251023112fa7147b92948ecae3d2f797d8ad08943;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5fc79c1140614506dbb1c972c583e6c90a17c115b02b4740f5fd4b8176617080dd80ef5dfe56c51847b5fb8dd0df3c038aed25ef3849e0e9fcb452ab9a694de5b9be9a76ff99541498b749b83c309e5558bbfa40adb820ef946e2b9059d60f6bd0dc81eb51323ed2bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h118b5aaf2ce8bcb25bc753341f51a49efb61952ba198a1a61eb0cd85e11282492586822c5b3cdbd6c1d8c63867f76b534992151c786ea5d54ccb0827f3572f8992a021198da9c17bedf19ee4cac92b52f04efd93201c6efe2786cc8c5d584f27e6126a42a9efaa3d0a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h738325efa430c4ff2e0be51afe5a1a28a4deede2dc619bf10e56e1d0023c9d04b5165847fa9cb29ac7682b740bd07684f93a5316516556ea8d992dfb17474cd417c62ea65e671599fc9aa68dfc8bda270754d6a29ba36fdf1b93f27c24be309e8f54b4c1ea56a2c95e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc05c5f6e398fac150ac3ad54dfb9d32ed8e9445830d1539d043ea31b0017c5a9583bc37c68eb2773551a0603a4bf127d13d1e3db62820954744c1c265b69da68bb213bf66b74ec8e4cad36fa8472a5f753f2d69583f8a19c9341e1e545f4d88c2f3f5575bc3dba7836;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b9de07bd0d8727c7d23f47b42c46ba55a7924fdbc2b2423c6ad104b3d6b3abbac36e6d9c1efc17189e331bb520340dedec3e220b247bf1ec3d0d26858879aafd5fccd488e7107b9dfa5ce69913046928b151757063f634bbda76705c029f5efd0d82c1fa32a7ffb8fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1116cbee87fe1f37731cfa3832c8492b0ccc0117929ca4f0f8e114d2df2109fde9c0e21854d56a2a7f1b887e6478e0645738fa7e6b44a86f3094ed032415afecf5fbea4ad31bfda5af19f79814c0c921ef707cda6031c0d4a64780ea38db8baf50a8e6fad4afd55f7bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha7fa689acf8b03b2a0e40bd4c97b6976b2269399a49411ee57d45115a3f7c0918a7641c746c024db6c98a2c14d31d3b8d4ba5f7d313f922925098b32e430f9406befd880fa8df562f7e4b58bf6ceb6b545dc49b95c33f606804b795a79e93ca3fd40a74f51948b2e32;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b19828967fe580cf39b3ea5aefb3316417695d389ac0667ed3c3bcd7a7c25fb9022b104fb2a419d709374f2bb70f643c7181bf184fa2b3205a71518bc58975f42a1db555d49f4715e18a8079466ab820739feded5bddaf406d98b04d6b0eee09f8422616c21a229bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3fe20384ee5a8647c502087dcc799d6e03a819318a0deb62f385ac7453fe9ee23ccbf193638134e825f3dd8c01ed2273776b57ec07e2c67da70eef75c806aca269afdca9c0752a42107dc90cfc08ff001f7cebe0f0f1eb62fe524e259fd38caaf14b995e7c30e859f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0ad39e52ed17d0d21008c2535a3d3a69296708b1f8bfaba52f6848876358864d09d249588ef60d183732d76b4521bb0acf3c74d20f8dff32da2bd7371fc3965a8898488d0c83a8f4eed96dba2001dc024a1e3b40db3354b3c7eb01089618bf52a61588c2b3262169d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e86414f95fefcadd2d48f8c29fd84ae85ae1eb7514dc6b6f73ba9d076cbd588301d2c819ab713a54bbde24ceb9cb3f5bbdeef5bcb08342774e5dcd2ab827cf01e2e5953cd14e646da25c1febbfca9fa59af451f06419378b3c1931000b4f45d58200085f922090b649;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1707b46dba037e6da04f3d0624096b28b91aaf4c6c8a8b64cef75a3f51f2aa3812299e5a71d2ecd900aec041c7aaffde9bf6d72cf8241542263425173616ec4eaac04b58100327f7e0397a5181dc7a481ef51f3ade4f987ca276a8805574baed9623a8e4ce74b3d03a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha866010878f6ad787e0355c438272d4dfd7df399308badc616b6cebef7dc1318c0e500393d99f38a7e8fbd33bc9f1e2c6cc673992898af6a593802aec7ae8aa3e9b5c312678a3738ae24f24e915df680b4722989eacb60e82ff42475d57f25b729bea6dbe48b0af4ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b762bb624fa4a7d4ae4d0bcd27a582fea36eb05d9a20ec11abbf2c1490ae1b0dca2b1b3ea905396e0f78cc607b7b4ea1a897ac0496d69d80a7df02d3170261b617ea36d45d1c20acae59d9e6e2c65bf0add22f30c223e50af441abeceab111bde7eccca44b248fb4a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h856222072c49f91e21924fd356a15037cbe1f103d027e9c378e7ee8df0f08f0d3ba7f002eaa41ce4600d01ae3aa2fc687d4a11a9258ef943808ec3ebcaa71b868a8fb05ae63ca50becfbc0ea659e1bbecb6964e4f91e8f32633b8e2ba51951d3891346808fb8a4c97;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15e3f586e68121e00786a47392e39887cb8f7ba598944ac99734058ae9bf53a867f651f838d0c0b7e2801fd556d920bd42866ae783843d873b037fc153cd02272e2a51dad84307f50a8f3be0a35cefbf3608a99bcfdfefd782de025137682e4e125bf5d31b98dbf3cc0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bdf2d9b1647cb45780827c8cb8f3c119e4a0ce082f09975e181fc87244d80536995374b44a69f233b15062ccfc2886be68bbe9987841de465daf29b1d2c4a58048e20b4fd51dd0154a4e8c357f4c63f1ac485989eb13720bdf3612e6e50fad612c2a385b75602f2324;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1211ffd30d43ac4f8b562982d1d2cfa614f9818972828e3b65f738d2eab9b2ace52fdd633ce2aeb3a6f37e1a84e92f17c269946be3cea993a41bb19f72fa907d5c24c6eb9229ac256880e9da9da4cf1b415fee796003fb9ee1419b1413e9a1e3c5229d7f48d67b78edf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae803a5de67ebe2cf42fe422f7141ba8e962cbced1e87bc1825c48595ae086e13ec8bd8ae8f0bf04a40c49d49eccd8c3b2175882fb82c989fcbf19ce899d7e4d81603d8add64a34c8927b91760e4a57addd6a8e4a11c09a4365527598027508128d167f9458e445e2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbcf9a9580f2d0ec467cc1ace7e12cc6e6762baf002b0d22795a6b4023227b2008de7a1af44ad1ce3372da89842d410ac24dc7afcab9884b032e3ca0730f91a990b25385d172f66b6842cfdd67016b3f3ed625c49ffba9ec1e2e7ef85c53b3d04d5c5d9e94849faf8c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161bdd2b6a5344c61178d97d6068f30243e7306491d3b2d28ed8de04c516a2327e8a38f4f2058bd15a8af09dc07e626a13fdc5a68d8c21734512d3e35726bac1bea5f8dfc682889357976e8072461b4d7e46171d0b3c4f702f3ee7299c4437520322bbe4cd6c6dd4be1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h66778c89514b1d431898859ba60241f43e635d13fead973641f8a10a411aba49d9b8e8b415c24100e69be7ee2739b8f389f60effaf347a63c667a7668ec70e4b92b4f80c011a23a7ba617bc926e307f0376a7138b67a1af7763ef79fcc6ec6152eead669edeca13231;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96372938d00ea03438e1100115e84f9239d234130876374d8ec71a443e84a75946bb8bb6ccd16a8d43c537cb64f6c896ea989b6868e9c40a7fb896b3da19c64cdcf183acece2befe94f88aa3fdfb599aad1ce52c119a2f796ad22fb45192ef4d27b88f55164655e3a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdd171feff5b92312c9f6987ec46f4ec85147dcd3d4b195b3a55635331a6a89318a0e060a38cdd06f2a979b8748c59049e666e66aa49bac14d2848968df15fdd4d2b12d6c076e755fcac65c35c37256dfe5aa4f7df301b70ce2d7d08b4ae87ff86f9bb633d972ca2f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152434cdc7bc6ed716e69f1686b849446401852c39a8a037bc4b526fbb726c7e80f2c101a18f64706a7b22d7d4a840f68bd5427866dff4ebe28237be3e82a58fd53fa72781ac4bf16a9850128c5a5d9816b4635b8d15df781ff7d0c3f3738b65e106d770ee2ef440285;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h44f5a0b12ab9ef736bbe0f71320767b1eeff50efceb01397edac93419f696b8b26a982a5acdb358a19c8f0650ca483974a5cb2a70958ab956469884630d63b375c573387380c20e1f8c37b862de83b1fdeafed5b1b07c87d79e908f8065d807ec492ee9a45b8b846ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14c25ed4a10eb0834cb5a1dcc2569101436ad588ecfd46b0758bebbeba9845a5f564ed63b4e8bf9eeb8b76c1221f2780969f25971520170eeccc5dc4e0644546f57d11f4598a7eb73b3b010c4015a5e9a89a95f012b4fc6b042e0f5a84d54d6454dd3e6bb20491b3d64;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12ff5396816e4f741dc709fbea1c02d3b0979bb89a45a6b6c194d67a6e22bfa17971772469e68606acb5852e5c5620074493e2b15cbc892b51a09c079e64654d9d5269e2ec8cf8777f3054753257ee894786c31fc323af57973598b53be71284ca9947d6960b3f580a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1606e9c524aebebaff3f4686e108d8d979cfaea6dfcb745a6e5d373ed72e2efeaf86d5d0e583ff285af7c06d1c033b0fa25aa1aff1506bbec51ad002f059653100ff37495fc8030fda1d21b308ef9fd667cb0a0012c725c125f527c971c5ebcf05f44b3ef22a6562566;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100b1521a99efc84f03be5840540fca5d9c5bd3d938e53c6704dc58c061bce8d005c33924838cafebac7a7e4de98dde4dde6d644da7c7146da0ceb8fff605b7e0f12fad8750d70a1692b1b119e1b3c3b56afe39103ba48f73eec242bef52e8304e375edb3f9835a1c82;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he1833935d403cbbd2de606c07d142af8dee081292b48c5ba5ce6d28a7a5f59b44a5daaaae3aae1a6cb3608c98d5652887e050ed6c66572d8c475d07c87cf227524d5232c6ffe45536df2002f764d38f820cd45d4469bbcbdbcc56351dcade204881a2acfdbc094f966;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1968f78ca3d1a8978b9bd51b91b6c4a47e34a2df0cf55e55a4317400a9020d59e19a9713b2fc756fb9a7c41d0d387ac133d0349038007c2d99e794b76f43fcf5fef235d4dfa748e8b8b9bb8e8f3fc240125c14ef10b98aaca36da6280b63433f63285a26f137c96cbcb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15eee961d26a64ae004b2b9930d011769080583be1d54046815fb17cb49ccbd31a952439bf4a9213f0c95433a88e987a99832389a1ea5746c4a16d4d4be9438c9a058da615df27d90769ff90a90ef2f2263d9d3c24c42209551315b9cb030ac96d567a980cf60b17fd1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h30ee76e198b151e91307ec7e7ec85643e0a3bc361493052f72e75063cedbf480cf2c01e3b13ce4328422e45b09a8a44abdfdd770eec65d0a5044b16feb02c9adc986acf3547d31c177c8e50b78079a1b817e026ac86f3f0eff281d28cf441a82391c54a194f865fd5a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf00dbb4a4287e9a069e684cdf3c8c2414fca405003c7c4de4ff523c561642f872268ae80e2266608a805e35a2c788f8778cb54be53c6aff76aa37287c283c7b186f992a13f239984104b67d434fdc2bedb0a64a25e3a4dfb902027b89fa469d06777e66cd158bce36;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h33778c9be2a062c309ac2a1cbf374f98223670da99b7faaa87fb365336568613ddbfe671a4e2653aecb3d778fab5908a70090acc29636ebf1cda15f74431084b9fc87c6be3fcb18be34b97f5fe313a38617d6843706d86dfbc05d08dcaedf12de6863ca39eb04b4bc8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e2262f5bebb1e80afc9cacd301e29838de49998df80dfd1d749b8267958109615b507ae7f5e87136f1c5eaf49b33369aa3a397f09d30b9874ee7f7597da0e9740f895f7e087fe689f5a375551bf65f9e90576dcac5aa11420062b7129783f77caf15f2cca146da27a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bec6a9528437ee622c5da9b47af846bb638e1d43fe6e6613ccf74f03b7468f8d6bac28b76320a50e3f36fc6b35108af8a889df837e57c90517dbb155002f2a38a8e342f21e8515c005b94e0531a57db36b1a37154c674cc2778d916b28d851c98ce77efd7a350084c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2685504d0cb3d150309b6d1c543e133fd12959a5ab2a536c85bfda25735ffabe6d6f9e793c73aecda7857ecd95dcf78a0484573e563932bb1f37a400fc7914a8feef159316f05a0e8818cf751ace98feb21bdaf86e931f66a4502e65e50254ecbbce40582653b3e05e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h224c5ade1340effc84821e7ddfad86a8be57ab635de265f0aea8e1a806bc0ff7988128f565b4fb24a19ce6c542a8dc2148800b84d6b0c62957821693fc1f2ddd4b270d742eb35875018be634a63b92dae8e65ee8276f625d5039c5c04fd6f604d8b9d61557614cf834;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de50630f405b811f344c5519b8f590743f16ed1278f4e3bd25fa4e611bb5076efaf93ca80967a82ee49e57cd41dec5c5794df7e3cc9e66aeccc95cbc144b061f1aeaf69074b95e0937fec0a03316bc017a4f376170e8c99079e05e65e08ac87abb8c3c61479041c3f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62e1e73c3feea9d565db44fe1e0c2b7c6feaa860e441db8b3f69fce25c5d6e5a579c2a257f0830e206c2c64eca9d3e3a074602eab78333a996f8dd17f607e0f6cc147d589827c29fe5d6860dc79624d917b27d50a109697242f105733200ac0d7d3c3a864c0287aa2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d4fedf0f12cd3bc80e0b549e041bf5a700527a261a0a24c1a51229f75a63c616c8e45a0cc05fe1207d9f1d8a5efa4c282f7df402b4de40664a74a818fc58a64fcce5b820e161e750c6bf1f5b5957dd2aad314605ce640b4241c89e2395fe11de65979dd70d89eef1f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h187acddaf8e3b9bce32790e378079a4708e0e3f11e0f193af21b6326eebc24270a662aaabad773ebbc165635eeabd49bd2c12845a7fb88ffb49254c2d445d2179a33cb2c2469fa1a25296a2896cd9bb3f5257492b6da383f040cb6928b707d2bc06f29a7a8ff295f5ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa980244d374e377265d4bac4e9aa5b841790003409173439c04008c869ae45ee991c2ccb5cf80b3a0ce39fab1426fb928e451075ef6ed1dadc7f06d6918b5207c6a0f93af030d3a09e2cf47d021430d71e296ab5096de3403358f4c8c4609d8170f0bdef5ace80417;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e377f652fd8e86eab17ea5b73db977b9b7c7a2709bf76f1fa8bbbcd2db3077185ddb09587c800eb393312921d124d363a1affb59493639c53bc7a08a15c0e7e3cd362066789bdd7825bff4972d751397583de1f6b64c65d526de90f835b290f20261414eefff9c99f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a3d13b79e4247992eb4cf54276b28844af4a32e7489e0b6fae55d872cdc0c87349b4d3cf334321df9c8df8b7c8659f59967f00078db6386381ba6bd7fcab0542ab02d42bc3fc3caa57a0f944cd95532fa8b9d07040c45cb29bc08825f7046d3977d209eba798746a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3f11a83b7ac95766ff490737583ea79e4caf77125170f54ba8ef1866422a55c41e5a06ee4a2928243369a737f089da8f8233108b97c3e875b93b52217fdd2cee5cc96df320666f99c35efa81bf711d5fcfdcbc7316484e748fc0668473a007c0dca586d03522580b18;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a512690873013bedb2e0e2818b3ad29c0802d9ff235f69e9a2691297dc6d356a9c3da14b3e783b51fa32e11fe1ac489ef7ab818289e4e72b51988a3061867586f8fb81aa02adce39d9d301d4a3a9111107c5aa3e91d21dcca5cf7b6bf1d021f630a783dc9c8c6e18f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h186c2639a57a5d257bbe06400bcc353f3462e31aeb00d681c0c57444e3095f1d4ee772236f3c7e90efc2a0ac1f90eeaf16c38ad4da867c2f786ad6724588e1f990a83e3a84d3624a3d950aeb17fb7fa6bb2657f7a68d5db6ccb595879bc6139d8fd90b13f20385c4980;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d420ca49cdc4518e1dfce62c2eac9dd88677bfc7be78a6f27932810aaaefa037a68a63d0e708d5ef9146c068c37ed196c9a171ec56b7953ad55cae0077d54850084ff397fa2a9b7c7e392ac7050a9421bbedadf8a4a6b8f5e31a61d07e375eb0e9e3fd7361e164e507;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc476c6c1e470e6b866646498087105218caba29cd38f0b8df2b7d39e21bc91a5b90a2a0f25af6b0c9d961f5d1622ed8f58b95cd11ff95e515a788d5ed655e78fdcc89ef5f79cc9152c66dd253dbe3bdf80ac3418b6aa60339e921f28c1ab91e1f09efc98add53db2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a65f9ac2ed518b9de01a7854bde7871dcfbdea07b20a959712102fc24adb123d9f5762315129d9a66543f67e93d2ef5ecfa72fa47126a3313e7f4d1d40dd9967d758e9d1347513ca398a63cbf08babec2966a3c4e66fe1e06b71ea862246b1098f3ee60beb637172fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a1ae06ce028edbecc46d7640a9576e9bcfd4ca29d0a87a23c2f5ec0a5bb46dba5e289f7b16e8ee08d75b9cb7685f40e55d7fede46e5685077566f0ad3ca768e173c1499f3522a4c85e4c80e13197f66aef61b7b488972c57810fba7bc1623c90a6233387ac97ea5f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8fae76b756cbfc4675a4a01f9fab41805f6ba502c215ba2d479940b30369ff9c8593d97d56b08627319db4da012d0153b25d4f05a76b3f80d70b2b3be644684f3502993aaad26e960ecac436fe48e07b030a93311622c7da4a274b378c0fba56435647c0f4d1c09e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1061d1475466296986950fc077b464beed565e26ca51ee14ce694293e7782969c44babac025266a01b2ceb660c34e6fd75993029c34f0fbe8b0b8f7ef6d056aca92fa0f51e48ed5b66c9f9695993d19b3d1af8cb52d89291c14811838c9e944dc7d129dbb831e732049;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2566f0c534f05a5bad15c0026685349a6d286055fa7602351b5fd6aa8b68b66a80225e17c7c84330595db46e1d5884b7116cc4980ffcb58ebdd52e09ee2bbcf4aa43aba9c69f7f09d595fe066979ce9992f3f7fd5ad5def0b84bbfb1722620aab7680af7b320b232a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb17b043b3856ff7c5685bd54b8e00fff25aa3acdc7a719e71dc70c3b741ad773408b0ddde2d433c9e9af9c8ca45e34cd6a2aeeb04a82b72670f945692ce62dc272c63837630fdec0353b3cca08427044950df4846b430d797a424543445cfd85d35eaa090243b810;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf209a8471a0daca0a7b9defa63da82a7a98509039b856eccbe0c839de8d845dfa5f03b7ca81b329fdf186e4cdd32914a7909f691086b2647c43fb2a41826d8ff70d83a2f54c8fa638af2a3ee2e31da11ba89ece0b80069cb01ccefaa7d1c605da2ef61b4e0d76f0ed7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d6dc520108ef827ae83d0df43725f3ffc5291570c57827e392fe4028f91436a387cd2ff76069e2772c9a21987b0479e3e994c81f68404d5f3fe45c0f3bdb7e39b54d0388d05231e8037b73022eea08bb23e5829f0f773969dac8c0c19f73c99969f1745f5da5fc7b5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf902825e2bc14bfe212ece86258fe8b2185c098eb18fa475e2ac94554606e0b96a1a15079e5424a9241aa04fe1ddab76feefae783ee123b36de818f7a08dec8cc7379847d8a918491294d648ce6efcdf0c58b15e7f723a027ec83be1f34b88d0be588764289b36acfd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff5310c497a459133913ea138d33cf6739e040cc3c9c93be1784f81ea09f78543053d235f5df9e2ad988bdd7c134878ea4240c86e1910275ab2bc6d42d02cb1ccfba022e246f1af3c4ceebc4580e62e4953fab5ba1f37b834a5706c4a8a3982c856dc8224521c9aa97;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1465972058ccae79ed064a112d0b217420ba6bc5b4594d6eaa1bf865d37673ac5be8cd24f223fe9df1615db39e71e8628bd348d5c2b698d27e00a67a1fbbbda84688e37c222d621263ba86fc151d13a98c8e209bb644cf41fe25533a12466bcd785f84dda3f8689fa12;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1364856b528ce2911663a3965e2c7be94a66e2fa2cd6664a869526c720ee900d98c814b8935afe8417788556855de9a7a272f8a9d32ff0454be5e292fb2df17e7c2c45a73cca3576c76a4ac216480d050a3e3588033f3a63d95184f81140b895814e834de9551ef2bc6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116327c23269a7963c710ec3a2fb5f26265e1bd15163761d0eeac0e4c5e1d47b76388c297d384d3bd2189fb0724897208d4a43b77cb84bfff902bc5a0d13f15068f4fbb3de8e5f769625b5f5947bd285347c3e0a1a331c274b6d1ea280ac88647660f998caca764cbab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb9eea4ffc1fa7f5445f35634e8e09398204173d06e4adface1d88aac227c7ca4f2533abcb78227b3b38c02f687aa3902150fb6f22643b9dee12b61220859dab46d81866c6cacf31027dc6e7bf06df6484cd4f59236f80150cfd632334cadab3d8f4fed6332a5510c2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h92ce9f265f861ffabd1997c8c48b13821b8cbef3e72c55ba4d3ea7c1e1392a42faf0252467026785bbdf3b40156a59a8123aaa9268d9a9720f9848e79fceaf6e6ce76734cf34507172d82857ccb9adef744344564496703edb128d8e4ed64ef1d581ecbe272c6fdd36;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4efffbbdaa19061234f7d29d329dc17eb7abe330acbd5d5e9e339423aafdeeef196c4ad2a8d44bc96353320105dda85fc8e3cd6c5047308ce3d05be1bdda23947d068bf080c48ece4a4a693762a4247c09924fc5990240d0568791b10875377d915de12a7ba464ad5e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18f3d9b60b17ba3f608566694c8c1e7dd4fe246d1af44dba11fa375ef379287cdb0293895d55aa0f1d9a3cf101338670181dd34b21fb8426104ae27b786e87cb1b191064441af73fec4aada66e0a680a8f54011d3af1a0d0fd6a0fd225b215df77231e5b96490a22316;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf21b875f1c79ceaeab14088dfc0e258921905587fcf882069803a221f35d72bd9d76b56482137609c870d4a4ed042ba7ea8f0965ccebf7568f85f7bd96331c959254844a771c1feb2b8a3bbabff476164a1316a931c762cb4c531cca30a2721a8eee3ad213248e4282;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8aa31b170451bf20c230ed229ab1e095bed35d46d2ceb4d9b8779db25b299f95841156b84c5a9204943ab96ae003da8b684ff530df6e0c0c5ad4ecf1e9cd3619bf68c839bc85b05528db2e4cf52d1837d31c6513505b61b344f5c422a4ae69623fc4e382b87096631;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11193e3b004b8677782f880ca734bdad67f57bb6b4b706721431457d4c912feaf227122fc15f6c660ed21cfcca4c0ec6d1a872ffee868afd3cc763933a3a1f895596e9cdff8a55b14102c9ee1a55421b0b84cf22ad5820fd455a9658fa488fbf73393f53ff396be7e34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ff09722df8cf48358c1d84aa8a9eb3316c7ecbb663626d07682eddd80602c88b32c7778a6b20e3a78e0efd5212dbf38b5491be2a4393fdd1207848ab63849ac7416243cfa783c3c56fa404912a5859f6388698bfb2caa3df2e640587e8d0646f842357b2ffa7d9210;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75bc65fdf813abadc414981d25227ff286c6f06c2d2c39b6bf46e5b24a220e05320c6797b3443a462a7d06fb7d8589fe48df717ffadec4405198202f2bcd4a836f2da71532aacd33e4c15f573d528fe00c4f968ff4299cfbd5e8b2c3de398c470ebaa39c388aeded62;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15327fe6599bb53f023957509fc22160964d21f50f0acda901e902246bb19262df3af3cdc7ebd2566625d485a3404cc311ef344cef87d9b78017d6a87f46b89b4a92d54936fa3326034c6284eb62d5d223913e941b33c60cdf421839a3745a6a4532949f95b2e8b896b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3f5a750304337ca6406b2a4808724d57e75f5c97369b647314b96222ee7bd8a12d087b3015c414afd7eb06d9b0880686dbb934641d5e2848e91c312e97de09c4b5927342d8f0abc96519f206c1cd3bec60284918140d8e6e396057cdf46cb37d1e3d72bf12d9b01461;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16259db960ef33ec083947a0a5466b2a3c0c387f67efeda92572c188ddf2d960bad6118dff8daa7679e85752815d4233d85a41f4860d0bd087f25827c4f1e4579a33423e71773f1aaa67406b4a8928822fba46b8b3000c933cf8a576ed2741cf87eef46bf401df97697;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d58fe7052f8b99fc07b5658e059a53f834a9fb43e13913b76e677b3302c1aa867653cc7a54d5cd2ea547c208c69e81d51af5c02865d50e225527277f078aa1f58a075aba093fb2d84a36121a60c4f63bfee8dd729eae9d4c844c65c07d826631f9bebbe0b1f97da104;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c8688d53898f79658ce6f361b160aba06493df434ad16c5ec5cd2c91257f9394a325021ce978ec20d25ca12aa79e894fa180d965b5e5fe6cb8cb955811fdc98662db82042e203d7c7bd20cecfb4a915b0166a63525310d33bb03b5dd5582546ad0662e182f60cf8cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fd68d56cdd5cf20aded5bcf9930d8861497892d511319e3e8b8054cf742b1fbd99941ac0bd206a0ed3d0dd65b2163ee7e7f001f968abff465e62888b15929aeeddaa149aca306aee9868aa4f5899e2cddccce8d78c33736cd4e64a83e1eadead5628b79d42f7cd16f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10589273f14b8854a2d600f4b2b0ffd4865b32b3a1eca84eed9a72cafa9fa98062a32aa60d3523540e09a447d955ee42d9bdc3b2315df9fc761fdf11798cd0c9c04b9f0e4ed3f7f1d9a1f355ca3ccbfa0c4f40175211474a06f82437cfe7e056d2251e1c05afda44fa4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ab299d4646cb2548c36fce27c6a1a57db05cd86af2817810c681283ef96540aaee5a229ffa72e513275024dd227329dab0efa3e443b87e7befc793fcf8d8e67099eddcd957a6adba8b594a17e7709dae7ecb5aab38e8eb2db26715b012a035a4409721a4e3fa641699;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c73fc1e13094276e7df360ea446c9f7c570e5c075c5285636f2d6494f1c5d4b6f55aebc024bc3ce658a56c1238f9d27c08b7be1d07b86fed9215241f8539c2aab4975530a84c7b2d5cf23d36c6ff42109a6586ecccfd09c5f303bc95fd6c3ee30c92f6e3e04bc1db23;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde0857a397d0d9976041668384f004dec8ffa20d415900cc5faad4a8d709c922b2bf129ecdcce2e880a1010a6364502d00c902feb5c0f10604ec18c96d981c220fb0580f3f34697b6953679c91b1d554fcf6baac6c904a9d38baed0dddbd21245259595451c26b39f8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d3c7e956e8d827526a5049ef4ba8eaf6677ff4548a80ef583f05c338831eb479cded793000809443407f8cb65a6c9d607e3a0ebd7f4ea0314714684b687d357198e6f6587612fa7c60131dfd4f4838c9ff36a6379e4b39bc82c54502608e5ed32f94e095d5451b607;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53ed8e453b3de8c2c5fc4c59dded19da91cc8953b80b8cb9edaf292af869995485178e12f8e2563b57908c5767f6cd41107170a47831bff18ccd31e1856e7c0184b2c7daf09aedd41e1b68ce700372bd253d83f77e7b58d638e62e97febcd18ef8f02b3df2e7ba6565;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h159f7b96584c500b65b7c23104a2f54d35d1c0b7c3b1cb19c51dc2f93b33492c0c43762c0b21725ad711d6141841386b20c26c43562a09f4ee9bba84677e648ca74dd95e08a2983d0ea4bda55ad9e6a1295cc80984241f1b414d5073acc5ddb6a9cc3897db660049bb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5b85c524c5e4e9eb4bbf82cf7e492d772e5fd6195d1889c5d4a59c6bf4753a2ea7f05ec13c2b92896a1a9da1c51bd31e4dd9e1d439beca632fcb4c0e0f0fe6b557a4025df49c8c11708f50fccc62faab863ef6f673ea8457045faae8b6d59b6e24f0b7572b37559bbc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183e4cd14771344aeec1dbd0b8383c5b36423e967c659bfbe206f70d7ea656efcd3d754c9374318e84c31adab4f2f6ceba5533ceaad850383a946d845129aed6cf7a551149e23134b2380503bb56e1f945a46632cd42e2251f19beeab2b08b427efa5436aa761f6b4db;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc69da64ecde084731e707d7cecc3548ba54c6ccbd15e8b5eac058eea1f17bb00903185d643385af87e621a68d154d1613a4faa1300a1673c8c4bf549b0f577d0d2c8f18debe0a548b678c353a49ce5ad25a1fa9e059f536d9f67c43fb2c91670c23cc8a747f8f04614;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ad4daa9f7bbd9e8243fa835b321051b3469b5bd6fae958f7cd92c4c0b9e1785e8c88148afb1468ce9842e23b61aec89e967e9cc20c613d16c22e7f4f8186388b4590c6d077237135a124c3761168fad4de8beb4ce89c8c3188fcfdb8c340fcc7295e76530de19b68b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d7ba8328cdebda3a3860db207409506abcb188b0fe78ac17be9d73a9cba0ca049535678ed16083dad107be29cafe7de4b7e75d6ad2de907f03e4b739d2a2907701755a8031600cf257ca6b323a58e09899a08472eb01a034f8f7eb0275900203e96cb4a202488a25b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b29ea584225c9b52af97508d33d5ee4eaf10dd1771cbe9adbae485a04262606454f976fcde252dad5d74ab800716233db5ed90ed87e8e394c817ef572c573acb5212c99c92d827db1187ef1e814ac0a57441537161f342c85e4caec9f3bbd87b574f959cf383d4562f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha9cb11d6ee03730e0a39458cf080c4ea8c17a4745bcda8b08105d9e4f640b82c3032e4d1fb870056acff3842a977815d2dbbaa397247247c4ca2c06424002b018e5c7ac88e87e2bb6a4ae45b0e070ce877d79f25a2392a91895930d7478a48a6f84cf1dc0b4eeccfe4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2a5ea51f6e2b354f4c470c696bd2fd142a0b312bdaabd7af78ada5e3c1e06ba9bfd195a44013de9cb9f2541aaa5fa6496d5afb2a1129af121f4d48af4a2d28852a92f6a30d4760decfac7f545cf9c2f79c047f4b4d81364e73cdb98026137234013894969d72ecec9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95974c2afe33ec9c18a82af18730b563145b73d1186615cba6dd5af525d99bdd777c97f50acde66cc4ac1cef2cb542fd58f26315c5e6f6064afb62cf92bdf0930fba53a0cf94fc40e9346f97439b32c9abd1091f6e5826511aa343363299efcc8d84ceee66d7ab5178;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c56f564ba2357f305f3566e08aff46480364830c7c0e5eed25b2f2ec52ff933f9e0a60d75f4a6e8b4fde22c7564dc0e6b72317412930dfe9fbd8c7e5715298bf5304c1b1efe556c58f5e76031fb52109aa3461bc3f912d891a7dddcf98a4b35b6c2e626bb5cb507d4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h170d7b80abf7469b1f02f6605aed9d36efcedf2c006d45bdd156a48985256d06d32b8c9e061f90b8c16de0d75c0d73498d60df130c48a73538b0110aa06000f7ad5a73dc43097623fd3516f324816d3757bd43bb14db1c249cb013d51cad13033fd0d82006a7b904c8a;
        #1
        $finish();
    end
endmodule
