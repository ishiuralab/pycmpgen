module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    compressor_CLA32_32 compressor_CLA32_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
        src12 <= 32'h0;
        src13 <= 32'h0;
        src14 <= 32'h0;
        src15 <= 32'h0;
        src16 <= 32'h0;
        src17 <= 32'h0;
        src18 <= 32'h0;
        src19 <= 32'h0;
        src20 <= 32'h0;
        src21 <= 32'h0;
        src22 <= 32'h0;
        src23 <= 32'h0;
        src24 <= 32'h0;
        src25 <= 32'h0;
        src26 <= 32'h0;
        src27 <= 32'h0;
        src28 <= 32'h0;
        src29 <= 32'h0;
        src30 <= 32'h0;
        src31 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA32_32(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    input [31:0]src12,
    input [31:0]src13,
    input [31:0]src14,
    input [31:0]src15,
    input [31:0]src16,
    input [31:0]src17,
    input [31:0]src18,
    input [31:0]src19,
    input [31:0]src20,
    input [31:0]src21,
    input [31:0]src22,
    input [31:0]src23,
    input [31:0]src24,
    input [31:0]src25,
    input [31:0]src26,
    input [31:0]src27,
    input [31:0]src28,
    input [31:0]src29,
    input [31:0]src30,
    input [31:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [0:0] comp_out33;
    wire [0:0] comp_out34;
    wire [0:0] comp_out35;
    wire [1:0] comp_out36;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out36[1], 1'h0, 1'h0, 1'h0, comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], 1'h0, comp_out0[1]}),
        .dst({dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      input wire [31:0] src16,
      input wire [31:0] src17,
      input wire [31:0] src18,
      input wire [31:0] src19,
      input wire [31:0] src20,
      input wire [31:0] src21,
      input wire [31:0] src22,
      input wire [31:0] src23,
      input wire [31:0] src24,
      input wire [31:0] src25,
      input wire [31:0] src26,
      input wire [31:0] src27,
      input wire [31:0] src28,
      input wire [31:0] src29,
      input wire [31:0] src30,
      input wire [31:0] src31,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [0:0] dst33,
      output wire [0:0] dst34,
      output wire [0:0] dst35,
      output wire [1:0] dst36);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [31:0] stage0_12;
   wire [31:0] stage0_13;
   wire [31:0] stage0_14;
   wire [31:0] stage0_15;
   wire [31:0] stage0_16;
   wire [31:0] stage0_17;
   wire [31:0] stage0_18;
   wire [31:0] stage0_19;
   wire [31:0] stage0_20;
   wire [31:0] stage0_21;
   wire [31:0] stage0_22;
   wire [31:0] stage0_23;
   wire [31:0] stage0_24;
   wire [31:0] stage0_25;
   wire [31:0] stage0_26;
   wire [31:0] stage0_27;
   wire [31:0] stage0_28;
   wire [31:0] stage0_29;
   wire [31:0] stage0_30;
   wire [31:0] stage0_31;
   wire [10:0] stage1_0;
   wire [14:0] stage1_1;
   wire [11:0] stage1_2;
   wire [12:0] stage1_3;
   wire [18:0] stage1_4;
   wire [11:0] stage1_5;
   wire [12:0] stage1_6;
   wire [20:0] stage1_7;
   wire [11:0] stage1_8;
   wire [17:0] stage1_9;
   wire [11:0] stage1_10;
   wire [15:0] stage1_11;
   wire [12:0] stage1_12;
   wire [14:0] stage1_13;
   wire [12:0] stage1_14;
   wire [17:0] stage1_15;
   wire [12:0] stage1_16;
   wire [18:0] stage1_17;
   wire [16:0] stage1_18;
   wire [11:0] stage1_19;
   wire [12:0] stage1_20;
   wire [14:0] stage1_21;
   wire [11:0] stage1_22;
   wire [13:0] stage1_23;
   wire [22:0] stage1_24;
   wire [14:0] stage1_25;
   wire [11:0] stage1_26;
   wire [15:0] stage1_27;
   wire [16:0] stage1_28;
   wire [13:0] stage1_29;
   wire [22:0] stage1_30;
   wire [9:0] stage1_31;
   wire [7:0] stage1_32;
   wire [4:0] stage1_33;
   wire [1:0] stage2_0;
   wire [6:0] stage2_1;
   wire [3:0] stage2_2;
   wire [4:0] stage2_3;
   wire [10:0] stage2_4;
   wire [5:0] stage2_5;
   wire [3:0] stage2_6;
   wire [5:0] stage2_7;
   wire [7:0] stage2_8;
   wire [12:0] stage2_9;
   wire [3:0] stage2_10;
   wire [4:0] stage2_11;
   wire [7:0] stage2_12;
   wire [5:0] stage2_13;
   wire [9:0] stage2_14;
   wire [5:0] stage2_15;
   wire [7:0] stage2_16;
   wire [5:0] stage2_17;
   wire [5:0] stage2_18;
   wire [10:0] stage2_19;
   wire [10:0] stage2_20;
   wire [11:0] stage2_21;
   wire [5:0] stage2_22;
   wire [3:0] stage2_23;
   wire [8:0] stage2_24;
   wire [7:0] stage2_25;
   wire [5:0] stage2_26;
   wire [8:0] stage2_27;
   wire [7:0] stage2_28;
   wire [5:0] stage2_29;
   wire [5:0] stage2_30;
   wire [6:0] stage2_31;
   wire [6:0] stage2_32;
   wire [2:0] stage2_33;
   wire [1:0] stage2_34;
   wire [0:0] stage2_35;
   wire [1:0] stage3_0;
   wire [0:0] stage3_1;
   wire [1:0] stage3_2;
   wire [3:0] stage3_3;
   wire [6:0] stage3_4;
   wire [1:0] stage3_5;
   wire [5:0] stage3_6;
   wire [0:0] stage3_7;
   wire [6:0] stage3_8;
   wire [4:0] stage3_9;
   wire [2:0] stage3_10;
   wire [1:0] stage3_11;
   wire [6:0] stage3_12;
   wire [5:0] stage3_13;
   wire [1:0] stage3_14;
   wire [5:0] stage3_15;
   wire [2:0] stage3_16;
   wire [5:0] stage3_17;
   wire [1:0] stage3_18;
   wire [2:0] stage3_19;
   wire [5:0] stage3_20;
   wire [3:0] stage3_21;
   wire [2:0] stage3_22;
   wire [3:0] stage3_23;
   wire [5:0] stage3_24;
   wire [2:0] stage3_25;
   wire [1:0] stage3_26;
   wire [4:0] stage3_27;
   wire [5:0] stage3_28;
   wire [6:0] stage3_29;
   wire [0:0] stage3_30;
   wire [1:0] stage3_31;
   wire [3:0] stage3_32;
   wire [1:0] stage3_33;
   wire [2:0] stage3_34;
   wire [0:0] stage3_35;
   wire [0:0] stage3_36;
   wire [1:0] stage4_0;
   wire [0:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [1:0] stage4_20;
   wire [1:0] stage4_21;
   wire [1:0] stage4_22;
   wire [1:0] stage4_23;
   wire [1:0] stage4_24;
   wire [1:0] stage4_25;
   wire [1:0] stage4_26;
   wire [1:0] stage4_27;
   wire [1:0] stage4_28;
   wire [1:0] stage4_29;
   wire [1:0] stage4_30;
   wire [1:0] stage4_31;
   wire [1:0] stage4_32;
   wire [0:0] stage4_33;
   wire [0:0] stage4_34;
   wire [0:0] stage4_35;
   wire [1:0] stage4_36;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;
   assign dst22 = stage4_22;
   assign dst23 = stage4_23;
   assign dst24 = stage4_24;
   assign dst25 = stage4_25;
   assign dst26 = stage4_26;
   assign dst27 = stage4_27;
   assign dst28 = stage4_28;
   assign dst29 = stage4_29;
   assign dst30 = stage4_30;
   assign dst31 = stage4_31;
   assign dst32 = stage4_32;
   assign dst33 = stage4_33;
   assign dst34 = stage4_34;
   assign dst35 = stage4_35;
   assign dst36 = stage4_36;

   gpc1406_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[4]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[5]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[6]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9]},
      {stage1_5[0],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc615_5 gpc7 (
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage0_3[10]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[1],stage1_4[7],stage1_3[7],stage1_2[7]}
   );
   gpc615_5 gpc8 (
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28]},
      {stage0_3[11]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[2],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc615_5 gpc9 (
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[3],stage1_4[9],stage1_3[9]}
   );
   gpc615_5 gpc10 (
      {stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21]},
      {stage0_4[13]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[3],stage1_5[4],stage1_4[10],stage1_3[10]}
   );
   gpc615_5 gpc11 (
      {stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage0_4[14]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[4],stage1_5[5],stage1_4[11],stage1_3[11]}
   );
   gpc615_5 gpc12 (
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage0_4[15]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[5],stage1_5[6],stage1_4[12],stage1_3[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[4],stage1_6[6],stage1_5[7],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[5],stage1_6[7],stage1_5[8],stage1_4[14]}
   );
   gpc606_5 gpc15 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[2],stage1_7[6],stage1_6[8],stage1_5[9]}
   );
   gpc135_4 gpc16 (
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16]},
      {stage0_7[6], stage0_7[7], stage0_7[8]},
      {stage0_8[0]},
      {stage1_9[1],stage1_8[3],stage1_7[7],stage1_6[9]}
   );
   gpc135_4 gpc17 (
      {stage0_6[17], stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21]},
      {stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage0_8[1]},
      {stage1_9[2],stage1_8[4],stage1_7[8],stage1_6[10]}
   );
   gpc135_4 gpc18 (
      {stage0_6[22], stage0_6[23], stage0_6[24], stage0_6[25], stage0_6[26]},
      {stage0_7[12], stage0_7[13], stage0_7[14]},
      {stage0_8[2]},
      {stage1_9[3],stage1_8[5],stage1_7[9],stage1_6[11]}
   );
   gpc615_5 gpc19 (
      {stage0_6[27], stage0_6[28], stage0_6[29], stage0_6[30], stage0_6[31]},
      {stage0_7[15]},
      {stage0_8[3], stage0_8[4], stage0_8[5], stage0_8[6], stage0_8[7], stage0_8[8]},
      {stage1_10[0],stage1_9[4],stage1_8[6],stage1_7[10],stage1_6[12]}
   );
   gpc1343_5 gpc20 (
      {stage0_7[16], stage0_7[17], stage0_7[18]},
      {stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2]},
      {stage0_10[0]},
      {stage1_11[0],stage1_10[1],stage1_9[5],stage1_8[7],stage1_7[11]}
   );
   gpc615_5 gpc21 (
      {stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage0_8[13]},
      {stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage1_11[1],stage1_10[2],stage1_9[6],stage1_8[8],stage1_7[12]}
   );
   gpc606_5 gpc22 (
      {stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6]},
      {stage1_12[0],stage1_11[2],stage1_10[3],stage1_9[7],stage1_8[9]}
   );
   gpc606_5 gpc23 (
      {stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25]},
      {stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage1_12[1],stage1_11[3],stage1_10[4],stage1_9[8],stage1_8[10]}
   );
   gpc606_5 gpc24 (
      {stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31]},
      {stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18]},
      {stage1_12[2],stage1_11[4],stage1_10[5],stage1_9[9],stage1_8[11]}
   );
   gpc606_5 gpc25 (
      {stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[3],stage1_11[5],stage1_10[6],stage1_9[10]}
   );
   gpc606_5 gpc26 (
      {stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[4],stage1_11[6],stage1_10[7],stage1_9[11]}
   );
   gpc606_5 gpc27 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[5],stage1_11[7],stage1_10[8],stage1_9[12]}
   );
   gpc606_5 gpc28 (
      {stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23], stage0_10[24]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[3],stage1_12[6],stage1_11[8],stage1_10[9]}
   );
   gpc606_5 gpc29 (
      {stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[4],stage1_12[7],stage1_11[9],stage1_10[10]}
   );
   gpc615_5 gpc30 (
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22]},
      {stage0_12[12]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[5],stage1_12[8],stage1_11[10]}
   );
   gpc615_5 gpc31 (
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27]},
      {stage0_12[13]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[3],stage1_13[6],stage1_12[9],stage1_11[11]}
   );
   gpc606_5 gpc32 (
      {stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[2],stage1_14[4],stage1_13[7],stage1_12[10]}
   );
   gpc606_5 gpc33 (
      {stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[3],stage1_14[5],stage1_13[8],stage1_12[11]}
   );
   gpc606_5 gpc34 (
      {stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[4],stage1_14[6],stage1_13[9],stage1_12[12]}
   );
   gpc606_5 gpc35 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[3],stage1_15[5],stage1_14[7],stage1_13[10]}
   );
   gpc606_5 gpc36 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[4],stage1_15[6],stage1_14[8],stage1_13[11]}
   );
   gpc606_5 gpc37 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[5],stage1_15[7],stage1_14[9],stage1_13[12]}
   );
   gpc615_5 gpc38 (
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22]},
      {stage0_15[18]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[3],stage1_16[6],stage1_15[8],stage1_14[10]}
   );
   gpc615_5 gpc39 (
      {stage0_14[23], stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27]},
      {stage0_15[19]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[4],stage1_16[7],stage1_15[9],stage1_14[11]}
   );
   gpc615_5 gpc40 (
      {stage0_14[28], stage0_14[29], stage0_14[30], stage0_14[31], 1'b0},
      {stage0_15[20]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[5],stage1_16[8],stage1_15[10],stage1_14[12]}
   );
   gpc615_5 gpc41 (
      {stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24], stage0_15[25]},
      {stage0_16[18]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[3],stage1_17[6],stage1_16[9],stage1_15[11]}
   );
   gpc606_5 gpc42 (
      {stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[1],stage1_18[4],stage1_17[7],stage1_16[10]}
   );
   gpc606_5 gpc43 (
      {stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[2],stage1_18[5],stage1_17[8],stage1_16[11]}
   );
   gpc615_5 gpc44 (
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10]},
      {stage0_18[12]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[2],stage1_19[3],stage1_18[6],stage1_17[9]}
   );
   gpc615_5 gpc45 (
      {stage0_17[11], stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15]},
      {stage0_18[13]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[3],stage1_19[4],stage1_18[7],stage1_17[10]}
   );
   gpc615_5 gpc46 (
      {stage0_17[16], stage0_17[17], stage0_17[18], stage0_17[19], stage0_17[20]},
      {stage0_18[14]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[4],stage1_19[5],stage1_18[8],stage1_17[11]}
   );
   gpc615_5 gpc47 (
      {stage0_17[21], stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25]},
      {stage0_18[15]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[5],stage1_19[6],stage1_18[9],stage1_17[12]}
   );
   gpc606_5 gpc48 (
      {stage0_18[16], stage0_18[17], stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[4],stage1_20[6],stage1_19[7],stage1_18[10]}
   );
   gpc615_5 gpc49 (
      {stage0_18[22], stage0_18[23], stage0_18[24], stage0_18[25], stage0_18[26]},
      {stage0_19[24]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[5],stage1_20[7],stage1_19[8],stage1_18[11]}
   );
   gpc615_5 gpc50 (
      {stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage0_20[12]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[2],stage1_21[6],stage1_20[8],stage1_19[9]}
   );
   gpc615_5 gpc51 (
      {stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage0_21[6]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[1],stage1_22[3],stage1_21[7],stage1_20[9]}
   );
   gpc615_5 gpc52 (
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22]},
      {stage0_21[7]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[2],stage1_22[4],stage1_21[8],stage1_20[10]}
   );
   gpc615_5 gpc53 (
      {stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage0_21[8]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[3],stage1_22[5],stage1_21[9],stage1_20[11]}
   );
   gpc615_5 gpc54 (
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], 1'b0},
      {stage0_21[9]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[4],stage1_22[6],stage1_21[10],stage1_20[12]}
   );
   gpc606_5 gpc55 (
      {stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[4],stage1_23[5],stage1_22[7],stage1_21[11]}
   );
   gpc606_5 gpc56 (
      {stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[5],stage1_23[6],stage1_22[8],stage1_21[12]}
   );
   gpc615_5 gpc57 (
      {stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25], stage0_21[26]},
      {stage0_22[24]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[6],stage1_23[7],stage1_22[9],stage1_21[13]}
   );
   gpc615_5 gpc58 (
      {stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31]},
      {stage0_22[25]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[7],stage1_23[8],stage1_22[10],stage1_21[14]}
   );
   gpc606_5 gpc59 (
      {stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30], stage0_22[31]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[4],stage1_24[8],stage1_23[9],stage1_22[11]}
   );
   gpc615_5 gpc60 (
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28]},
      {stage0_24[6]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[1],stage1_25[5],stage1_24[9],stage1_23[10]}
   );
   gpc615_5 gpc61 (
      {stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage0_25[6]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[1],stage1_26[2],stage1_25[6],stage1_24[10]}
   );
   gpc615_5 gpc62 (
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16]},
      {stage0_25[7]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[2],stage1_26[3],stage1_25[7],stage1_24[11]}
   );
   gpc615_5 gpc63 (
      {stage0_24[17], stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21]},
      {stage0_25[8]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[3],stage1_26[4],stage1_25[8],stage1_24[12]}
   );
   gpc606_5 gpc64 (
      {stage0_25[9], stage0_25[10], stage0_25[11], stage0_25[12], stage0_25[13], stage0_25[14]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[3],stage1_27[4],stage1_26[5],stage1_25[9]}
   );
   gpc615_5 gpc65 (
      {stage0_25[15], stage0_25[16], stage0_25[17], stage0_25[18], stage0_25[19]},
      {stage0_26[18]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[4],stage1_27[5],stage1_26[6],stage1_25[10]}
   );
   gpc615_5 gpc66 (
      {stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23], stage0_25[24]},
      {stage0_26[19]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[5],stage1_27[6],stage1_26[7],stage1_25[11]}
   );
   gpc615_5 gpc67 (
      {stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_26[20]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[6],stage1_27[7],stage1_26[8],stage1_25[12]}
   );
   gpc615_5 gpc68 (
      {stage0_26[21], stage0_26[22], stage0_26[23], stage0_26[24], stage0_26[25]},
      {stage0_27[24]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[4],stage1_28[7],stage1_27[8],stage1_26[9]}
   );
   gpc615_5 gpc69 (
      {stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29], stage0_26[30]},
      {stage0_27[25]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[5],stage1_28[8],stage1_27[9],stage1_26[10]}
   );
   gpc615_5 gpc70 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16]},
      {stage0_29[0]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[0],stage1_30[2],stage1_29[6],stage1_28[9]}
   );
   gpc615_5 gpc71 (
      {stage0_28[17], stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21]},
      {stage0_29[1]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[1],stage1_30[3],stage1_29[7],stage1_28[10]}
   );
   gpc615_5 gpc72 (
      {stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25], stage0_28[26]},
      {stage0_29[2]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[2],stage1_30[4],stage1_29[8],stage1_28[11]}
   );
   gpc606_5 gpc73 (
      {stage0_29[3], stage0_29[4], stage0_29[5], stage0_29[6], stage0_29[7], stage0_29[8]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[3],stage1_31[3],stage1_30[5],stage1_29[9]}
   );
   gpc606_5 gpc74 (
      {stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12], stage0_29[13], stage0_29[14]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[4],stage1_31[4],stage1_30[6],stage1_29[10]}
   );
   gpc606_5 gpc75 (
      {stage0_29[15], stage0_29[16], stage0_29[17], stage0_29[18], stage0_29[19], stage0_29[20]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[5],stage1_31[5],stage1_30[7],stage1_29[11]}
   );
   gpc606_5 gpc76 (
      {stage0_29[21], stage0_29[22], stage0_29[23], stage0_29[24], stage0_29[25], stage0_29[26]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[6],stage1_31[6],stage1_30[8],stage1_29[12]}
   );
   gpc615_5 gpc77 (
      {stage0_29[27], stage0_29[28], stage0_29[29], stage0_29[30], stage0_29[31]},
      {stage0_30[18]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[7],stage1_31[7],stage1_30[9],stage1_29[13]}
   );
   gpc1_1 gpc78 (
      {stage0_0[27]},
      {stage1_0[6]}
   );
   gpc1_1 gpc79 (
      {stage0_0[28]},
      {stage1_0[7]}
   );
   gpc1_1 gpc80 (
      {stage0_0[29]},
      {stage1_0[8]}
   );
   gpc1_1 gpc81 (
      {stage0_0[30]},
      {stage1_0[9]}
   );
   gpc1_1 gpc82 (
      {stage0_0[31]},
      {stage1_0[10]}
   );
   gpc1_1 gpc83 (
      {stage0_1[24]},
      {stage1_1[7]}
   );
   gpc1_1 gpc84 (
      {stage0_1[25]},
      {stage1_1[8]}
   );
   gpc1_1 gpc85 (
      {stage0_1[26]},
      {stage1_1[9]}
   );
   gpc1_1 gpc86 (
      {stage0_1[27]},
      {stage1_1[10]}
   );
   gpc1_1 gpc87 (
      {stage0_1[28]},
      {stage1_1[11]}
   );
   gpc1_1 gpc88 (
      {stage0_1[29]},
      {stage1_1[12]}
   );
   gpc1_1 gpc89 (
      {stage0_1[30]},
      {stage1_1[13]}
   );
   gpc1_1 gpc90 (
      {stage0_1[31]},
      {stage1_1[14]}
   );
   gpc1_1 gpc91 (
      {stage0_2[29]},
      {stage1_2[9]}
   );
   gpc1_1 gpc92 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc93 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc94 (
      {stage0_4[28]},
      {stage1_4[15]}
   );
   gpc1_1 gpc95 (
      {stage0_4[29]},
      {stage1_4[16]}
   );
   gpc1_1 gpc96 (
      {stage0_4[30]},
      {stage1_4[17]}
   );
   gpc1_1 gpc97 (
      {stage0_4[31]},
      {stage1_4[18]}
   );
   gpc1_1 gpc98 (
      {stage0_5[30]},
      {stage1_5[10]}
   );
   gpc1_1 gpc99 (
      {stage0_5[31]},
      {stage1_5[11]}
   );
   gpc1_1 gpc100 (
      {stage0_7[24]},
      {stage1_7[13]}
   );
   gpc1_1 gpc101 (
      {stage0_7[25]},
      {stage1_7[14]}
   );
   gpc1_1 gpc102 (
      {stage0_7[26]},
      {stage1_7[15]}
   );
   gpc1_1 gpc103 (
      {stage0_7[27]},
      {stage1_7[16]}
   );
   gpc1_1 gpc104 (
      {stage0_7[28]},
      {stage1_7[17]}
   );
   gpc1_1 gpc105 (
      {stage0_7[29]},
      {stage1_7[18]}
   );
   gpc1_1 gpc106 (
      {stage0_7[30]},
      {stage1_7[19]}
   );
   gpc1_1 gpc107 (
      {stage0_7[31]},
      {stage1_7[20]}
   );
   gpc1_1 gpc108 (
      {stage0_9[27]},
      {stage1_9[13]}
   );
   gpc1_1 gpc109 (
      {stage0_9[28]},
      {stage1_9[14]}
   );
   gpc1_1 gpc110 (
      {stage0_9[29]},
      {stage1_9[15]}
   );
   gpc1_1 gpc111 (
      {stage0_9[30]},
      {stage1_9[16]}
   );
   gpc1_1 gpc112 (
      {stage0_9[31]},
      {stage1_9[17]}
   );
   gpc1_1 gpc113 (
      {stage0_10[31]},
      {stage1_10[11]}
   );
   gpc1_1 gpc114 (
      {stage0_11[28]},
      {stage1_11[12]}
   );
   gpc1_1 gpc115 (
      {stage0_11[29]},
      {stage1_11[13]}
   );
   gpc1_1 gpc116 (
      {stage0_11[30]},
      {stage1_11[14]}
   );
   gpc1_1 gpc117 (
      {stage0_11[31]},
      {stage1_11[15]}
   );
   gpc1_1 gpc118 (
      {stage0_13[30]},
      {stage1_13[13]}
   );
   gpc1_1 gpc119 (
      {stage0_13[31]},
      {stage1_13[14]}
   );
   gpc1_1 gpc120 (
      {stage0_15[26]},
      {stage1_15[12]}
   );
   gpc1_1 gpc121 (
      {stage0_15[27]},
      {stage1_15[13]}
   );
   gpc1_1 gpc122 (
      {stage0_15[28]},
      {stage1_15[14]}
   );
   gpc1_1 gpc123 (
      {stage0_15[29]},
      {stage1_15[15]}
   );
   gpc1_1 gpc124 (
      {stage0_15[30]},
      {stage1_15[16]}
   );
   gpc1_1 gpc125 (
      {stage0_15[31]},
      {stage1_15[17]}
   );
   gpc1_1 gpc126 (
      {stage0_16[31]},
      {stage1_16[12]}
   );
   gpc1_1 gpc127 (
      {stage0_17[26]},
      {stage1_17[13]}
   );
   gpc1_1 gpc128 (
      {stage0_17[27]},
      {stage1_17[14]}
   );
   gpc1_1 gpc129 (
      {stage0_17[28]},
      {stage1_17[15]}
   );
   gpc1_1 gpc130 (
      {stage0_17[29]},
      {stage1_17[16]}
   );
   gpc1_1 gpc131 (
      {stage0_17[30]},
      {stage1_17[17]}
   );
   gpc1_1 gpc132 (
      {stage0_17[31]},
      {stage1_17[18]}
   );
   gpc1_1 gpc133 (
      {stage0_18[27]},
      {stage1_18[12]}
   );
   gpc1_1 gpc134 (
      {stage0_18[28]},
      {stage1_18[13]}
   );
   gpc1_1 gpc135 (
      {stage0_18[29]},
      {stage1_18[14]}
   );
   gpc1_1 gpc136 (
      {stage0_18[30]},
      {stage1_18[15]}
   );
   gpc1_1 gpc137 (
      {stage0_18[31]},
      {stage1_18[16]}
   );
   gpc1_1 gpc138 (
      {stage0_19[30]},
      {stage1_19[10]}
   );
   gpc1_1 gpc139 (
      {stage0_19[31]},
      {stage1_19[11]}
   );
   gpc1_1 gpc140 (
      {stage0_23[29]},
      {stage1_23[11]}
   );
   gpc1_1 gpc141 (
      {stage0_23[30]},
      {stage1_23[12]}
   );
   gpc1_1 gpc142 (
      {stage0_23[31]},
      {stage1_23[13]}
   );
   gpc1_1 gpc143 (
      {stage0_24[22]},
      {stage1_24[13]}
   );
   gpc1_1 gpc144 (
      {stage0_24[23]},
      {stage1_24[14]}
   );
   gpc1_1 gpc145 (
      {stage0_24[24]},
      {stage1_24[15]}
   );
   gpc1_1 gpc146 (
      {stage0_24[25]},
      {stage1_24[16]}
   );
   gpc1_1 gpc147 (
      {stage0_24[26]},
      {stage1_24[17]}
   );
   gpc1_1 gpc148 (
      {stage0_24[27]},
      {stage1_24[18]}
   );
   gpc1_1 gpc149 (
      {stage0_24[28]},
      {stage1_24[19]}
   );
   gpc1_1 gpc150 (
      {stage0_24[29]},
      {stage1_24[20]}
   );
   gpc1_1 gpc151 (
      {stage0_24[30]},
      {stage1_24[21]}
   );
   gpc1_1 gpc152 (
      {stage0_24[31]},
      {stage1_24[22]}
   );
   gpc1_1 gpc153 (
      {stage0_25[30]},
      {stage1_25[13]}
   );
   gpc1_1 gpc154 (
      {stage0_25[31]},
      {stage1_25[14]}
   );
   gpc1_1 gpc155 (
      {stage0_26[31]},
      {stage1_26[11]}
   );
   gpc1_1 gpc156 (
      {stage0_27[26]},
      {stage1_27[10]}
   );
   gpc1_1 gpc157 (
      {stage0_27[27]},
      {stage1_27[11]}
   );
   gpc1_1 gpc158 (
      {stage0_27[28]},
      {stage1_27[12]}
   );
   gpc1_1 gpc159 (
      {stage0_27[29]},
      {stage1_27[13]}
   );
   gpc1_1 gpc160 (
      {stage0_27[30]},
      {stage1_27[14]}
   );
   gpc1_1 gpc161 (
      {stage0_27[31]},
      {stage1_27[15]}
   );
   gpc1_1 gpc162 (
      {stage0_28[27]},
      {stage1_28[12]}
   );
   gpc1_1 gpc163 (
      {stage0_28[28]},
      {stage1_28[13]}
   );
   gpc1_1 gpc164 (
      {stage0_28[29]},
      {stage1_28[14]}
   );
   gpc1_1 gpc165 (
      {stage0_28[30]},
      {stage1_28[15]}
   );
   gpc1_1 gpc166 (
      {stage0_28[31]},
      {stage1_28[16]}
   );
   gpc1_1 gpc167 (
      {stage0_30[19]},
      {stage1_30[10]}
   );
   gpc1_1 gpc168 (
      {stage0_30[20]},
      {stage1_30[11]}
   );
   gpc1_1 gpc169 (
      {stage0_30[21]},
      {stage1_30[12]}
   );
   gpc1_1 gpc170 (
      {stage0_30[22]},
      {stage1_30[13]}
   );
   gpc1_1 gpc171 (
      {stage0_30[23]},
      {stage1_30[14]}
   );
   gpc1_1 gpc172 (
      {stage0_30[24]},
      {stage1_30[15]}
   );
   gpc1_1 gpc173 (
      {stage0_30[25]},
      {stage1_30[16]}
   );
   gpc1_1 gpc174 (
      {stage0_30[26]},
      {stage1_30[17]}
   );
   gpc1_1 gpc175 (
      {stage0_30[27]},
      {stage1_30[18]}
   );
   gpc1_1 gpc176 (
      {stage0_30[28]},
      {stage1_30[19]}
   );
   gpc1_1 gpc177 (
      {stage0_30[29]},
      {stage1_30[20]}
   );
   gpc1_1 gpc178 (
      {stage0_30[30]},
      {stage1_30[21]}
   );
   gpc1_1 gpc179 (
      {stage0_30[31]},
      {stage1_30[22]}
   );
   gpc1_1 gpc180 (
      {stage0_31[30]},
      {stage1_31[8]}
   );
   gpc1_1 gpc181 (
      {stage0_31[31]},
      {stage1_31[9]}
   );
   gpc606_5 gpc182 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc183 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], 1'b0},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc184 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc185 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc1163_5 gpc186 (
      {stage1_4[0], stage1_4[1], stage1_4[2]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_6[0]},
      {stage1_7[0]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc187 (
      {stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[3],stage2_4[5]}
   );
   gpc606_5 gpc188 (
      {stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[2],stage2_7[2],stage2_6[2],stage2_5[4],stage2_4[6]}
   );
   gpc606_5 gpc189 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5], stage1_7[6]},
      {stage2_9[0],stage2_8[3],stage2_7[3],stage2_6[3],stage2_5[5]}
   );
   gpc7_3 gpc190 (
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13]},
      {stage2_9[1],stage2_8[4],stage2_7[4]}
   );
   gpc7_3 gpc191 (
      {stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19], stage1_7[20]},
      {stage2_9[2],stage2_8[5],stage2_7[5]}
   );
   gpc606_5 gpc192 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[0],stage2_9[3],stage2_8[6]}
   );
   gpc606_5 gpc193 (
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[1],stage2_10[1],stage2_9[4],stage2_8[7]}
   );
   gpc606_5 gpc194 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[2],stage2_9[5]}
   );
   gpc606_5 gpc195 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[3],stage2_9[6]}
   );
   gpc615_5 gpc196 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], 1'b0},
      {stage1_12[0]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[2],stage2_12[4],stage2_11[4]}
   );
   gpc2135_5 gpc197 (
      {stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage1_13[6], stage1_13[7], stage1_13[8]},
      {stage1_14[0]},
      {stage1_15[0], stage1_15[1]},
      {stage2_16[0],stage2_15[1],stage2_14[1],stage2_13[3],stage2_12[5]}
   );
   gpc606_5 gpc198 (
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[1],stage2_15[2],stage2_14[2],stage2_13[4],stage2_12[6]}
   );
   gpc606_5 gpc199 (
      {stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14]},
      {stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7]},
      {stage2_17[0],stage2_16[2],stage2_15[3],stage2_14[3],stage2_13[5]}
   );
   gpc615_5 gpc200 (
      {stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11], stage1_15[12]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[0],stage2_17[1],stage2_16[3],stage2_15[4]}
   );
   gpc615_5 gpc201 (
      {stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[1]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[1],stage2_17[2],stage2_16[4],stage2_15[5]}
   );
   gpc615_5 gpc202 (
      {stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage1_17[12]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[2],stage2_18[2],stage2_17[3],stage2_16[5]}
   );
   gpc615_5 gpc203 (
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage1_17[13]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[3],stage2_18[3],stage2_17[4],stage2_16[6]}
   );
   gpc615_5 gpc204 (
      {stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18]},
      {stage1_18[12]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[4],stage2_18[4],stage2_17[5]}
   );
   gpc615_5 gpc205 (
      {stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], 1'b0},
      {stage1_19[6]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[1],stage2_20[3],stage2_19[5],stage2_18[5]}
   );
   gpc606_5 gpc206 (
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[0],stage2_23[0],stage2_22[1],stage2_21[2]}
   );
   gpc2135_5 gpc207 (
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4]},
      {stage1_23[6], stage1_23[7], stage1_23[8]},
      {stage1_24[0]},
      {stage1_25[0], stage1_25[1]},
      {stage2_26[0],stage2_25[1],stage2_24[1],stage2_23[1],stage2_22[2]}
   );
   gpc615_5 gpc208 (
      {stage1_22[5], stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9]},
      {stage1_23[9]},
      {stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6]},
      {stage2_26[1],stage2_25[2],stage2_24[2],stage2_23[2],stage2_22[3]}
   );
   gpc615_5 gpc209 (
      {stage1_23[10], stage1_23[11], stage1_23[12], stage1_23[13], 1'b0},
      {stage1_24[7]},
      {stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6], stage1_25[7]},
      {stage2_27[0],stage2_26[2],stage2_25[3],stage2_24[3],stage2_23[3]}
   );
   gpc606_5 gpc210 (
      {stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[1],stage2_26[3],stage2_25[4],stage2_24[4]}
   );
   gpc606_5 gpc211 (
      {stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[2],stage2_26[4],stage2_25[5],stage2_24[5]}
   );
   gpc606_5 gpc212 (
      {stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12], stage1_25[13]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[3],stage2_26[5],stage2_25[6]}
   );
   gpc606_5 gpc213 (
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[0],stage2_29[1],stage2_28[3],stage2_27[4]}
   );
   gpc606_5 gpc214 (
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[1],stage2_30[1],stage2_29[2],stage2_28[4]}
   );
   gpc615_5 gpc215 (
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10]},
      {stage1_29[6]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[2],stage2_30[2],stage2_29[3],stage2_28[5]}
   );
   gpc615_5 gpc216 (
      {stage1_28[11], stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15]},
      {stage1_29[7]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[3],stage2_30[3],stage2_29[4],stage2_28[6]}
   );
   gpc606_5 gpc217 (
      {stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11], stage1_29[12], stage1_29[13]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[3],stage2_31[4],stage2_30[4],stage2_29[5]}
   );
   gpc606_5 gpc218 (
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], 1'b0},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[1],stage2_32[4],stage2_31[5],stage2_30[5]}
   );
   gpc615_5 gpc219 (
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], 1'b0},
      {stage1_32[6]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], 1'b0},
      {stage2_35[0],stage2_34[1],stage2_33[2],stage2_32[5],stage2_31[6]}
   );
   gpc1_1 gpc220 (
      {stage1_1[12]},
      {stage2_1[4]}
   );
   gpc1_1 gpc221 (
      {stage1_1[13]},
      {stage2_1[5]}
   );
   gpc1_1 gpc222 (
      {stage1_1[14]},
      {stage2_1[6]}
   );
   gpc1_1 gpc223 (
      {stage1_3[12]},
      {stage2_3[4]}
   );
   gpc1_1 gpc224 (
      {stage1_4[15]},
      {stage2_4[7]}
   );
   gpc1_1 gpc225 (
      {stage1_4[16]},
      {stage2_4[8]}
   );
   gpc1_1 gpc226 (
      {stage1_4[17]},
      {stage2_4[9]}
   );
   gpc1_1 gpc227 (
      {stage1_4[18]},
      {stage2_4[10]}
   );
   gpc1_1 gpc228 (
      {stage1_9[12]},
      {stage2_9[7]}
   );
   gpc1_1 gpc229 (
      {stage1_9[13]},
      {stage2_9[8]}
   );
   gpc1_1 gpc230 (
      {stage1_9[14]},
      {stage2_9[9]}
   );
   gpc1_1 gpc231 (
      {stage1_9[15]},
      {stage2_9[10]}
   );
   gpc1_1 gpc232 (
      {stage1_9[16]},
      {stage2_9[11]}
   );
   gpc1_1 gpc233 (
      {stage1_9[17]},
      {stage2_9[12]}
   );
   gpc1_1 gpc234 (
      {stage1_12[12]},
      {stage2_12[7]}
   );
   gpc1_1 gpc235 (
      {stage1_14[7]},
      {stage2_14[4]}
   );
   gpc1_1 gpc236 (
      {stage1_14[8]},
      {stage2_14[5]}
   );
   gpc1_1 gpc237 (
      {stage1_14[9]},
      {stage2_14[6]}
   );
   gpc1_1 gpc238 (
      {stage1_14[10]},
      {stage2_14[7]}
   );
   gpc1_1 gpc239 (
      {stage1_14[11]},
      {stage2_14[8]}
   );
   gpc1_1 gpc240 (
      {stage1_14[12]},
      {stage2_14[9]}
   );
   gpc1_1 gpc241 (
      {stage1_16[12]},
      {stage2_16[7]}
   );
   gpc1_1 gpc242 (
      {stage1_19[7]},
      {stage2_19[6]}
   );
   gpc1_1 gpc243 (
      {stage1_19[8]},
      {stage2_19[7]}
   );
   gpc1_1 gpc244 (
      {stage1_19[9]},
      {stage2_19[8]}
   );
   gpc1_1 gpc245 (
      {stage1_19[10]},
      {stage2_19[9]}
   );
   gpc1_1 gpc246 (
      {stage1_19[11]},
      {stage2_19[10]}
   );
   gpc1_1 gpc247 (
      {stage1_20[6]},
      {stage2_20[4]}
   );
   gpc1_1 gpc248 (
      {stage1_20[7]},
      {stage2_20[5]}
   );
   gpc1_1 gpc249 (
      {stage1_20[8]},
      {stage2_20[6]}
   );
   gpc1_1 gpc250 (
      {stage1_20[9]},
      {stage2_20[7]}
   );
   gpc1_1 gpc251 (
      {stage1_20[10]},
      {stage2_20[8]}
   );
   gpc1_1 gpc252 (
      {stage1_20[11]},
      {stage2_20[9]}
   );
   gpc1_1 gpc253 (
      {stage1_20[12]},
      {stage2_20[10]}
   );
   gpc1_1 gpc254 (
      {stage1_21[6]},
      {stage2_21[3]}
   );
   gpc1_1 gpc255 (
      {stage1_21[7]},
      {stage2_21[4]}
   );
   gpc1_1 gpc256 (
      {stage1_21[8]},
      {stage2_21[5]}
   );
   gpc1_1 gpc257 (
      {stage1_21[9]},
      {stage2_21[6]}
   );
   gpc1_1 gpc258 (
      {stage1_21[10]},
      {stage2_21[7]}
   );
   gpc1_1 gpc259 (
      {stage1_21[11]},
      {stage2_21[8]}
   );
   gpc1_1 gpc260 (
      {stage1_21[12]},
      {stage2_21[9]}
   );
   gpc1_1 gpc261 (
      {stage1_21[13]},
      {stage2_21[10]}
   );
   gpc1_1 gpc262 (
      {stage1_21[14]},
      {stage2_21[11]}
   );
   gpc1_1 gpc263 (
      {stage1_22[10]},
      {stage2_22[4]}
   );
   gpc1_1 gpc264 (
      {stage1_22[11]},
      {stage2_22[5]}
   );
   gpc1_1 gpc265 (
      {stage1_24[20]},
      {stage2_24[6]}
   );
   gpc1_1 gpc266 (
      {stage1_24[21]},
      {stage2_24[7]}
   );
   gpc1_1 gpc267 (
      {stage1_24[22]},
      {stage2_24[8]}
   );
   gpc1_1 gpc268 (
      {stage1_25[14]},
      {stage2_25[7]}
   );
   gpc1_1 gpc269 (
      {stage1_27[12]},
      {stage2_27[5]}
   );
   gpc1_1 gpc270 (
      {stage1_27[13]},
      {stage2_27[6]}
   );
   gpc1_1 gpc271 (
      {stage1_27[14]},
      {stage2_27[7]}
   );
   gpc1_1 gpc272 (
      {stage1_27[15]},
      {stage2_27[8]}
   );
   gpc1_1 gpc273 (
      {stage1_28[16]},
      {stage2_28[7]}
   );
   gpc1_1 gpc274 (
      {stage1_32[7]},
      {stage2_32[6]}
   );
   gpc207_4 gpc275 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc615_5 gpc276 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], 1'b0},
      {stage2_3[2]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc277 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1]}
   );
   gpc23_3 gpc278 (
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0], stage2_9[1]},
      {stage3_10[0],stage3_9[1],stage3_8[1]}
   );
   gpc2135_5 gpc279 (
      {stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1]},
      {stage3_13[0],stage3_12[0],stage3_11[0],stage3_10[1],stage3_9[2]}
   );
   gpc1415_5 gpc280 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage2_10[3]},
      {stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[2]},
      {stage3_13[1],stage3_12[1],stage3_11[1],stage3_10[2],stage3_9[3]}
   );
   gpc1163_5 gpc281 (
      {stage2_13[0], stage2_13[1], stage2_13[2]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage2_15[0]},
      {stage2_16[0]},
      {stage3_17[0],stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[2]}
   );
   gpc615_5 gpc282 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], 1'b0},
      {stage2_15[1]},
      {stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5], stage2_16[6]},
      {stage3_18[0],stage3_17[1],stage3_16[1],stage3_15[1],stage3_14[1]}
   );
   gpc1163_5 gpc283 (
      {stage2_17[0], stage2_17[1], stage2_17[2]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage2_19[0]},
      {stage2_20[0]},
      {stage3_21[0],stage3_20[0],stage3_19[0],stage3_18[1],stage3_17[2]}
   );
   gpc615_5 gpc284 (
      {stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage2_20[1]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[0],stage3_21[1],stage3_20[1],stage3_19[1]}
   );
   gpc615_5 gpc285 (
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10]},
      {stage2_20[2]},
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage3_23[1],stage3_22[1],stage3_21[2],stage3_20[2],stage3_19[2]}
   );
   gpc606_5 gpc286 (
      {stage2_20[3], stage2_20[4], stage2_20[5], stage2_20[6], stage2_20[7], stage2_20[8]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[2],stage3_22[2],stage3_21[3],stage3_20[3]}
   );
   gpc615_5 gpc287 (
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], 1'b0},
      {stage2_24[0]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[1],stage3_23[3]}
   );
   gpc615_5 gpc288 (
      {stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage2_25[6]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[1],stage3_26[1],stage3_25[1],stage3_24[2]}
   );
   gpc7_3 gpc289 (
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5], stage2_27[6]},
      {stage3_29[0],stage3_28[1],stage3_27[2]}
   );
   gpc615_5 gpc290 (
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4]},
      {stage2_29[0]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[0],stage3_30[0],stage3_29[1],stage3_28[2]}
   );
   gpc117_4 gpc291 (
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5], stage2_31[6]},
      {stage2_32[0]},
      {stage2_33[0]},
      {stage3_34[0],stage3_33[0],stage3_32[1],stage3_31[1]}
   );
   gpc2135_5 gpc292 (
      {stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage2_33[1], stage2_33[2], 1'b0},
      {stage2_34[0]},
      {stage2_35[0], 1'b0},
      {stage3_36[0],stage3_35[0],stage3_34[1],stage3_33[1],stage3_32[2]}
   );
   gpc1_1 gpc293 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc294 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc295 (
      {stage2_3[3]},
      {stage3_3[2]}
   );
   gpc1_1 gpc296 (
      {stage2_3[4]},
      {stage3_3[3]}
   );
   gpc1_1 gpc297 (
      {stage2_4[6]},
      {stage3_4[2]}
   );
   gpc1_1 gpc298 (
      {stage2_4[7]},
      {stage3_4[3]}
   );
   gpc1_1 gpc299 (
      {stage2_4[8]},
      {stage3_4[4]}
   );
   gpc1_1 gpc300 (
      {stage2_4[9]},
      {stage3_4[5]}
   );
   gpc1_1 gpc301 (
      {stage2_4[10]},
      {stage3_4[6]}
   );
   gpc1_1 gpc302 (
      {stage2_6[0]},
      {stage3_6[2]}
   );
   gpc1_1 gpc303 (
      {stage2_6[1]},
      {stage3_6[3]}
   );
   gpc1_1 gpc304 (
      {stage2_6[2]},
      {stage3_6[4]}
   );
   gpc1_1 gpc305 (
      {stage2_6[3]},
      {stage3_6[5]}
   );
   gpc1_1 gpc306 (
      {stage2_8[3]},
      {stage3_8[2]}
   );
   gpc1_1 gpc307 (
      {stage2_8[4]},
      {stage3_8[3]}
   );
   gpc1_1 gpc308 (
      {stage2_8[5]},
      {stage3_8[4]}
   );
   gpc1_1 gpc309 (
      {stage2_8[6]},
      {stage3_8[5]}
   );
   gpc1_1 gpc310 (
      {stage2_8[7]},
      {stage3_8[6]}
   );
   gpc1_1 gpc311 (
      {stage2_9[12]},
      {stage3_9[4]}
   );
   gpc1_1 gpc312 (
      {stage2_12[3]},
      {stage3_12[2]}
   );
   gpc1_1 gpc313 (
      {stage2_12[4]},
      {stage3_12[3]}
   );
   gpc1_1 gpc314 (
      {stage2_12[5]},
      {stage3_12[4]}
   );
   gpc1_1 gpc315 (
      {stage2_12[6]},
      {stage3_12[5]}
   );
   gpc1_1 gpc316 (
      {stage2_12[7]},
      {stage3_12[6]}
   );
   gpc1_1 gpc317 (
      {stage2_13[3]},
      {stage3_13[3]}
   );
   gpc1_1 gpc318 (
      {stage2_13[4]},
      {stage3_13[4]}
   );
   gpc1_1 gpc319 (
      {stage2_13[5]},
      {stage3_13[5]}
   );
   gpc1_1 gpc320 (
      {stage2_15[2]},
      {stage3_15[2]}
   );
   gpc1_1 gpc321 (
      {stage2_15[3]},
      {stage3_15[3]}
   );
   gpc1_1 gpc322 (
      {stage2_15[4]},
      {stage3_15[4]}
   );
   gpc1_1 gpc323 (
      {stage2_15[5]},
      {stage3_15[5]}
   );
   gpc1_1 gpc324 (
      {stage2_16[7]},
      {stage3_16[2]}
   );
   gpc1_1 gpc325 (
      {stage2_17[3]},
      {stage3_17[3]}
   );
   gpc1_1 gpc326 (
      {stage2_17[4]},
      {stage3_17[4]}
   );
   gpc1_1 gpc327 (
      {stage2_17[5]},
      {stage3_17[5]}
   );
   gpc1_1 gpc328 (
      {stage2_20[9]},
      {stage3_20[4]}
   );
   gpc1_1 gpc329 (
      {stage2_20[10]},
      {stage3_20[5]}
   );
   gpc1_1 gpc330 (
      {stage2_24[6]},
      {stage3_24[3]}
   );
   gpc1_1 gpc331 (
      {stage2_24[7]},
      {stage3_24[4]}
   );
   gpc1_1 gpc332 (
      {stage2_24[8]},
      {stage3_24[5]}
   );
   gpc1_1 gpc333 (
      {stage2_25[7]},
      {stage3_25[2]}
   );
   gpc1_1 gpc334 (
      {stage2_27[7]},
      {stage3_27[3]}
   );
   gpc1_1 gpc335 (
      {stage2_27[8]},
      {stage3_27[4]}
   );
   gpc1_1 gpc336 (
      {stage2_28[5]},
      {stage3_28[3]}
   );
   gpc1_1 gpc337 (
      {stage2_28[6]},
      {stage3_28[4]}
   );
   gpc1_1 gpc338 (
      {stage2_28[7]},
      {stage3_28[5]}
   );
   gpc1_1 gpc339 (
      {stage2_29[1]},
      {stage3_29[2]}
   );
   gpc1_1 gpc340 (
      {stage2_29[2]},
      {stage3_29[3]}
   );
   gpc1_1 gpc341 (
      {stage2_29[3]},
      {stage3_29[4]}
   );
   gpc1_1 gpc342 (
      {stage2_29[4]},
      {stage3_29[5]}
   );
   gpc1_1 gpc343 (
      {stage2_29[5]},
      {stage3_29[6]}
   );
   gpc1_1 gpc344 (
      {stage2_32[6]},
      {stage3_32[3]}
   );
   gpc1_1 gpc345 (
      {stage2_34[1]},
      {stage3_34[2]}
   );
   gpc1163_5 gpc346 (
      {stage3_3[0], stage3_3[1], stage3_3[2]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_5[0]},
      {stage3_6[0]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc615_5 gpc347 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1]}
   );
   gpc135_4 gpc348 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0], stage3_10[1], stage3_10[2]},
      {stage3_11[0]},
      {stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc207_4 gpc349 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1]},
      {stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[1]}
   );
   gpc606_5 gpc350 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[1]}
   );
   gpc1163_5 gpc351 (
      {stage3_16[0], stage3_16[1], stage3_16[2]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage3_18[0]},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[0],stage4_18[0],stage4_17[1],stage4_16[1]}
   );
   gpc1163_5 gpc352 (
      {stage3_19[1], stage3_19[2], 1'b0},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage3_21[0]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[0],stage4_20[1],stage4_19[1]}
   );
   gpc1423_5 gpc353 (
      {stage3_21[1], stage3_21[2], stage3_21[3]},
      {stage3_22[1], stage3_22[2]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3]},
      {stage3_24[0]},
      {stage4_25[0],stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[1]}
   );
   gpc135_4 gpc354 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage3_25[0], stage3_25[1], stage3_25[2]},
      {stage3_26[0]},
      {stage4_27[0],stage4_26[0],stage4_25[1],stage4_24[1]}
   );
   gpc615_5 gpc355 (
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4]},
      {stage3_28[0]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage4_31[0],stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1]}
   );
   gpc2116_5 gpc356 (
      {stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5], 1'b0},
      {stage3_29[6]},
      {stage3_30[0]},
      {stage3_31[0], stage3_31[1]},
      {stage4_32[0],stage4_31[1],stage4_30[1],stage4_29[1],stage4_28[1]}
   );
   gpc1325_5 gpc357 (
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], 1'b0},
      {stage3_33[0], stage3_33[1]},
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0]},
      {stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[0],stage4_32[1]}
   );
   gpc1_1 gpc358 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc359 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc360 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc361 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc362 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc363 (
      {stage3_3[3]},
      {stage4_3[1]}
   );
   gpc1_1 gpc364 (
      {stage3_4[6]},
      {stage4_4[1]}
   );
   gpc1_1 gpc365 (
      {stage3_5[1]},
      {stage4_5[1]}
   );
   gpc1_1 gpc366 (
      {stage3_8[6]},
      {stage4_8[1]}
   );
   gpc1_1 gpc367 (
      {stage3_11[1]},
      {stage4_11[1]}
   );
   gpc1_1 gpc368 (
      {stage3_18[1]},
      {stage4_18[1]}
   );
   gpc1_1 gpc369 (
      {stage3_26[1]},
      {stage4_26[1]}
   );
   gpc1_1 gpc370 (
      {stage3_36[0]},
      {stage4_36[1]}
   );
endmodule

module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [36:0] srcsum;
    wire [36:0] dstsum;
    wire test;
    compressor_CLA32_32 compressor_CLA32_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1adfacad51ea8361e9eaa04f3883a3e9e913fd8863413e5b3c13240e393125b63ff843d3f69b225d1bee71409822ff71e5f6e57b77dc36c7f9f1d52b304b72b6c3ef12b1b1b17d15518e22668b4b0043521490669f36ca5e98945d9c93f7d226d48b5cf93540bd17ed35e4a1cc765486f4f8604a4ea4d9b1723df49ad562138e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3e9b5366cbf90780e4fe10e035e9594d68b5cc8ecc7f1fd2c7d48cfa83d23a15348a5d62c006b04ba5eb191819b387223520d7de4fdf1e8cb0c34fb1b57cfc4e14a2789cb2379dcab1a744d245b2808a64e027235388c272f27bde88411f0152fd788bd1a83918ff9b637f61f84691ce4bbf6c57cc012ed9e0fa109b634de4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7a7ba0a741c2006c68b6a511d573f3084122ad4a108def7f4c2cfd212cc88f42a4e3ee878d2faa322ec80230d0596661423e232d819c11745006d37301603d4ab462fa6a44fb99831c77b9de12d922b06e4fd33a8e47fc5fcb729b8c037280c1cba71b0dde5ba5b1438a871ea65e363e34642e1ece7b64d69ad7a8fd30c50dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9ad120cff3851ac35712c4cd61674c57e273f768b2719ed714486bec4745a22a835f36c1737f544dc33e8eb17368591ef103402b96b8c0bec7d7610dc2a683497ecab6d298359a28a8cd6fd445d007e1431e5741197636c3c3f537c0fca86eebac677b1f3b3270cb5bf5d17cc3507540a829cee812aa30627491154e1b4cd15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfac6f67fd3e92df501994320fadcd7b607d1329d7ac1b792ec5defe08b76aedd3ce8194d487a7a0d84273e98dec70e11046a26f5868a8c13f2735f9dc005a9d6b24c7c88610c29eb43e7dd6d1608b47cc5495acd3fb8f12812af0b5df9c2c5e0e46b1ef74d0d3abb00617e36f3c9c246966d3ad67adc8639afc48250e8ecaaa9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fadff39c9ee3c506aa1c0757ac9d95e1f52cc0834a0775fc3fb9087dea424694d836f32f567b20214aa3467b2d043b53ce665943b0c0f32e123f8084623e1d38a132c1d530246ae64448e9b701fc5aa77e7ae6eec57cd8e113504a9897338a3975566fdc3e3e342ac6a5955b3b3564799878ea4b1b2f577bae010dadafcef84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e9968a2f2e3c21454ae8a1cba89904f0b3d3fe91d1e1e6c9f9fa83f650c6a11f2c3ea92440177f6c7b639ff53ff968726306ae9589ea6a52c37f881edafdab2894790579ff52777af892ca1f1a03558aabfac810e9eb775dd412173610e4b41cbbcea32c6af6f7d25922bb348b30f3cad39e9e64587004189ecf852433832c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc552c20c40b5c614e7d4877cb4096b11da19898da66143fb36a4bdb6ab92d8ecf3aa96b8b6d710f3555c5058772062bb65090289dc3132a16fbe4423441586cab8a2c19de1b2ec8ab6825e493354aaec3bdfce3e556e9d567632fe45105569d89e796ffab157fcb86891cf5d49db57a413eb182936312f9f072776f204a64f19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h568f6f918204e27b83a1c43c2967b60d8bdb0913366a147a97b3f2fb16602c72a9accdc6d56f62adb8c3d628c034b2459f40e94190b4a623f0a60740845c4b0009f2760bfedb006f6062d5cfacf4c63a4946f406fa93d75d6815e8d26156a9fb406499d7aeb64f805f0decc362b8a4191d99592852380ec66ed9c6786a882e67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h857a3c19aecdb1f73ac827b3c22866d6cbe173223dc8b892581918e1e9afc3b1f37a3d454da9fe07552e7cca6504cef2ee7b4f5be068340a98fe739eeee3f60aad9e91afae34ad9cfa65f412e6f93c5645b664395b0d90deda3a211b9a9aa1fd2056400a95f8c2786374e6b4f0520005e49c344be66e574817e51a1373a8e7c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55c857fceea4d70cc5fcce5b7fc47fec5b433619de7ce2769937b65b5c912d9f570a2cfc1c7c5086004e37384606e04808659f7aab465eb1569cb66c72338407a6c054d78f6a16b373cadebf00197b08d79a7794f221a0f670228542270bcfc2e0658293451a7cedf8a491f81cffd98f1959a7bbf597bd949a094c316312f749;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed97d180842b387b9b2c1c64b8a843d07be90351ac4b65d57583a31046de953bea353ed788613a1cb48d77138069be1f59d10c9dce106470ae722d8dea2ae4b12aa6f611f2b77d844fb5ef7d783daa579304cdeab76418908069dd9524d70043dd32fcd2c3ad6984f9fd0e45edb531ee5a608aa814802ce81438b29d38d1ec53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h667aa3fb8a1193ffdeb7206c7b559a5a9e013d85e49068d88900b5b33f253f35fddb92b8d94c7dcd4c91d643ad4c00d9f1d8f206a751353080ff2e55179d9ed853c7fb7a997ff4c02d1c97af5fd4fa6861e674435a02073baaed6942c8973c22b25a8f0da4af53ccc8d5878754403e1be6604314b784bffc696992bc9007a1b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdce4b6cb21b1899965d4ef36b40d04b55eeab461c9968dc17d9f4d0dd8085627e720aa9e4f20d65d2b59cec339f272b3b5c8964ee249ef584e1e5fdcbb2cf39b921a4c51d4d9933d4b76be8169576c7c64aa1551863eb936261392203a376931e5d7674ece15665f4e11bee4eb2ac5f02de3eab00bbc71217306e773ea4abf69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d5a5d23bfad488bb146f1c75a12100e9694c4a61010b83e3385cc45c9c8fe1d366c57966efb7444791a88a03be285b82c5fca478d4cd667923c69921d50f306a8ad5ba7bc0be78dc56909c85866faef658c126f92ab06bf88202d2926dffcc9afe9462194cc9b34c7eb4d27c3df2d197b435c983626e7b57766cda6565bec15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd222a5cee9d891750bfb8c5083417dff875bdf45c08ef93382908a57937fbde06ce281c04bc79f2a943c3646fc0be519b02fd5bada9f9944eb11f4e3dc4c96164206711176cf977282d3010d354460ecd0b28e463a1a51a78d9a61f45fb8f7b672fa45d74f64c4cdf1760a6a5c7aeddc09223346c8c1c82eea9e8e6eeb3d670a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1022a6eb522fe51dda07bc7243057236b3a846a1231b29b925b9c3e2917b882dcd19cf192e41d946a06fb499d7cff77fac1c19a6df0dea477ca75bd87d27a0d5049284b38c4cbb36bbcbf9238cf8b167f1c4cc040696e511a65e8384f8f37a5209df1b532dfb70d4f7c93a061b27c33ef031e86dd61d8414f596bbc8f3c13160;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd787a57830c5b1ca748101506e0b289b7afa94f93f466c946f236e1b3164f4f133c316d5ae1a37818f888db0ee490570899fd40f64106795505ba6c2a8e57cd2a0792f6b36cc908b41cb63bea0b18530bb0a1c7ccc525377924c19458d446e8089681f0abdf7d66618f077f58250d16b50fd5ce876f7cb4529aaa41fe6a4c130;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40d6c2578951fa43db2031c8d94d2ed35a81e2e94314258a49cb1c21aa17d2b6deb47158f15efeabea88147362b9593a0b0c22703d40c52c5f5f4189827b4f58d529a02aac2b151c8d92f4449c13b46d2645091feb0f6c57ca2d726c6037771b584c62462b121752271bd8bbd13648cbbe9ef2d90ab235a871db0576d4dc421a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h988072f6d3d0e6c3c3dceade928c2114dfe87fa1741116e87c3592135230315935da5509919187576c8c235f6c9d50d8df0792c109b79dec473377c851166ab048195a307fcac981410aa027483640051bd26b66a8ad413a741815b9ab3c239469135af4b7b6dc399358aecae1cf79d8630098335123737984a98dbe8cbac6d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84cb4d93b7ed8b258ddfe38049fae3bca657d001c6dbd3c6861eb84fb81a07e13897d62398cddffa250aaf63789d1636755bf7442ee7fcf8fda7ab0f7c8e1c86059fa6730ef5bcb74c3d4b7a9d4fac0c8c1c982229acbe34f05831e583d9dd8cca3c5b75d7af2127a4efe2a2732375dbb6a908f76a85169ba4cd08a9b41fe27b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h328996f1c0857cde862beaa6a56fbd006e503978b4cf54d2b24b94c823a8588418501140af84faaf7d2558508e78033293667d08b87c106e64322f75de578864869eac42be9189f87920625300cccfa8f31b3f4297b056974af7cd7c4671a102a3058222a5bff5fb0c163bd317f4f05c9b4c6e056775c5ed5f6946e53d100227;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd98c30e08ebd1751c2ddee9a241c98f0396b0b0be39f0b408dd3fa76df2bd9c6123c35ce7fedad60a99f382f780f6c8e7e1e807dca52ee5cf24bb5f942e2448c4e0852d0ec4413bea34e3d43b238f8a8d3c9ad1d4a621c401ec7bd119e702a4709179304d05803812d27247ea932372c7fc68989879897fa16517fc765b547d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6456439cf478cc4ca973812ca2cd70ece703041fbb82bd4b6ee83f9b8479294a24b8e920a1a7c957bd2b8f8a2899c9a58f152175bae926c9fcd4a7c38ff2536271536ba0a8dbaeee8ca6827b281844d84918edf920ec69ec7aaaeaf52bbc0e675816e6c04388f9e0a4ba29124a5171769a20c42c61f993a329bfece67d84e67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h522a609f20bbd98ddd219c85ae018c2f96ea2fd399f06254cccb2ac70713d8d35c873a9dbc6f65d72751b8ace3e7f677915690afd415236731e25c0bce673eb9b6f3fd70889cc8c8a72e89ee2cd82dfd77b5963768233857d02233551e84785bee809ceec3ba65ac693f42d8a86e501fc3c0ce86232f0da92c20de1d18a0427c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14ae7a1a448addec5856bab4d52958c1553a972c276e5f43fc2ee7ac71868c4ecf1d53a235aa7163fc94df3c03bd80818e226ab79e71c3290af0f703aaa48abaa6ed8b4d9e684f16a7a2714f3d4127642bbfefb8b53676d0df6e71dd1db62da8f57bedd70b25041b3ace96b9c853c7c4acb516b495ccd0534a7ce8141a413ec7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h241f7cdf51665c975b7e77b6a01696612ee54a5eb51cdbdfed48eb275a0487289a8a617fb9ed520b7f95c759dad887242262ccf48ecbf9cc8c9c63ce65db5277544e1785acb49822428722d06bd03779c4f6f6a88ac55020ad910471feb1f47d3ca1fde230d89ea3ee42f8308cf38820db4e6a06f64c99f1414954239f3bfa4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cff4cdfa54f30c65cc701b377470ee564515ab64e313f3decb451ce2e60828e4368e9d61a5b0562896d0b0645e9d6643179a16a5884b80f4174f741e95d868d6d3638528555824791cd164e595564a81cc4cf34b31d2c1c1e74823fac54e29d0bb3e0982373cb288c58261830aa2af923346460b8478e0b4e455238b527fe65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b4ee16251371d8c414ef232816a30330126d0a45febdadb90b1cc617c02c1a6121d11c3e4b4c32b0b677d8c0cf60af3bee83c3c9e4d3121fdac58720801dc0d4bbcba8c06826ffcea0f011602261e8332474eedafd98edb9557a6e031f64e0b24e62324a49e507bbc4d91fd6edf430f81ab884ee3cc06fa798006404e167642;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87fa9041f4901f918c1340b363e12f6684e8dd0a788b65551d9cf6196e211eda610f3e4691cd394175aa5926f7bbc0070084a8ccaf99d924d320d2b97848afda3c312ff79b79bb4142e41e9cd1721802d4ece971fbc34d3b5c1442588d4b5ecb75e0ca33bac16db86839b9a254a80571754a5ae61848f40c06014535e953e115;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8a31d422c9053e428832da5abb1ef0a7342068bc2ec89470178f7dcfd86c16ccde981cc080e0e2abdc182ae7b65089cc4ec483d1c66c503248a8151546d80268aa8a4bfad4d2cbd6cebafb79ecceea7351de00252ca3bd0431c64e66d3398d8967e9d2408f013ee8e013ea53b66ed1ddcd64ad43b5ab4e5806140fa3b6d80bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fba7aeeca5cc5a615e35d393db24e77d15fc15bfea90c8f2c5dae085a238ebf7b39963c8231f631fd646042402c69ed73b9896a3b4e4a2cb90d2f729da70566cbaf813340cf7d6681e592254b08431ac9ac5ed82ffc4285fdeae422697abae93fdbab134d833c832fc141b022a7b660f7a056c0f97d3c80667c970b85e04a76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3fccfd9c001e5d554a7e2ca2fd73f8740b82aacc245cd0897f8d7c42000ba2a2f932ecc772d2cc32202c67c81d377a1ed074eb7d5ed064672d17d7ae33c7cf489b4ef54c23666a1d79eacf0dc0dca0ed33148167f65b9984bc82e1109d64441b740a7f00db753e634bfa7beffc39934dde663be1e4e4c02d3f13e433b7c8719;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b1d2e996b225ede54e00ed6bc06e3c1d695f2302a2e674794728a34882451e861387bcb46a689582d515d952092eeb6ee638cbaaa6bdd054e357a28e7ed8000b467b8aaf0ee881f745085ca4592303368be6fd7ecece9401c76ed3f1c3bc99337b299c31fefc3a68299641e544096843a6518ab86b4d4a89476f1759b4254dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he862d57f66c848d21a37bb25aba6428944cc9932f631196b60f9e48cde4642de780b8cdcf25acd4f5292aa35b52d5364852a0db1787a253e114bde3a19b1e7424fbc887f74602649020cfe0624982de87c7bb2a1793d03513525f65c4027003f2714c8ae98a5b1686cfda1f4ef46f1b60640534e939bce4f9d945fe112440b5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h586015c0f2c2cd64eb8db35450c71561efd45a8723e3f1be343dbd130a1c24a8297fbdf4d0948bfaf377ba4d5bb9b696b950a85a8492a51d165564a656e6af692b76b72b769ca6ee9ecf18e5e47801e4fb8f00ef826bb5149c9302f47289ea3369acb15631da9ec5948c22101c4af30a65de391b69fc5450f47db6d9ea3cf8e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfeeccb7abffbc64bb168fec032516ada19c0e6f30bce17885d90a87345e0b67192243271ec504c882971ad1cb9029cfe4f6b405cefc5a8c11acf091102eb6b264918c9cf5e7fd41d7ca746d388cc7681e266d16bc0828b024bdefbd141cebaf8f840b1091dacc96b761fd3ae27072b1414cf93bf2d41c298751ebe06871d178d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc22444f7de89ac27a1e582d9b33cf45f295bd6a908665290ff38cb167483453408cefb0482f15fc2f88a07f6618c2bffdc0c7e7fe4ec6128cd31927e203ad60ffa2f7a3372288073290652ac0f922c8cae18dce7db29fafc373bfe8858dee835575ad11e93e88232a49c8be1ef96c221906f007743ea3b5ccb17bbb0371092b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11de320b738495c54740dcc7b2d302a5bcf412dedfbdf551fc85441ce188e0e352bb7e19f894f6274db7d82363e19316711493bd9929a80cb2e57ab5fbffeb10aceea1db39f3b95569492d52242c618f9c26e229a6f1b3c7ec6df873b1ca483a8a5469ab864292cdd684afb9e0d33a30ab118d2e758a1a7a8da0a2206ca8cfa4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1db5f6154a851a2c1cf1f64d9c027be3844aa11b7a6b5d9d58b6b210467b013586836492dc67842045ed24709c6bf7e8fcee2b113b3430df08d2a5fa69922cc313ba05d7f7c6c2b15c7725c856934bde32e9791f3223f033423423700dcdd565cdffe30ee73b3d161caebbbb7695b72337dfe39bf0ec4f3658fc9efc010a4af0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a248ce9482a34651284d37a319122c091b06042885509886e0cd5a802680629ac05faa2071c4f2a4a9c352f4cbc39d9d541ae37e34c8b4765005b7eb4038bfaa33c833259ac7bc9627cc65c9b4cdc23ffc71c87f00bc98c0f8eeb552db0ca024e107f8a463e9a754f9c971f4e88977a6b87b51c2f401cb1a20ba0399e5a462c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cd0fa7c6ae9341994d1ab015759212fd68b818a38ec89a4cf19657d2fb92d31a219866141ec80890183d18769d794484d478d6d3e51b2f35dc61d83065441f4b1dafd7589f766c60a123987790ee8a6b553e5519dd3308260f0bbcaf1ec10bc4d1c9a832ba7fab3dbab4f0b24c50dbf82c2ff1dd10fa6469706ea9830011c60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2c599bd815a3845f8cfefe6978314f4f53ce0d00021b892ee03bae0c1c83198ce4eb97d8fd80b0c3d31813df78d399afa59a5db66b0b944378d6be68431e843cdbce5f900badc8cb1e73d8af3f8ac3f6f910a48c71b1a8af201730669efed934fb41b4b27e6417e07c2bdd7a8340edc3b988dda76dd228356ccc32655f9345;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77d72bea7b560f40e0d223e2d05537d18ccc4165597be8e66073281bdf3ad625a9bc427c3a14dbb38c6887a553e8bd667b90a0c712b50f15c6f373b88e84a01b1b60c927e02d9d7dcc7c770f229582db34b5bd5eb37596c2d038a0cf7e2ccbd3a390397bcf4ca80afd10e9accf1289a5ef10a09677f5bf6aa8b07abdc3cde935;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d80c2c507663720137dd09a8e980c5dfd5ce47438c366ae11ad9497f59c9f82a8a7f3f9eaa9fa67cf5676313acbe085820b294a196ae53555bb1d0cd4e8b30a0842d0c47bc809b70858f33060af3a914edb87fbbca74f18f9ac6a95bc795e681229a954b71823f99567c5a405ea61bf59b7afe2a63c5d7c726da662cafe1167;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3cba1aac33d020116353628745cbd62d1c422a89d3e9f8beb4e31f25d4f1971f881f3771df5908fa8a64a7c7ddd5d9a111253161b3fb6c8533faca61be2555b786a431a997334b93baeae7ca3ac435cdf2fa9365cd67619857b507446d21750d315c468fa025b3143a5e7b0e60018da815fdfadf65f87bb35bbd8c7a9f86fce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a28ae186b2417b8ef53f58b16ec0b1b1e659dc2fdfd080e9e25fde86b112f5e94647c8c3c73cbbd6edb47802f9cf320abd40ac72b26d9f1ee415cdc0b84204df86ef4a44da80d21144cde83e9ef657d1532e6ce841f9ed44665d5a2e63843887e37288318239ae54ff103c082bd1b3287c3f93edcda7fcd2386296c760c79c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he35e30d697d15bb8526a685e2a4edd8a8fb0f4b7c853b8a5f340f9073783866c0ee97f0966030b986ff16dd0b684d387ec6093e39cf360db8a14ee7d7e7d475d24e56ee976fcf3d4ce7b11dbd616db7e708dceff95ee1bdf5e8d43a32e87c1616317b321983055eba2f2ed73634243f4576b3a4f1ae206b0f4bd00521eb6fa22;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54bdde1a4f4cb8ec5c3a7366627590daf973c8c5d793321776db3d1ca4bceec01c2bf87765f2571baad874d934f661ad4cfb4886da00ee6fb514cc6cf359ec718ccc10b4e2945009bfb8c417a4ec9287b4e96b65876055bde728a8623f09ebd37632e4756d75ff9f42f41319c40b912accc7f1422ea66edaaf44fde64ef814de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b14243d826ffa32302e928813989902b2a38670688ae7efcbc19aac8203718e610282ff5d0d70f3e9509f85e9989e1ae57325fc208a454dcfcdfcdc0b3854990d0bfdd1dae111efbd8f3da4d2eb145f475270abed00860a8b6784f5127b04f6d267ee9c88cb8e7607c31de2789083ee78de923f1d4514932a2e7f625d42ba37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h102f7c83770fccdddefd4d45b04794a25ee94337ef8431f8a569d69d9adf23eb71e6eff5a8cbd1b1652fe09fecef926bf4662693c2cb7a8991f6611b9b3927bb5b48736303ef98d8e294d8266ccf02711e016cf673ddbfbc0f400f4061f75e33e3b2261668a7d0be438b0c01a76b362dbce439e4f7b60b76bb9df8dd256b62d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h757de323c88c5ac83092bda1d43e6001b4ad6589c0972f4857a138cbf8f33bd28f59445d68576f2eccebc83d7440d5a0c02af9b5fe0f9c2678718a82030ec8fe5d7835aab3ff4704715d67bbc79a50a8f29b69a14afdf1036c9afe0ac27cc60d01ee802b61b6ad1717c2df0d386ce9bb34397a0508055485c69fabbb350c4e2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38e2c0a5873bb39f1dcb277918cbf28a4b2489ff95f4d6f526d04accae9eda285c55d00d11fbeff89304629496cd6a4b18acd466f0e2850a91bf41c0a0abedf7816f544fd962e2740d786a8a5cf283edc6464e41a0bef5d706be2bb8d001a909e22e1e0e47a4e5089a5e30b5fd8a9848a4628acac4db72496d6b8a14071bcc35;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8548c3886d16f141a5fdea49f77f1e1b8882a1357239d4e39fab9bc8c7b4916033b825c0fb5a4b284917d82dcf60ba2cb2abe370c9b80dbe103de76214ad085375ae4622749b757d2837b5729a536506a20017b740ad281092d79fc4a6593c409ed4a052d2ff14f9b5ccdd23c2b3b6891cec3ce8dd95d1b40860394d57233ac8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11d8ca476a4eed79e3f0085956da162b79fcfd30c7d38cd3f25a0382ee4231324d6239394c8129eaf2db62c3845eacfeaeb8437aee97b7d9e400ef75b25895207f2821dc115f249d9d34abee457457d1b956ab4e93f05af009fd63c2c4a8d0cc322c9caf7d067a3a0b8bd115dd5b3d562f481c3d4914129848474bf6e08e506b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26bbade3ff8fcb4cc400273a1e80c811aec9182c55a5be3983be61302bef714ebcb4f6d615173126b53ba0ee01d286746a9e996a3d41adbd43450fec51a176847bb2659a87f80354ed55453c13d9ae1cb66ea2fd33fe7a209b8728be77d631b46b31f61f2eed9b97fd87c7f17850a4a42179279fd9201c9f43301edfdcfa497d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd77fc237fa357a56494307d0ab52df2e1f8ba6fde112d27f9fa977aafe5089f30119ba86e44ee6be4feab972449404bcc7894f22cf524efb98733a287e86498fe2de93f90138e264cf43f6f1b012339a28a22a4761b41f9a5dc0ec22068dac0cdbc9db909b2ba65c2421660d400f5c6df4985869c9d1c28449fd16330d3f59a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h609d62343521270d9c4c47883047a68be30a69c4f895d1402967ae2263e997b1b14c3ab4eae5a545e3c455bc2412bf5fed02cee13bc2a2e18be0e3fe9aba3b4a7e277d65f50547efe3a51521f06ddca33b992c5338277be0f55cfbec3f853725c7dbc44529fa4cc29a15e25ac3366687c515baeaca07349299feb8990089edfe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf84721a1fbcf671270eec901f781e67d46edb964db39f87c3173df65e242097f3071bf1fb98ca982df1b8e6eab8cd7fd1eb27d6a52de7cd7eb7bacbda9fdeb212c8e1c522eefb5865fbe413916ecf9d48e64ede249d29731d9fb2a3c83ca26f9947b273e13ac501d267555c67c852e851ea8538e260d689ed1e836f2f6309912;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7f72cb3485e47fc66de71114f9a89e2c06922f53bb301fc53bf4d1141a0045ec34d52aa1870349ee8644715356444d3af619720c06f4f74652c00c2f889f8e83b37b20e213668ea6c2fa37871ebdaa0c6624411abb6a4dd6f113c18cd102cad206c7a532ad0e9e3375ab9f8487b4ab58fdbbd1a4139f72a63e3622100a1b868;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b4d2d2c157e31a14727c91f56f743e597dd9f14472fe0e6f4f25a3a54db81d7f063bc5ed04dace51b82100ee6df76eef039140e56686bd553009ba1eb56181d42742ba3a4dcf7aa1479f841b7d39931afeb76e77d615c386e602148eb660260290252dbd54aa3f7f14f811a7abf485a600fbfa77c1f2a20fafebe7f75fbc80a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h693003d2d0444d6ae8c622e849047e4e6f8e20eb40b140d9e1e65387ffff25a2b634b742e7c16da582427c0fc588c833ea91f462315e8258404d6ca179da847409df5f30aad791bf7631d6dbfec037b598b05fb650b13f09d82e11db0747dd2d5c7cb856bf6426a68998a12597f43d1e8ec0318585d22cb4fa7d49ea0850fa81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdafac8896f046c24b5742c0bf7b9d9524a237ddebff882531753abb97c3ba6b00a50140796684eadc1db9338801104b3668ca3f3b2c3b25793d0a50db48525359e572f8657920440acfcb02e0d1469f8346ad4fbd9dae51472dba727b7e30ca13839b6bbb89416c69f3d2b543e6a5d42df1d2cc3e19895dc2e172966c975f67b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h217f80dfd5a0422ae257a338088f5fd1838477c1349e07b9607dd0ede570907fc0030eaad5c797c4e6a59018a69303f399e85ddcb12907d85bc469b36be5df4f910dc20fd0641b7e67dfeaa03ea42d6c835cd9bf27ae2fe1354975d3109b7631934cb37bf10a3af1272ce2441e00de05eb8abb39a23662a4494f0c009e14dd99;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc72e2a30fb638f61e9490409fec387806ec7ee324c78036ac3e507780fd2c9ed6c76cca79610b1e2b52e31e2e6d9505f66526f94a19a42c8b9a19542fb83085188ca95f8a3ea5e8677a069ce621e9f179a07a201a04e18393a180599d9bdc835a90fa5e13a594eeb9a35c9975b92afb95cd030c5afc5ee305a44a3a8186c939;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h837965bd5150fc1c5e0b7c0f31b5e67a7d6526527fa58a439f3a6605ce5ad6ad2ecdae130434521e10dfb4844613242c0b5d8276e680ec5aa5ab52a4b57e531807163f5f2c9a2a4a063afbdc4121ca8386a391efd4032057b3d413b66aa9acef1a2db532960338157a602f2cd75416532cab1f9d9ae5d24e9e86fe1c0d133c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9733180c74660b8e245bb681adad6de89ac1c93c7286314f174bcd6bf38e5347b0c322005c075a1e4c5874d2f03ac56cb999face1940e3937cf21934bb8ed5af85a71720b5b0c2a4650ddfe87dc58796b750a23764ba1bcbcf45712ba2ec5ff0a1e992f22ab5b39bf90a8f9b94d1bf702eb502a2e663a9567099884af774177;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ee573f88fd4f36612263e7ecefff5090a7d77edfda83540ddebbe0f59926d5a64bff7e200fea7d71e57aa70e08ef9c54b3a212e299c90dbad3fde8dce602bcffa7a4ad2833441be1af95903e156cd2beb916976288f20eb93f8eb64586b3a561c45a03fe2ddf01a8343b0602a4118d3faa06ae3e0baf7799b4b3a0097d9a400;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12bb62470b1f35d0029ba089638b12359a34fd631299f91e911e9b6e7d5690dbf8ceeca2a9e7c346feff70adf8abd9b8b7fe8ccbece2dff6dbd9c9a00ccaa9368aae0f8632a03ea07b88428801cf412ec0fc02c48f9e3948124ecd041873b02c4d3454e949b3130243382ac60d11c87f50ca3f595871ac048802cce76332871;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3351219c95f13a019a27f306294a9a0ac3589cad248faa667f46c1152530bf2c5ef8b444d2089cb82e60d7932b22281f4a46a32958d77e2f4124adb544fd80f0c07e7e8039d3988451f7d0a494b85d04535f0154696a8a43ec643b6b29093b688a19b98651027f30e02c2d5f49f9d86d1888f00174cfeb8f745656eb4917b87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc00f6dd20c52ea6e80263bd04fe817566d22e1d855735fe5080ae593a3faa1d614b0dd7f419bdde210eb254a123d929c62a88852ce2456e6bfd76567d8881cfef741f0867714bd82e7efae560c0fee2f233afb23a62fc1baa93ead2eff8c12c76127b6e0f09c949bced91103327f7dde3b3e91dd97284be7284ef433b666464;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f6b1014f0e65752cf6042e8c32b6bd9caa0c335582b03949e08408ec51c1082423d9216b95eb9c06f44674f01679de32c3640e9ca7c25325eb4a37cfb9e1be7d51e338e8f8696afe739b84a2eece5f16083fd82188d28d02cd24c5d641d93e3d6c487a5f350a82a1176c434f05036131493bef391281b8bfbf4979d1ccd68bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7e2da4f6b0752bd4461242683cdb87a228c4244dcc7e59aee0b9f40f391a92c1455c7f8dc2afa4835d506ca299d8ef44d6ea2add9b18a0f46e4e295a276791d8184df3c4fad6418d774de247f66d67b1325fc6f81cf0c0d1a7a6584462d0db70fb0fe4e9f70ac4babffbb92daa33b6a1818fb4c93255d21564331a17b28ad2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdb58bb889ebbf5961d3d982f3cfc37190b0552194c0deae738d7f80d8dba76d211c490a51e0bfadaa2a7a97ca05b38e64033720412da7120d5e0e6b643fae25a3da4559bd4851d433d8469a005ba5e90d4d7d45c5134bdda493358ea72bf35b9fcd1c9172f6346d0cec133bac4bc10793f51e070a57b7778360fc84056b50c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f60e8d85c9fe828b628654eb446a6c300df7194d738259934fad0618913e670c333dbc4972b8f6cf75254580dd4a1288424b0e5b488b9076602b88f29029c4e99f9335da961bfed831e3b721a807ca93bc38995a7d4254b212d11447f522190cf5022b8015ff3d80ff7ef37b598e91aa072bd95147016dd1f417285ad5101d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h434a46eb03f55b93cacd623957d3ddc32c002c202125ee6934089d51ebe58cf5632148044f97606a0653915f889ee69455a0c3c6a579c070a8a61d17ea46516c202bd7d29367270b5306a47afdab5fc708a485d34ed73be7e51e2bd072304727532d06efa88f189f6cabe8d813697fe73cedf741201c39ff1ef1037e84eb16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8e96e77690aca1194feada1c22a6804ed6394f2f94425a315d58f0530ac25639a3e464f4d2d44f8fdcf381f9bc84d688e27e74ec630be8f2f3063dc648919e6d290b50ee215d14157222a6902329e76e9ec3419458266bd56c6254649e2f45a6b9924c60deac7d9073c4c4d2b8162661f289ae476859b44486d625448f0f7e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fc1b4c6403cf0b9db6649a5aa2c70314f07db72ffa457c5f43247a84c2ab13da7b41a2585e9ca6a289055ba35ea060ce8ec94b1a699b8d15c8a842ad16a5ed590a56d615b1da0ce0d36af5f284d1b1edd4b4bd0a01142f38aec95958ab8e6fa91a59e59a770771b0cbcdf3c5e2135a631b02dda71e8fb8aae915ab1355d873d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b4aa373e4ec73adb6be8f4d41604033a3ae8c091f413c1402a31328b0d18f0e1966a414d9e6c5ce9238e6f434a28ab3ec9646b177267b322cf58ef7065a98e5007b7cfe2016ce5d5fa3c010ed1095c5d52f34e9fc35cb9b38c30be5cf9f7b6b7988ff1cf553eb1070d170684f7220373affcb9272f9f16b2e440964eaaffd08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57519cfcd0994dc3984cfa917cbee9ed7b80681066e78bd69709857fe82365ca14b361919fca07805532b15683842c94dbf19810e9613761533732e48f24f61659f0d1bf1cb179f62dc4a5585c01513f7bf55c0c1b67981d58d64e1c72223a310452f575980cd5ffc1684bef20cc01913cc9c60979d1cfb5861e013fc2918e82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2546ff5e07692dd265ea348dc09b43560eb1d18239b9695d851bc853e21d7a1c489a5e0bb64f07c2c0e79fe01cbc82b97621338cd2de4553e3009fcad426e040fc9cf239cd0830b81c5ce830bb4dea5da9d62c728c4bbd80780c713d0a841f0d9bddee8a836b72945ccc55c8d14ff665438888cdb3aaa89acde487c7e67c0c69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e6a6b81b5bc486caa249ea7859eaa32c3f54ff6d609dbaaca8aa627159d8089925150fad49eeaf45f11a442bad6293a68d8e7f15312f2dfe5a0c2fa155dfef86510c9c5ad2433dddff7876891c518a9893581e4eb735936f39de5d7c2c1d4d0652f36d68c209de26ca39e1845499af246e7d06c03c6c43e71b8499b47ad5b35;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd79e23f2a165738c80e2d0a1b5f0087019b9b7d239b1578d6f9cbc864ee5c646b2b86e947a490b3e80f3a780362a9536a24937bdae7af8923e5994c5250d2c07723a85801717eda7708ae535d312f8e24e86a65a48eca6bc5c36bbf1c9dbd09b152a0284e6345f63f183a96cd20ca0f943c10245fce5dbc50980ea3394c8fd4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76676109af6c9d37db694a89cd19579912dc76328055c4804528f74f48df09ff9adab8c0f0b091d3f56891cd189024682b38177629e7b29ec9b267a934951f834745a5b2d30567fde7a9229dca2de844ac54a0df731340a1ee11c226cfe1c624d61ac9dd5da9905ecbef70ff3d59eca8f6451cdd1e4472f1ac3c173cfec08f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b1a56427e5115725326d4056fbe00b025e2fe054796ee297bf39604d884509c14214e0cd0d4a5abf950464d27b3fc3c718767f64079bfaa906f5a9be982642b3ccefba15ffa6b5b27076ef52c28af24779b17d46abbd8485098cf0307c8697f55c0963bb0d415e13a9c95e0687beb80591b344e5adbb2c0c65d271fca3fd0fd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha73d4f71b83f00d4b2f4aa2eb9b38ab03760c1cc11ea440582080f230477be69ed13009079954d8ade51e9291e522aa2663e78dd5d3fde763f6a681c9d3e6450354b062d3f7498c812dc4662f6bda0268979e5aecfa2d72b86f0e72708a31fbeac0ff8d75f6b02f7a27ae7e4560a5e79b547f37deb9c68a2f782ceed01e4342e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1860b702b6268b96f6d992632a59eac8c3bdbfde382c1810a20001d5be2ceed6ca3bc10adab11582b893a699c60c08008241d0511f61d8a167167244413263cdabc49d6f2f2f97751488b52e4da27bd24806bd971074d7038a08ae218cba458081c43953bfd3205bf52642ac685dc236d88bdc8e4d7a5895c14a682be05cb6b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cb5052ad161f516d4594d145f1401d0340981e90a280b2c6ca6104fdcd03b79c29ced5dad569af8981fecd059a3e99b0842986a00826cf632dd5eb18355bfbe111c66b08c18222475a375bc540d85e6e018b9e5af4e5606e522f608bbee328a9dc66a6bbd1396a50cd03a7b616fd2bf863fde37dea41ff2a93cf08ed77b3e8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6abe88733948828582fcde81f5336c564fec4bd2cf0498f5dbfc54422b677b5ddac9ae61c6439b899a6b3496d45a30c4d9e8bc926b89035f7805aec21a2a4be7438f2949ce91abe7eaaaad8d7dc714b120e4224a11ef2e56631c134d14694d0c6f53f2405dd68d0ce323a2989c4a37a0e60d94ecc36df16c2a82ca4560a07b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f6bec65b56e2572506fbb1665a5b900a74d2ac2320959b0c0b87a6941556c20f8f84f2ae444e33e50ddb167ee441d7f08449b2bac057401fdaff090da48d2715ec397ff89c1f8ea498414c66a809790ef6a5f056a7768e670d75261e458456ba11a79f518a29a424840dfdb4187ce49bd7680e0816cafe4740f045a4b6a783f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb75db3d9b3516c3e7e288a63f224e6368bec68b24d52627d298994c5d6bb63c3d425f379f353823f0e5743d364b13b8a5a11e3aed945c05d06cb07f44156421fc22775ed807cf58a88f4db6f40212fa5cad087a3e51a36a6d5c505150be8f6126995f82bdf3bc09eeb2ccc1604d4084ae95f016d133bc5f38418fe8af224e188;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd08b20e5fb2e750ac5faa8b889a7153502920633cde727b56449dda832e40a594a9921f5dc2c0706a1d01f9b434b54cb9a9e9b3b44e741c60e77b4f7343ef5f1d6a6f419ffed7c908cf7c35e47116b9fb81c1fc986a757a70f6929bb011012e885e09d83668e6ef4ad71e6ff5b8a8fd5167f65bab39cba6d32af96cadda969f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3903ec16972bd58659de7f48b89b0a55344c74ac46918c795dbe94b96b3df1a8f5cbeb95fa59a5d79cc93e653526d1e7d95339d01cfd6b8558bf5da5d04ff77f8b950a2779cc357e8925f51b4c95f8328862a4fe745c4d3f03217f44601403c47140699a57a50b68b74b7f5f71d7656f8b8a4167b165023655285dcbab846312;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8255b7985a0638684bbef212e83ab19e23cebfe2b5d72f02aa3576fb225e8497c40be863393bd85a35c8f194b0255c8a621a92a81c8990a8dd8363a78e516d250c01a4937263549623253db223bcc07cdea1b79345a761915ecd2c8d445bf267ee4b315ac56f042d9195d70fd6343f91726fff3fa84ae19432e7f97f4f63474d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f2174e7b2dd3aa2f9e7b4f078dee2457297401ebdabf111a111809065cad56740e2d0137604ce71043ddde932746c24f25479419bacf84cb575b26713eb4a46ebc6b1587dc4f6c53eea4ad74c2cf73b006187b098124f50364210904847e4d004b0d3dd36b7a8e656b85626eaf6579270f3e7549029853b2f39e21a104881d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b9059715b56c573c0b62f6b8818bd8ad5f17e726673d8757be220ad7225358a63b56d3880c61605f96c27ebc4da31e963aaf80155b49de71a085cde176cfd6e91b7c725b24e40df9baa9f3e499a1017189bfaeae67a6e198e2d7cf76ef29be7b660176f40fc4cf2e5ac9103b68dce03a2a31563d502d0b35294b78f4f15edeb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3991d7a6405767f43d606630aca64c98a90a4d5e7a441b18b4ac0de7d81af736f3989b25addfe0662d835f6b96699827def37588c1eebb75eb94d7965527bdb22628a4859b4c64c560f699b465e058dacc78a849ad04b275f4e7c9191bb9c0c4c9311e96c0122f04fe95bf297e6808bbccffed484252c222d7c091ff44f52e77;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ebec98379c8be7bb665faf83a2f04459754c9f6c702b2d124620cd45c25e0fe6996aea98c72e61f62e56b905ce4462a551e9875a3016a9d55edfc35ca6d8f86c553eb7ce4123d769388016f88790fe58f28d292d020352081131c4c95cf9ed103d9527899ab9a40fb6547fc74c767eeed76a90ea849e7d6cf58208a3432d73c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cb505a1d7fdb9adad08225d2d954cfa58136d237f5d9ccdce09ec104304c16277e2072120d15f0caa9667161ddeefd454e17f43aa4a4c70c62ad95fdb5ae323c89cf34a9f61f0e8da3cab76225d066f395f632826fd595a88c57d4159e89589abe947e82cc6ff64a860d2063d20b9fc04bb189c37d7a57898bb5429ae1eaa5e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f4074989cb5c101d8c0674cc495ab68c8dbdeb000a785bf7faa4bd1eb2b58b6ec66fbf2200b74508395b37c8b9efd7b437bf28c18a76f6df8ba412a26a46b1d42763da8c2455eaae9cae0dab65f03a68024853641fcd239bade13efa9fc903d01f8f2ae467a433b8e25c4f836ee19d4ec310f7dc681bc1a261039b30120bb26;
        #1
        $finish();
    end
endmodule
