module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [17:0] src19;
    reg [16:0] src20;
    reg [15:0] src21;
    reg [14:0] src22;
    reg [13:0] src23;
    reg [12:0] src24;
    reg [11:0] src25;
    reg [10:0] src26;
    reg [9:0] src27;
    reg [8:0] src28;
    reg [7:0] src29;
    reg [6:0] src30;
    reg [5:0] src31;
    reg [4:0] src32;
    reg [3:0] src33;
    reg [2:0] src34;
    reg [1:0] src35;
    reg [0:0] src36;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [37:0] srcsum;
    wire [37:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3])<<33) + ((src34[0] + src34[1] + src34[2])<<34) + ((src35[0] + src35[1])<<35) + ((src36[0])<<36);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haaee5b7bda11023e0956b6e27d43a7d59fd62c76f6b3e09f4cdcd32bccb83cacfa7809874b99526f262a1cdc03;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15393b55968ab31db67884d33d4a185be7c50fbc5ce281333ec8cd6caa7052132edb895ea0b36cd8f099ac0b4f9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h713b4a91d0830e846ac69ab8dad018bbd1d2bbeeefea65441204396136b1f5c93a9d7876b2499130847de15478;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc26a1e1c96df7cd0990f495b94e3d467fe50af35ab1c4052ef282710a9dcab98fcf3472cb8e0556d42d0b593da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f167459b5f1bee1ceaf8d9122f50726b069d201a0a5225c25d9f18d160c1263f3ae8f827321886d76d5ed307c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168613933152432b4a7f77f417ffbeb314fb6eb7deebee460c00a1c32fc89cc174adac7b7b51ad9466985fbdcf9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb7edbffa76714eca2457dcaedcd2eda019ca4610a4f1c34982450413776dc42bf99ce034e56fff338f5707ea8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a19ce528a8a80639a5ea29438ae940fa32cfcc8dc11139cc8457414768bbd59d1d393d8c0dc7412d4752597ea5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h713c01608f172027646d2cdc0e8804e285344865320c21e82ba64f4af108ebf1392c0674cbb888f3cc0678a4ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149ab2d9b82100ec5818ff0eb0d7ab4d33b881c5f1202699867ff98b6959223661e9b9c54429a3eceef94b835a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1481b5144fc896625814579f7c5aa6c483c4c0978ea9b3e29785090fa6a9eb01eebd8e0a1537eb5cc37671ba7ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha69372e2b0fbbdbe2a0d72864cb2e0c2563eeb32c22f69d278ed12b1351232ea8da371d3455a2835358117e34e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b9e8627c22f59048815e7150cdafe5ee9c63e323cfe6cbd0293acc77b462792f4e9c8fe8331bc086c0aabe233;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76fb1f282b52b46280e14a425120b77a10b81bd74592da1cf6213c182360d8fa7bcdc18923d333a3b6c0476632;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10214bc2d901ea6fd3145b5b79a640d185304e4f2446ee8146966e46fb71b124e311002b10cfe623e16399c6c7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d32bf8f9cb3f6628f64b14ad80d71eb68f9000566d838628e1042a3a172931c15c824dac3a82843323a068f0f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h83a93ebf8f153d26d5a94a65892439e74a79993f250c3f7c6c777fe838f30bca114e4017bb4b726534b07400a6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f6241babc3f09f75f0750d8c42583bbfa98b19b968310879a4dba24d39fef2369731f79f954381dc48bd5355f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a794043b7835ad393d169614024c65865cc4809bede667ea0d636c84a2cb395375ac43313f8462fda3fdb56037;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5446c8e9cb2f28dcb7db4fcc11381e0802edf31ec08a18c83b57cda87f70d587111d25e87cadebeba256408e64;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67b037fb7b90c439748bbfffbdb7d98c5717deb2f21f94d9f4cc9a64d8328a53e44838b0d85eca5781ba6b5654;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cdce0f7e117fc4092b7fdef9c8e430f8b34dcb7cbc03567808302d2350adf6e50162ef9f6a51ac46c5eeedf0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc5a7f2dc98a43c0b76435a7b679ca16fd65d949b5f947de3dd785b12145ccd488804b5003f5799c92f6e63e2b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121d727c8c8b40ecb7e4dbec9d5e04d9982e26f629c35454c4045fc63ec8bc21be42793b96b7b01a3d718ec93fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187cd40dcc888eb84b9632f352447a81d641757f9c7a66643d116428f3966381b9ef1e4ce870dac8af38788366f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3307412bfedef8bb8c6ef90fd857cc8af0e6a516ffcdf7d53bf670d699494a09ff4f08901039b9b752644f0c12;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dfb8af3221d847b8d6f43023b19eb4bfe5ec1974e606388beefed9572188a31d1a37f27ceaf8789a12761a47ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48903047b10ec7a2c3be503a417176aacb39e8cf2dde5e77e858cd90baaefcd86922d5fa6a514b8934f572d9a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c206632b3146e597bc919dd4085341d3209cb88027dbd2739153b56b8d983590801dc57df09a451cd49192050;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1993c42b3b6560a0c96fb642af8c0cd89e8624cd40cc2847d7e46fb75b62808463ac82fdff33f70b422436db0e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13051a4f69fab213e592b8099b75f928197e1b1e51b175161b0bd79cbf52cf7205014ab0649a454aab62b2bc02a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54592c9db52cd0aecc9f24730475a59f2995611479afbd303fb5f98f58086538d3d4c4e78be4d9a6cc2f92e556;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h59c903662217bb0830ebe8e6e49536b72ae29ff340280d54e080cfe92bb5e652d02a3b41f1cf823fa66bf5bf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189bc0892b3f7b31576b2b492c7f27ecba60021469ddef3ee533939910bd70d8933638956e74657c3799c610ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b3941865ee766696b6a11479af13a591f13579db68d7e18d72de9fb7b2262246c3648c2953f5690015137f8e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d731ace967990d0a2a0e2fe3c0f09b72a45cb0e9fbf85d607b8a9859d197c260513f272b4f8aeb7715655fe46;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80d53809264b8e5be418331493fe7f4e4ac22c8fa5dc7d2977226c23cb4db6f8613b6a7b62794d50493a604ae9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16d15ae832ee6174f847afeccc9a6a647e9cdb32cf532f0af77c7a37b5c6d591d471a8f4bfdd035de9fda91c0fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd6ed5273464653284c327fd126a7a3cc9aac9b21da5e196814fc521b4049c9e1bdeb1cdef9f40cd74d2d9096b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3de467e7d6ca7d7eb68186a5630d2ca2004d22c1cd213376fc03f2168e3f2c70d3e4fab05cb73798f073ac0b7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138e1e1e19cf3813c86b001c2aad2840ca8cf33aba1d0740c2113e26c6ed6555dbe640cd182432d79000a4010d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a4b66a1eb4fc8e58e12b30180fa861f1cda3ede58e99cb4e967a77296168fb99ba322abd3e67c75b1936c1638;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a57007a72a031d45969aea45e0c137494c1d8503afdcaae69a06aba8d7dab96737ccf7ff4f6deb4876164a8017;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13db4befbecd8503237632bce3ef2e19dd8ab84f807a9fe13a9d9930cea5e316abbf4b274dd9c004e0fb3f4e9ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f3f564e4c74ad3f32fd19f47c2a98580440a37c77d10780a3110b1376f9fc8e4d1e5cb4f60153243a1202837c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb005bf5871dd18c4a8fdf5a13cfdce6a0dba2a55d0be359ff6f91efa9e6fc373072180beb2b19cba38344c3f3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b58eba3eb26fe13b5dad9d942f4b316207f26036fa48c0a2510bde4e135eab8792f51181b1adf5ab8c581b873;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1855f42ac15aad94d116f1b6b70024a2ea14a82449af75c919cf9a3c291db10b0bfdd33f4114230f55eef47e7f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47fc12da81f60979ec7501f4cd2625804c458f695027ceb1f154bf4180fcee98c557cf1b09551be3b230bc5b88;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c7ec67a0ed4384c375771eaf2c2ed52d1a0a09cc38707d32fcfffc8d7270b04251944b85bdb0744f1767711ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ce0431159ec530ba560d1b5900dc68cde4932c620f3fb5a229901581e15cd30b1ea35a880e5ddda536e05be661;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde4a912f64cd1a93ec007e87c16fa5a393da93224f55925284a2d6ca4ea5188adf49360ea4f067800938f694e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18528e8045a4632dc229bf15defbe3075fc3eac6db8d13827e623edfa3fa81a7027be37ae23e06dcd0a1bd07372;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcfdd7c9f6446ae8c823eaa2c1d76c5fce42782b0709785d081f362eb7dc8f1a9386731e1b645492a886c50496b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2b715ae67c233dfe88e46950f9df7e725bd2c109db653248e2a0ddbc7555431b5ce84697cf202313cf649eeabc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163725f93ecebff49ffccddaeb5cd2156c6fb394248cd865a471827ebc6caeebceff89c84ca025650aff046cefb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dffce7c34b93553bcefaf9d9ed6b7473065c2a9ae889621d2106d92abd591a681128d8cc1d0f7c313226fa6f9f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbbd9ef1e131c5cc29ee10a8135ea5fe22c18cda94595a04950e3a8bf7b119201366dc5371004cf57c1bbf0fc74;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bb0081267d3ce7ca79979058cf9b0f699c492f4d3b608c7be43059b65b47cbd73d1ef272769de510462084558;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h558770cad82fd606fbaf41f954ef3c4522bf016ea921749ed4b972cb5d7b156a6c512823dfdedbf4b696a682d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175b5f3fe9f1f10b98d52e98677e7a907301cca079adea1906b176735a236a4e88d2deeaad51e74a1258c99539d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f27132d6d77857029a378d2575f2b3167c1e7590eab270e9b4143eec62f3c0bfcf1e94ed974d5f7a28c349780b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h975b6cb625b01126a530bb0dc41608046571e5750183fbfae1e3276bcfe51089acf07c584e64a86bacc239fe62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12feebe9ff6bc62170ac1c31bd50774902ff4349b2b8eec5d255cf6e848ae2edddcbe677664f602aa581dfdf18a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h797db2c524e693fbf1d441edab21ca5ab7ec8caf87a061e5a3ccd29b729cd7beadec9c4d879068cc19408e6dd0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7fff824a99fdea6ada2d6614d96ae7db381777ebb94647e4df2eb86b05f5d718efb7f916c58262e4f645aee9f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69dcea172ae4b23710380da39c0b2140d39b195a6b401caed2a4d0838885d1522dc92beb9388657021fa4d72e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf57b1923d1cff9aab081d226299764a7f9c4ee0ba72c7ad02cf4a70379e17b3ba012c433951be833c04b8a8858;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h74dc4d1fc55760742ea17ae79e3a3802ef3aa0c8264b6050ed06d0790193bcefc45969d88755c2e337160c864f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf74f279812a9d19e25cb3f2d4b02b78df80272cbd702013f3505fe6c8265443a857a9f7e58b0bf5cff5ce801b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4656479374fd4365e8db33ff257bcbd390767c86942447cd2dd1fb2a7453b0058eb065ae2f72c7d022d1b2e2e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16999f81f06bd31f0b4461a0345464c390536bbc1a512202714467bd3222ac449037e793a92d71fc1cb4049d28d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha507cbe7e57d72994d49cad1a2489bd17a960717b267da88ba8bf3ccf09caf19ced7ac7746aaab7460c68941c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d4c50937075d3eec69e596219706a5ea50ccd2960bf8bffd05401560770b76903c7bdc4dd5e52338c235eeba5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23f8f3b245e52b43faf362513f63022aef1f96a1849092ab8e5220b17547a4f930f22d864658ff8dc1a68c589a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb14d754de17e2436f7190516e601b77b1d7802276fcc6c28683bb5c3e712b5ca1dfd8b29d42f543f5243ed555;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7592455251513323aa52ba7a0fbb5bed1600a9e83a022d0685ae53dd3c0227b05e143bcb754e34a14e8ed84b39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5f6549da4abd22af82b1ac63336c78fabbb793010c755bbe3d4d08e4d55dcb18b6fa24e932f2419735c4b7718;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h966f0c7fd32e09e3535bbb609fe3988a07caa5f9c5828b246a86c04dd6c6ac5dcf2a6849d2a5b73a24cbaf0fac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98610c2f44a652143aeeea6424c97498a70c0ef7478ee2d2fffe2d4fff0d375e7f04af964db45204f0a9bcb674;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hea68a0b307c48dde3b1b65e75b50b9faef80d93b27413dd04d0a0a34bce5b41cfbb9b09451acf47ed4353da991;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15eb06d0252dc6b6c55b0843de2c0b3063ceee729b6776667511589c2f7c640ca17deccbff024ae42318d1478bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hccc3bf7f33c46b2873ed7b8f9adf2894186855d50dc589863d6c9c7975b6df0510f8b2db7fa0c8d1d6e7e79ca8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e2187fd1b22dbbc5013fbb04bdff0ba317a50af5416d2225a97ae6b94641848c1450dd679d10c9ffba9107a95;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7cc32063cf02394b24c21a50de54ac1cc56e875f29baa1e1ac8abab0c6c0f589f0b2c922cf3b62eff7638fbb75;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h393ff7b8afc2b07b75ae3e38fb4d3f1184ded803cafd93bec540565766d94b36e0f39c7489b8630fca300af08;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h179ae758ec25c02f5b15c642217ee75004df900049aa2409be84b6c66eda7e3baf15fcf9cfd86abfddeea121f15;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1412a0902a0bd16e617e2a19fda9de48aa0fe195990d1d03b3bc74c9851f7c29467dc24478b3583433a440cedb7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15692669bc49c10aa3b3e8d982868178ba78d86c6cdcc402ec96b3e6a85c57a6bf1524b3f989d492ff5972333a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h551cefd318f3325ca0bc5b444d17df458a24fc6098f3b90dd9dc4d4e49da4596c357c2468e89c2f9f2511ebc3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3fa5934d854017a7b83be5d6c735646908e7b55e064d7d90dc6349bb730e112b2034046dfb6a8955d7212b98e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189b7588d2eca83376b8a12f07576c39b3c0045f7064b9b1fb673b39e5a352d60e40bec9566c5b887492edb789;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h192502d39f6cd23e351455f1d3f22cec9b193ec60593517d067c918c0aaedeeb44f9826df840f9a8fae7f4decaf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf316b5d29e547af13fa8c962300263ebb3ac895fb5b5a8b73464277a807bc6dfeeff61b17f041ce615409449a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1892880648ac6584ba26dccc9eace75a508f8747692cc6b2d23c5b64faad8333ff9f6b60658962e508ceb33c91;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3bfeeaf6e007f8b440e58fb41d71178bbc5454df49e02ed50f68bde705eb08267965dd41c81190bd2a9a8cfb83;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb388f680f2c67da01c6868ce95e06fbe80368bf17748636c0b237cf68b3bbbd13b3c431155283a9350917735c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14089dd22b09d610305b08908634400d09fe4a2b9fb2e0aaaac81c70275d3f95b01aa1f4f7a4aae749e59bfa21c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161d157bc3f4d857f5a0fc7f92a0919f01cc53895a6a5fc67dec5f868829e9c584b11400d3fe18251c84f3db3e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cce4cc7f77484c4be2cd8122c067ebe3e09fb33284c744875e23ee51f7f5576415736e862353b8d5ea768001df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e45a3f67d13061f1a8951d1eeca054bb7daf94c4ed2d48be3c2e5235812bf1972b1cba7f71967647a7441ff7c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h198144a115274325a06de2211f3e7b72a50461d0b95e85f524c9acebff0bc3430bb1ea93057318d941f6600b5e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a0d44c66f46560baef1192cd9039cec6f309f3f36a35f3a088f56725455bd056546337f556cba744b7630a87e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb83c35b31b019c7bfee673fa81357160ebb2ac7a0899bdfab94884d6c28ea1fb06d9c46de7f29642b97a7234;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111a2de2bc55d15d1a8f66d301a54a4fe65be32348d8aaa73862208cc4439660af6f81e45bea444e933444f42ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf01703ecec887dd53f2041e607ccb647cb13f042c82940954e3c68a79895137dd84be7759ae3ac09a98fb7166;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5051dcbc2f5af99786986a845e1e4452d4b01b2a9ac8834c92ddf40082acb2d565f5862d64e1481dd0003324b2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186d9acd8dc94a80dbaa6e45e8cc0a0b58550e67ae3514259fb6e8e191473a6cb891df80e89c88dcdfaa81d1b5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1daea1b127e9681490e86a4a682f03a924407f2554a8f0c3b9aa9f1b0400dfc8d9ef53bc02dee8255f135a838e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1223ad0372e7ad2530ffa763907786c174f0c5260e706cee707b5fa15394e3189a6c1d2f14a3adf0ad602d369a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e29e240feeddc1c584f44c443afeeece5faa1d1084023c3c5ec768d025042b3d8822a4a3ab50cccaf20ec7378;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54ea6fc049cb5f084e6c292a6e9e1fbc1d3cd096a4224af51c29514227ee1942a221f33ce111d4bfa9e375da2b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28da22a11f3115cebf9ec1c1e04242cdb1c0604a872709e755f3251878a9320e3fae94218f3ad42c732c84f39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d464a261f5ec4d8a9f818f2c46e46394c41c835065fa184325f3f0d7689e7bc1c39abd0aa5a22834e529b97f2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2be1d56df5fae9cd1437d43a9d5ab79c6c6b05dca3ea42664efa020a39cbebe5e26944d1f3a3b41fbadc909cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cc6d1f04835db8fe428e1f9880191ab3a366fa2718c41fe6584c219a7c8780eadceeb86b2395abbc8557102d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdbe02ed6f5c55af737338e86116b014f972088da13e058a7e6ebc10126b58762fb0f1c102b7e446e360c7758e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19e23c00ab2ff0f2dc868d8adb7d5a24889365348cd25122093e7e37062be9734adcf1fb8619b2f146a5c170a3d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd68c86fef7456e5704c0434fbe618c8e39970f5c226d552745167f696c8580dff2c963c7c24f2ee4a56ee1f970;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5cc4123bc32d5302e3907b5efaddc97e9e3e639170e947298c32f508c284417a0bd54c78ad224368312ae3d6b7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d2b61a47d34a8346df7f5421760c041373a270e3d7a5b08e1a666383e043fd2af43e68ceb62895b3082326a5c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19cce63caa732f9b753ad150bd8427b710351c1155fed406b1e0c0a7a95d98dd82792e7167b2f7ad16d41df22ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c16ae296764a46061e0d0c3d006388d8da927388f401211f982249c6855208aeb69f5d259df9eeff600c3ac0f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132e0a840f55ba2959b1e03a9ae14c435f613e909cb4162ee940f474891005aade45f01d1ead07e8f52665dee5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1630dc822228d1cabbfd4a2b2e9de7ef527e46aca484b64d89ee3ff7474fb1487e0cb71ab3ebec50ca2c3242a97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb61d9dd8a7df5814e03b6fb6feb125c2baca09e0924e9b7e82dd0ad775bcc603e088f67f2e82ada8565de7780;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff3c2baefa542a959eb152705421b97bd7e0ac83475120b51814386d2ee8e6887eeedaaf404a190d12443a842e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154c718d771fa5f4a10452a4bc96220dfc52d8609a5c27367020abd6e50e833440706b4f1214c720167e9faf42;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf5b5fe5f521c027b041f4ef8af84bcae18025f5a1a6675a77a5577ad4de9dd31993efd329e86bdecb0e94806b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a00d4a54487f01073933d7eb13956bf84a83410a32bcb8b942f3fbf22a1c12d1b2826bca51580b3951bcdf1f48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dc5991e617cbfaffd5b0ce5d3d388a431710dcbd486d8402f82a6c76e868e9ba88d6fa4ced75665041b4511bc2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16cb11f229ec248fee915f128efbed393f62ec44629a1bc93590800be99cf4e837f4bd4ddf98749dea4c3389c4a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c39ae2632ff6fb4d36e46c2767b74d4c3ab89e57089e992c67f59096956deee5e3e1d3e022c5e9a9dcd15df865;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d6931fd8264fff522c327f7b9c2f276865d6c20aa26c4b09b53589b54b322c3e1c2c5a5d155cb902ac03541a3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h174f3c51d2a5106f9f7d54ada98f5912d9a141a58a5f7b7763ff8dfb800541bad72e7a44007064b864a30f38f40;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3cc0ddad896fc22de7de865b3e9bef7d4f1242be0843cc630494bf3c3ae67c274e847f49cf7914cb3cb4000b4f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34d616ef902270793abf4be33838da70f3047d6ea6af61f9f614b3dec95f9c2e74d0400f7e172813295ad77499;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h169e7727ae95df07afc3c911473b1ce618ed6f2c568a7d07caebf515948b7f2f66ef335232b19084694c9abfd1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3382b53f487a541933e79e91d20fc43e3fa6cdc895465e2f2f418b188d05cadd9f799d1214b13b47ed5af72b91;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25acdc7876396efce55c7760a0d5adb7aa90eaeedf609b5a1549550a3bb068550085d657b7f357b0155c06df80;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb391868ff95c8f769ebb1debeee378129b286cf51c5ff0e725b316415be73784e13df8501f6de3f29aa8a769;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aec0cb791e82b6564c6fc2ff8ef0c1ac5007f73ac3e208379dc9a5ec51b5b4e4d395b9e9ed84f319a6dea7f99b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h596c4affa2c0fad50d90c6b50bf7b91ced0065a31ea0bfa3602c4ed4a3475f82e4d645952870f0c981507c02d7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff8b15101c6a519c4181b80096f8d351b5214d0c4a81e8ab1bad68c2a50d76b0f169fa5f66d902c0dd687aed50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1184291f70c79c18357e2f7385ec89e3b4c9c7af2e9e4cbb1f58220c329b714cf03a8f2a537422045e772b74c7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he33147f13a6ffa96a4f2361021b75e59a8917da7130517883cd8dd949e4a38b53c4e5ad78a65e0d080fd050b44;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ee9493647f282b37bf42430c3aabf2135a0ccb1125267b53c1f14ba510d399baef9598777668bd737c56451fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23c7d6715840c0f3459be5916678d44ac15e0372eacf63d7324c562a5ca770e087fcc43294f20066dad2a24ab8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58be4d14070cbcdbe2df2639543d13f89a897aff6229a9c934354683e46fa06355e405c56de3c4954a64c5d4e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1122fb401d5eb541eb1faef3d349309c4527abd3aaf557cd4031b35eafaf14daacbe1e31b9ed5013c32c1d8c15c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12aa70617add9f2abd688a299c97b1539ef47fceac89e0280a35f45f5b5a5c852fc557d319fe6393754c811a2fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2887ef5cf6ade26362b9472e1e7cf8fee3175c8f63eb55b1d31ac2c9380d792b370cdda0b67d35f8f41f3f9460;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc293112639cd419d770886d8e6dc8780279ad482e77a672a27baca82d602a3217ace397486f13d30fdc2a6d360;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9df27ff6c20fe2628a3949bcec19c0289c48f859d32c369aa34af16905df7fedcbfa643e9162cbb16a914ec806;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7d1e7f6d4cf9279f84a81439964769c3300015c7cf46a953d8a6ed642ee0b954ca5a2285186c2bb287e4fbce6a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfa2518a3633dfc97d85e168511e9711828f08b021ed179fdeefb22190e00596be514b26616f078ef553d834439;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbec930b2c22c1b4356c17991f0263df501ed02d4e6924e658819feaee306bb07d94df4662ad69baf22a4aa721a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a8843bda2252adf8a259f4d2526295b3e0fd93ced21d866e1fd32c86fb63fb5f25e773c4791435f9ebbe3fc0d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a2d6abe0dbc00d24fd7ce7dc995a7b00f8eb1b66bd5c93eae82ea230959f558fdc3928318042f4a5385f6c2f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a8dd382294aad09f76b1025fb1c17d6a6cc2bb32ce9d5ad2d44410125b0af2ec720788af5b75a4b473bb8b070;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc0abf025df62ba3198fb26202bdcd085fed2fbf40d02642c611d304d8d544af805db35140104d6c32443ea69b8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9cdd61989cdda47e2c0b2954d7711d4443a7ebdc7835b4a4ce54297ed3304f1dc7228e0582eb165c51868458;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e41f2f254450d325e384a7eaba4a50eab09fa0bd8ba8a0edf66b763abfd84f67d59dd9d31fcd3c66bd434b37c9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f971ac3d569a21cd6362a92d9420257f544e196629cf321bf53e5a5dd9b7d78ab1fd778c38feff6e86b910f25;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf9cc48289faaa797a7a62b6ef94d81bc0a9e0c159af501d37eada74fe0960c348d937b0400ade710bf7ee34e4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1391d24a4530c4fd6d961b92ff174c67f880aa0ee8f6fbe66b0d3a80e8ab48ab2c2ad1540ba4387d70985400d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h57584323d03c0f852ed23cdb1ff28d1f9a86df946bfe8e59f7537dd66ef93e33c86393fdbfda7835509d896bb4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ffe61d0a586227b095cd7fb4d3bfb29954200bc2b9b984ed41caeebcbfdbdc9491ff9c4eed854d573987703a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d67dfb24a838814f7295a0059bb5f8d4a27a22e37de309cc32aa8bc53d562811004fa94a02c71bef697f961dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191c153189beeee489a048daf9e3fb2720d6dc2f7486a78e0be71628ad976f5a829a4a8697f90af4631e131b163;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a22ef09a59a172d759443c140a6f08f5a97304e86a75602d3d967106a39877e0b9e6f49e087dc994cc06a095ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3510e847219fc9a849fdf099655b285e6451f5be88895e0ce263e80ada0ab6adf41286b1b398b3d2a034356356;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18502aeb39b74d5a5f56b266d4ed61b2f5d5fcca2dbbc0d93d420cce3818b08ef4d461cc1ac34486467b7231bdb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16f9db938e5d599c520bb6345a64d5498ffa231197c0e088e3af7d737fb11d2da705c6ffcb7fca6f39608ce5ae8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a745f8af3f69b3ac662d6ebcf5bc24ec0f4af9c2f2800ab7262ce31212ef7c59d09c44e395f0b0056e2e78be3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8158c6e48625af1bce414320642bd15957cec0b0122f1ba2fd56d341d96757054df827aaac2f2ce0cce46c281;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h158350c936ff6f589eb627a99e43534800d7625699eef73ab947c2d267f34d7e89c3fe1e7e9a3f545b54ccc496;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8382bb72974f9ee852aba8463d161fd71a780e32d548a62565c6a2e03df8d80d5a7d49331c8f8a9b54ebd0aeda;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10e46607256fde4465cfd1296d1d70fb67c97fb582a3992d8ce658fc8438df3a80f70e14ee66a6424dcda2b0d5a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14dc603f3164aeac419a3e2c54cc6b13f68f85f69899118e63b6edfde1f7247ed66b501bbc0df090b2ff5cc7bd9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff94ed2fa89911e926a860d74b6b2fd44f883961a61591f71b5d20f60ed73b6956fc5a1ba0f199915025147955;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ecaec6220801fb1445eab800fb835d0193bacd682f0e916d2b4763b960bdad75d567df0c13a01a9ab5552361f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164acd9ef4d2f711f270665d0f6b502b647df0acc15985560792d62b2d985f77e406193d9b49d75f1951b2651b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ee590d11a23c794187edca1130e0071fb23b35b138726755d7df894ccf9e047aa04c9b345c55191e1db78e38e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6ec25a519ad37cab952199dcf6bc95b29b26425ba378a82e2259b9a9f9e28c800bc57104bbf9e578bdbd6384f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf11c1fbbef022aafc7f7a2bf76cb751a33e7b965a21c1b6c55e55559b1d100a817daeed847d51cc22a905eebb9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h27db0aee52abfb165b49b3b4c866c37846fc003fec75ced38684a404b4b10f62022af26bde72b3ccbb67f7a585;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43da7c5fcb20d8c6f3929cc06a7bcb67aea9668f721e18da2f10a8fc5c6550bd486c0423f73861cfaefb7c222e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he524ba0d805d917960a021c72c6d132c1ea810b57ce6b7084c91bc949f6500bc62d6d2484bd3e9d8daf1a099e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1469322e7c288a7fdbe8aa9d419caa7b45dc6bab648636f6b69e7e48f317d766f04572055e7ab53fb2935afc1fe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d95247075c322edb65076d0abf3006fad30b42c37d3b05bbc999f711c97953a0270d4b301ecaab7e7f153031;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60ee3708cbc559babad54dd9e16db0203f5d27673b1ed777beb05887aa67bfee1ea45084ba30ccbd22ecb9109c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10e26a4ceb69f5efd9fa4eb836f260fa21dfc25ab2f9600e2f6371d348ae7c524832311219598c75aae94f3b6f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a0cd7a6e270451a9fdc713cebaaf0527b607c1803d6507a9878e9b55d65c3cdb55dae678c59f7066c0cfed926;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc96255787ef8f3042506f5ade4c74590b8d288298f4eeb118ebd948af1fa00cf9cbea1298f87b106473aa4b66a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d21967ff75f92ba4b255d0c19690c48051c2d31a298b4f193b0b1d0f722c50c98feea51f408ecf11e5a4daa33;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc983b079d53e31c94bb1613edf1f00116acc52f1b32c5d8129e25c03749f4cad7fbda7fcc3e89f78d13d02e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2da32f1db4303f872597c99c4f12680e4479c4e488652df0849e2f183870c92268c641c53d443db6fa22df0408;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19c7e5632f4f3d5a43393c9c926e5165ad7d872d15d918b8e97a1a9593dcd32fc132511486cf0b31370c4bec86a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8093a00b23d626a3ae27e3d8ba1f644bdc6b7e2debf5f0c84aca16f5151246f6f7ebc09436c119f9c59e879a1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1096613e85a7b17d19a419112d6ee726c64fc3a806518c27399626549babc4806653826f714f09d2e5f95f6ae6d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd8779224d7080ca755eb52e907329e255a9b8cfe6cd9032c47ecc3425f75d7110392adc6e4c80fa043a4ec3dd3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19370406eeeac8c354bb4fba2f304696494f9ec1907c4a19e31cd7c9a8088ef9386cb2ef1062750dcaa05b77972;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4bc0b9fb7732e21a33d37bd57b222836f08e559d72783b387020fa264aae07fa9905eaa17d47f0bf68e6433e14;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1094aa9cb1943f85047ca22cf5663498b11968f0648d9acc3068cce5976fa1626da8b0d205aa3f064e54981b5ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h975e0b249f25f139c2b79471f2d9419bf3d5dc47a9d576e0514b61287dc1561c6109989ab4191899d9a0a12e27;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e065350094d19b34138a0471a613d7fce3def2470bd4ba18442359f9dc3db699a7400f32dc9e87424da389e9c0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d72bc99670d8b38099ac8395076798db5fb28f9731e2d5aca1c7d91b200d643d8587be4d2cc6e4f5d6688591a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2186991f4d4ac3063b02d8a85ea400afb62799a2f2c825801786c0611c4ef1ee12eaec949b162ac4db51d7be15;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hafcce1d3dd82ceac25e5ffbff0dd6860e69c93cc84b5e4d013b01baefd6174ec18b679db98825316de2e03fde;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72a596a761a5ba158d18f0e9846df73c0168ce8e1887ee5fb7819a5c97970cdba153732d689546e2eddfa42670;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc277b12fc91eadaa19cce08ab5ba678b7536a848d253c016f0ff4de8d2782ba0f82f6e879bd5add1182fc6f187;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c9342821b34076cf46d3b4c8cc10ab7fcbbf68a9a38b907d84116d7fce18df2c10d67f57bea2921880aded842f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c0e58ee4e8f4f2bfbd6fd236d9d8c1287532d213893d02ae2917daac416801c33677c06e06f7dca6b288fece9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16993d353c21c0ee04458df75091bb83e124492261fde4381d29641c84a8404613ae15eb48c1d994686fe41a46c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dcac6b5957275a7627b3ccba3698e78e17e9a25b1406a68fb876836677009f719386e8e375fd497eee9c2023a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc6750c3f85a7eeaac8e6c147cc29ea2a33aab01c298cb5e2f7bb8b967dfd17a990cfa5bc629698cb79db34c029;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb47f06d133ee2e0a0271e6fec29714050086c05c5fc7a1ece703cbccf8e5ce0299c8125dfc6d40e5dae500f714;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e63fd056e10615cbfcf337550d32bb7f13944f4fd6a47c5938b54f819e8c2cd71091de85c214fdcad7fa69b9d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117a0a803bb23275ac1bc7242d3964fceaf17dd62dd837b4ef5639df9fe76beeb01714a2e897c334b6f7654aa16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed27dac320d29ba378403b46bd5809a85d21be004d48badd0ded25a959bf991846b536ee92ad7c72183aa8ab0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62b252ddd37b7eb6d177b90b798827c80fa40994dafdff8ad19bdeaa3759989dad956df44bb6c9b47567721a6a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9a2b2d04dc8466ebfe11142d2640230ba4788538b786d89e64794d546649e5fa225df7bc01c4ee0f6fba8436a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2b8365d16d4755f172d8a2539a875e0cc97cf2d779db22383882c6b34bda5fc8de1bf910f55d96a1139a2087e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h915a12fff750f6f167887372c1db4138866a9ef050f63f896774514904ae5914cdf241c951ef7a04afe0d0089c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18236671bf3f8016c782542837a0ffa54083902446a3b1bba622741cc0576f8efe20c204b4c4d03d7914ca8f61f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bfdbdc3d77ccb02a4233ba96343bc5decbaa767ae189204313e229544408add9c83aa7b93f8213fa3963052e49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce1581ccf999d12711e569a2be4af60f575e5a4832c25f7dde28f979aef5cac4a045096da6c40799247dc24d67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc37934558359ddf5264f1e31c68bb67f959feb07b4993d22823e273e6585be276d47b53d57eaac819d69289c4b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h97798125123bf15e17fdd24154228a0f34d0a4057ea973b87dab52b34c5831e7340c08f83c5f3850fac0d70fac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19bfe9a15118aa223b074d8ca54012afd6ed9d6b6d75eca7a1faa41b498332fd0e222348cdbd46f59540dbddc65;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hec3c512293069425df1975c2a5c9e45707af9e344f25e5646028750fca9df0514762964613fa24655e46e6ccdc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8132e117b0c8302acade5cdacbaee38aacb0239d4adb7e709ab0cc4787ce238d8c62516e5eb62d35779b7672cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5875d9da4d620ee249c798aad9b002ee60b11c178f0a6a606e7e2146d52585119db1ea16ebe4c754e01e976f60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h155bdb6a1709850cec63667d8a3ced290bf5a94351b0f1b5840f6bafae32bb7ce837da4cafef11c56b1daae49bd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h192868516f50dadbd236a4b5baf7570ad3c9ac86d83ee0ade91b35098c7a187247a6cbc8cf1792adb46e7f958c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe1b00a7e70fe7885e12918499e415cb3e5b81e63095358624db5228535e78c20f07ca1d003aed01f66a62e860;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c1326b9eaf8b39ac326f52975709fd2141ee589083847ea42d2bc90fe97e46002027f81e544c3cfefa04530fb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168118da140f28d4ab2f2f940421631876b6c197b9e8b87bba70f70a2af7621f317478e0168c0e854cb96bf1841;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1113d443d919f7420fdbca8b8e2d083d590947c6afa6fd7127d2ea9e07512f26728250103b555655a08f6071dfa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f86a945f0b80bfe21ab3dce57a7039f1b8206edd79174fdb56b0d609579952d31b22df7400f779abca3cd8494;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7fd05b74fd0399847dae9706d03ee67be8dace5b32df6b68e85b78b0eaccaefa4d2b9d657f650aaca8376ca7ff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bca567d2d99ae004ce00f9a51879fdbdf46942243c8d738b0ddd1c46fb50679f744e31c9676c605d39de5f5ec2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h52f906671e91c79dc3efe38b040aa1ffff71e7cca2090527f8da660a7934cb347d4626ab734f019560d5bfc9b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h439e17f1e4e926989828b9688e1aa85ea352b2341fd89adb3adf2f392eca6091f2e05ae4acc08e119b1deea6ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf638f8708fee6e7f0e45135c05e8c4bc0c3e24d49665aabbcbdcc2c3b7528c5ac17d7ed0d1244c0d497976a354;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3aa8cf1013e4d27fea3f83377b76f654815dd38cbb49cc593148c55349c0cbb04bb7b70becdbac015cb19c2252;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125805ca26bc4cb08d0ffb83205c83775e2d40743acc7c4911c0fafad24a1c1cda41ce5c55c43a949749c85be46;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb032533d52213828cf1e821a97d610eee17c4277180693b8e49a38b09978c6724aad4ae35437c02954848acdf9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h49fc30ae237bc62b67e3d9bfeabf1c911d1cb89c880fa57518724629f07d2eb58eb5085906f598b9f226a2ce8c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12e0a39ee1148dab92f75bfc8d688265f174a4a90f86c36544cac38e8844222218f4cba45aad96f578973e9849e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19e06f076cd5d1e584eefbd5707ede4e026719c720e42afd0a5c5f670e1cbae25cfa487c6e19f7406423d5cb36b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbdb75478c7788e10ddb862779cc38053322d79b5e256b6f87a0c7d5549f1c1a70c3df9f1827c22058b96b84a47;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9378dab4796a3a5a226f5eb84562833e799d7194d9a47edb066a3bcc41948fe86da9498d6071c683b7164a1d5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1516544a857338379a04af8273a0fb54bf0230cdb9861b31758d442ce7b0aedc99ce10e6fa3aa48646a20c10279;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36597d700f06b2ab1d73cb44ded31ba2b1abe30b96e5adb76379930c15726ae5d84225d57782a5ec76bf0d7837;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1491588bad6c4652c85f54a5594d1bea76fd5e4d2cc47eb1f9279253efe85c7333b81de08012bbcbcc61e047b6d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hadabc7161c2fb7e01f1406bf606a2a49943a7c318e73d75c3e7ed3828877d0f593a9a290f5c1e63f8807fdfcc1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d19c8ed7c7d8827a8644e12903c34a7a62513d58c341c8188e4faa4daf4767dda62d17073cb6ab3068222a9ca1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10fe27c51d13d1e3d8e7901e16f9878ae67ed403498146c6ec3d9fe9046f40f23a4fe56e4ed4afcfb0035e2ae50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b33f95985bb0c28a04109aaf57d4863c2dda5f6d852d15b3f289793216a9f5d716873ba8bd4e89ad89c859642;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12108a0e10ee2b8b19912c3888226c6212ce41923bd5f23764eb705b8f590add285730e3137c75017ef3541b6e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c615ed995d8f74e6bd8a799f73ce30cffcc97472f7b5c3cb4c55b027bcba5b8761c85577e85157f13ebe5ea9dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f5ca019aa11139ffc01e514ea2ac29eea178ff348798c3c4e27c827250da92bf5a2d411048b6d3701f70e04c6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heaf55a2cdbb3a19a03a0208daf9e82575ad30b7fc6ec6c8269da2da57dbc76bea773aa4af00acae5aef78dd7e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h879d84e5bab79dacceabc07bd772c2952ac35314d6e94494d9c5a2cc1f2d71c29945ea355ebaac6160d125864d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16431fe69ac616d23e87d80523f813d78305d560f03902053f9a8f8208d4efc3667ee251d1f25be0dd9cbc5f1d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1acd3c28cf5c082deb4ffdac07d992061d41c6881ce99e80367b0c2cc4f98dad2d5ae3b796a9fe7611d5a9c0759;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12270616cd41593d827258381bf33842f2be434f59a3ecc792c5d807d7cec5fadfbdfe152e90972519a8d09949e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ca0cee61a3c6186c04c8a2effcf2efdcd3055aba72110e8fff46e0439b4e2807e64339f482e11aa49d690e64f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f737886f28bb88aa3d13bfa3c0291dcc0799435d96365085327916d0a9dcefc39760bfd0402a9121582deff22;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163c848f6d4d4af9a15176132fb91724f51ea6fa8b5a30960275b9ea9cb5f9f8bfd75d05e7bbbbeb81c25a22fe7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1513bf723245144d57308b5073ec5f63c1cdab226f246c9c080e713fbe94d0d683076aff082b48f18aa95732a21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ccc31040a53fb78b705e25b78d1d90ef074466087d9329f3e9a6d0e5e72cccb13003a76d2f5b7626ce9a71979b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15eca36b00cbd1864ea889d923612e1dee3f8284da765e98f6e72382e796b21f4510b944ccac4b9cd78b91fa8c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d4b72928cef121558b762991cfdf8d81cdb05b0efe5fae16592068b843f5cc757d81ff64f35333c6924e914f7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd805cceba14a92d0eab0b1105b1b2c24604987e98ca8e8a93cab75d304a699bf620915ba9d8fcf21af6067565;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184d7d7219b6dfce55a72a927b334cca45dfbcb473ef2699983a8d748b244ce51ee5140da7792a542c99ce059e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcf521c58cf45a103a7f5fb0669e1fe4a84a1f5acd6eedbc3fd10ede1360e2634f84471b40a5078f8ac48ccdd81;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c9f6c42144073a46d7d7f4a82c16b769b9a4ab9ce2266657f56160f6ad79cab519dc75a4b8d69a6fcbeeed053f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h90690882e027453d1fa9c0f967cba85dfe77ab9eb4323f744b2c4714b6d71bdfa9010bd8d2c71a8dd7726cba2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181c3c118ed0c215cdf5b2a0b0cfad56b362716d53093593bddefd215f20d70e2f68d632997f6d5335d2dd3114c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141121bb113cf3d97da40bf109df842219eaf7f5bdb25b5cfdd6099b3d2a13c46c0dbcb4ac39b927ed2a7c0b5dc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf61eb20f95b4cb6f89862d9b9189fc52d194efc4d8ad1ed9f028564202072f50030e70f5731587611cfa0fa88d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec5a8267509db211d48abd14de0fca0faf4b1370f0efcba46d13e35e66bc3b33c51cc2032b83c1653999fa6b4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11784d353e991ed4e0fabd360f67c284131b4429a3c083f8f5d59b40bd6fe695397948a2475bd0647a04bf10f99;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8161e20062ec15c5956205946eece72cfc9497dcedc0779f763df2b5269326f44cb025c9569af3651bccdf54dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b92835c481ba5127e7d3cef5764ab0dc9851224fdbceed9233ee3d47de9c2a7c16bd16a801ddffecc8846d5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116c5d7925b62ac829eafe8d78db2af126efae38342ee3b13bdf3c923bc9c9a9ae0e8130e57c01a95d221c11efa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23926a670cc3d8f0d36eeb802afd9f695e98b37f3c9254dc01618c964ab29c863b572a56dd72b8e1a48e6d1b4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h222f9009af3162d6a5df02f616b961563377f58a56ff72415f27786671e40da75938d5c376c569ea8b53c4f7cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3d8608141a6578fd1f2ccd52bf934b4b5cc536d0615038dab7706977c317057b0b14f83336b4aba34c67d0620;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h145fb7df4aa344e186957278589a8b6271576382669acde4a6838558dcc68460076e5f59117a630a59e75a64119;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150bb0f6935720109b836b5dc67d0dd9c55116300d44ae75fdece14f16855d51a0a0f84548f8d11240ee2a22e79;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c98feba291be93b33a81782f124d0403a5c43ee61c23d1ab4a67bd75dff8b5a91fc250f4593e92beec15fccb0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8240aefe7ef259b7b4771ad64e2d5d940ce87e53236bae5a71f97b4c5d4100294964943681eeb73ec03489fbed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6073148ecbe099849b71fa350802351cc83e3d563427812b7fbd068c8396612b13cb902a56635ec33e6942a20b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d763eaf179704de01f287d7417e7196fd224709de162dfee4c00426116012a8639da497793f4abfef7691c746;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3104d57999158bbb63971603e02d384bd47187a29894406d35bc1944c7fbe418eed6b24125b7b290aae027ad62;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ab40fc85de45872947082037390f0cf4c3cfea2e74815613d2cb70889e5f9351b1af3f5793d1204f7a8505e7d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132ad678a6668bc90e3c6211b52c66bd56a849d6d73bbbe98e241ce5fa77eedebb5f2954afd066e86d6b83c82ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7b8c27755ad02dc2bd41c1b0b268238b36bec76b07227ea8e41f228f27fc5b16d812929b3aef032be2dbab485;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h762042d90f7f53f460049257cd09c6f24c76318e7b57d4e27ff54a93c8f6021265e4eedd24116c5ff2efe484b8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3746778edcf35fc8bb123ec43e0cc89ec859df22d9f18cacd7a90156cecbc6af1f65af4cd0d1977a61b7811d09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a73d5871ffb28c60dce3aa5a01c92a39b0284ee6cce735ec21f81a0b954bb2dfe44e5b8bd7f26e7cd7bda6baa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14967bc312df291d991f2085e67903c1a6a1b7f54309a8e5d050ae6da2931faa3e95ca9d2f38eed28f3adec7007;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h837a56d8e69312a431389ab440ad3138327a608eae5f3709e761fab05966ad9831049e1b07c789e323d3c5f58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf48c5ae41826623264b634c708f2f788ca3d0d296c321d56936aba53ada87c8e56e095ee596251bf6a519d542;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4064a2927089fa8133a38d5a36d0b6a182ec13a4345b8edb368755c2a4b33567cdbf946c74150097172f631c92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf4bcef5e24958bbe492b0752892ff049ba52ec2506954dae556e0d989cbd1348db0e7b135267d2de10779bbc9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h96d16b0c52145b624452747e285103d3bb5d2b722e887ffe514a9417c37fab4305b4038ce3423ccc094c672a2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f1a880ecd34c80133625ab9d42d8a00f26b320b8af28beb16f7be0e872f89781418a94d0316b03d1341e554dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178c8bf80a981b401b4321dec78e48a52efe86490c16b22c01bc5a124ce914a5c17db18f532c6c9c3d9d130bed0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db44a14077d78a2640d260b277bf76686762fd2042fe886173b2e2202527770f1c03dcf841a62d065881fef6ac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e9c39675338cda6f25b0157f0eedc2e1eb2f0ef2ca0929a2738704b3699a90895b74ed02ddfd2dbc544bca805;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3a19ff69704c0ee0c9bfbfe7f56957c9ca7d94873cd6b30b3e31cd7cf193669408b04ed4d633d8830fee2c6a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3335ee48eccf1af10d8c84ec33381d5aab101521d6274d91bce5bd376b91d403af850725082dee4d66333d9727;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h190ee985e2463c8a72430a96e0faf1fcfa11fe4c5d23400cf01a3c699c62e753fdbe87d8234dc0ea2a4e7a78c04;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad38b9c99efde26fa9ae3b529218c7b4fc170326db30020ceccdd7c99953edd64b7ba5e0edabe4069805a224a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f43109ee32850a9b943163dedcc4a9c5ed64cb2ecc20928eec04a57186b74316ceecabcecb7fc19945a09f3402;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb71e59640bbc3185ee39c3b97398808203cb630e2a9def6664901ae7561a9f46aa5456dea9a7f7f643483136f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a082f57f70b60e6ceae2e9e3deefb031c4e2580a20ebb6a16a81b41661d1f3cd8d94d9efdefb91621f98f9eab7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91fa764493eb7c86603eaeb4924c80c02eefeef6a233db100b7e0ed44234d2957d723e0167de22d484cca9223b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1927f8e1d84b4593e235bc488428b6fa1f0ec3912907d555e367124931c069794f929e5707c0fad858f45781032;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h232044d6489e97f2588f65eb9be3294e142c7748717cc38e07e31f22aa55e0c6f643a193aca9f0f2c0161587be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18286cbdaa53a837855a940c88c803a757f28080a820e2b9368b51eaad9421af086d351ef63c8f2a1b8e52ddcea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2bb2b4987df6d022cd05e43a94244a8f9b98cf8268cb993cceeba83f6fadf8ecc32f140edea530fbc645c24984;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1067c28ce12450c7f0a3d4f75595113d00ff93af5245346568ae336be216c7ce85fbca0261cfbb2e551ca10ef8c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f33cd36e80e8d3a2ed6a261660a488e71a3b6c81dd06d1efa318b1e21d1563b8402858c9afa9cff4f0b77a85f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h44df31083044c5fe0ebdb3d8297a92ff148ee78220259eaaa2313091c1c849e4390176a0b85239b6a0044de232;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9befe02f9b1379980899cfadecfc8178ada47ec4a6ae550ff66e914d36801d1c3f505ae339dd2bf7b513d1d259;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h105caef25fb932f9c1c72710730af7268ecf6380ef44a5503e8229823508d3868fc524f2c7a54f58ae8a1daf585;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7c8f3b6a407d01d7ff2301a853b65507fcfe3c0441110c9624d449ac2b65d7fc77e88bf0164fa03d795e328eb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15eea198cd0ed3a3fb261b22af140899e2ece4c3616f0ec72e1982778dca66c9515a74f3397eda67551dc2de538;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148f2b4a28ea4a316da4dc74562bbbb601818a8504cc338669ff1e44a7853981e80110dd48a2fafb5d4b0981600;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c54f44601b9bcdb988ffa573bd8fc958bd94ea700e2177b4f247d92a63ddcb1586d981c9e3a4f6cf04af31072;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c91ef28ba7effbca707bdf386d00a93640e2bc95877bea8f9ee3f79ff3b69944ed5044d80c4c4bbac9ed4afc9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c24edb775aaaf9e0dea2bb1f8644a2a968898828ee1e2989bf08cc576745e66a2d6e86e5f9e91e45fa90e4175e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1620595bac0cbd9015684a5d1bc9bb26c135e63fb1c2dc2f3fd0449784c92b1c4a51c441514cea9745a933f8c66;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ca8c4a433ffea5de33b61e5e43b3975bcdbab93f497b46d7b99d2e98dc7a08ef1b4f2a52e32031b6d68f7ab2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11522a5aebf12618489814c924b7ece5260a82090863333bf8fd3406956dc6851bb511cfbc4737d511f0197da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf4ad5ea5fef6d24bd348501ee2e9f9ff5042d0d66826992dec4b8ce323d4627a9a9b427b6f5718127cd12baf1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1365b497aeae70406b284e470eb6fc86f040763e764e8a3f5deacd7a7adb23968894407688f022c9241e10a1b3e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1244d137e472b876f3e27d148c90d07b12125296888166e019b1b9411acb80da7401f053e2f1f3b5f51a31486;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f2be1ecfc41b01692bd18fb961419c983d88ef830e07b619e3e679c29d0ca5ee7acd3b76f3db8a60e6b67d2d77;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170affc876b17af88609d523cd265ce92b2e70350f37ca46d9e8e97cbab2da7da8337aec1cf38c603c04fb59644;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h120bca60696424031c230726921c125cdd933aa4c98983cdf43fe99b5da08255cd84a38765d4127251cf410f860;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b694131bfdd25c0199a34dd5e825604f97b292350446c9111ff84f303524463cb2c71ae2b15dae35dc5559d52;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h886457fc9586a79a76344c73b6eeb89b0606be688590f2289f49735f62862bdeaa9cc721596a7384ba896a4f55;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ddf25830355a2ca40e431321420988d882ea0069f5bf654d62c2feeb1736d822a6f9ec284f3657f373a4ab0e41;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdeca40b46c065414c50154fbe95b29599c1fd83af1ce46ceb3978b4fd7961de87152a0a3fe89da66a63f8669a8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91ed03d448663b4647ad954ae12c7cfc780d10d1db59697beaa587f830ab03397617112d7d53c3c6068e4b323e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f4bbcf66447d685bd62fd39a4b1e70619c16b5e0ee310341ac48ad87d210f0ee23101228e4de696e2577fb150;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda9b08623a3750a8afe9a4f97d44c86b3ebbdb73da6a66b940fe5c3b6191a3954913b9c8f6498b583105263509;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f15cc0b0e5d2500fca84e012d3e835090cef42e31bf90a03aa7f501170d6aa8d6b6d10789bce750199789b49f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b2145dfde9bf220b2a258e545be2d99780cd69badf97597e40a572d67e8b32361d9446db71ba34b6eb762dfb9d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11fbb7b360134fa99239bbbf35974c9c3c048b52a7178d931cec8748e5f95905c96fdad6cc069bf3e59ce1ab15d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1235d7a111d924fdcf12ac5a45e794a8a0aa2dfdb0d216f055bf8f5123210f4cdc9835010e625aad78ae1bc3a89;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ec82aaebe06e918a4e551e0a6f7144619dd27f1a3568812a4041e2bfc763f8bed25db3979ebb58d8d709207b0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2cacdf110e7f1568bbf11932275596f624e8aa77777c17acca446dfe6c48e1ebdbed92e9e8ad38860ac66a31c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h95e3756abd98f7bf91e667880ce1de2a5e0ae2bffdbdf4ea3b3bee2d00bdcb1c5f78d19ce3d76b295f92fd44ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cd27712420539c3460d935bd62e6f26139170edf39090e19aa4ea8d25fcc58bfa5222911632c886a4af8d2b50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1401524f3b3d73fa22740c9bfca2cfcda569b0dc3aafa14befce49f430036b143fc9d97ac795dd5d63540eb1ab1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h32b2719668368b7883a5664b9a658a8c1abf6906d0fe4c910e5e5b9f63295abb6f8e6c9e4cb5283f8192bf1fe5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d74f6136d3313d4dcb2729672f84dfdccadc518d2fdce190eacb01cef8c8f0601f945e4b820b806025fe98ea09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a2f281b911e86c45e621c4aa4953ec1b75d37f33192456bf5f27d0564d34c8387e615d97ede5462fe44a380c2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h761beee1459bcf3460e29f3b56a5a4375c7457206826ac8ae37ad8af40137ca8ba761946d3537ad83b8e578dd1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47c33338bf1d00db944da782e464fb71fa79facb79afcbd7bcf90feda80c59e175c1d74b5dc46f1c90867f48e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3cec909c17cc1210902684a45f169277fd985928fec78bc7b666aa429a24ba9308794c4aa67206ab7c84c73682;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h107205e549e2efd2bb17e65e4ee60f74a36c7302516f10dca74edd24ce242d51b8955ad113361229890ff98caa9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1264f06cb60847af3012a0cb3c702a7fea1a9f286e1018f0bc09c435d4746ba089ea104faeaabfaacb29c8aba42;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d9d479cf9f610baeebfce16e95232100af7841108c8cad97d5d3c0c81fb7f4438f827f999f85e934cefde0e4d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f4399110d90d7176aade370c68d71b8a0cabb13b7cff7a321d3f303f1e4aed67b30bf2c0686d590f760c76db1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17661c235bb7b6c25314fdb7fa0786bc119079ac6608136768afedabb2fa7948529bd7a14d0d8a6d6936d4e6acd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116674a8d28f3bb612b3800d5b601541017aa902a6fb1653370b333eb8a26d577622d7dd5f8324c44beef64b645;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67647ee3ad6e17988d77bf0f27b4e4fad618b2ee71921e46e56dce883aaf2ef73d8c74340225addda53f4d37ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0fd58f799060a3b701dea0d36ea44c7e26f09a9766ece382a9e8c5cc97cd87133746ed5bd5cd0dd5361efce07;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b5380dca97720061ff9d2f93adbf30e86ae2189aa23eced5368b3eb9089d00bc3fe2402592fe25923bfc4368;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3dfd6fcc87e33b9e1104cb58cc6f36671e28f3d356e1d23ee38a561f270c01e10da7fbabb56c31c78cf7b3adc8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b1ded84e4d6817696b930398f224c1a6c34700070c6f9998d52408aa31c5510736a1894c22784498df7c757d1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1d0afed9b127c10c776d6b7dcc255dbc56daf423a364e6fc1d17cd052043b8cf41c11403f88675b96e7392f79;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed656e7e108b10374137a0487a185f4cc0a6acc895626c4a4973894cef43d1fa017d97221c3594776d5744368f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ce1a9f55376f23c99096189aede532c0997a888371da7ea34e306fe0522c6753e43a4b03599d8fc9aaf9237ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1973d4a68312e0a5ae2cbca674e70eab16df3f1c73f74cbf3e10e031eac2cd43efe517e3a232cc82281e3ca6d0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8fe83ea617c8d6d5824c3047b75df2b3b04d12437130abcc5b715408c4e74a6eb7c7041b7b48ccce3fb60791b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha61935e366fa421d6b385caa3edb05a7eea6999043eb2337c086cd9506693bd09e3d23a8769ba82a58f4519021;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ce8f5fa61759854e9cff813fc8363bed4fa4aa13ed4ae94a70893a80a6e783d2a28c9e35906c4c4402b474c1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a525e5b33032629323340cfef95684dd4ce019f876ef7c7425b6eee606aafac80eb2193774f48727fde677085;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18697aa0eb1ceeaa7fde13d856682803e46a03dd963da6aa73aa1ede085dede38c8d6f2f41e2c85a6b45f2b9cd8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f533ab4fb8a79dee08a6e06520383d79de9298edac1e8c6845cf384038cc45f26723213f091c1a98d7fc4939af;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f533ccdad9b1cf3e805d47a4ae0e4d50880e2ae672e69f129083392bd2ea9b1ec1ad4c250bebc20f7b988f7b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c0427616fb1a3f3eeba931dc0e69f4173b1b26405c7a0f9ea631c47f03dd1185eea0fe4ff17f268a702ada271;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2db0276b1a1ecf8d572b14a72e570adfc2fc2d62287f7c34206bf0549542114a890f94c22ce33bdb2cdffffcc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f30e7da514503cf9d97b551affdcdbadaa86314268795d8066e85df34df1c45139a88a158ed6445c258be0bdd9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haccd3852a6fb16c5008b25147cc30968bb836c9f5284a2ef8fc876898879112d461e117a6c9ea2ef2fa51669a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1732e141e10f1539c9525f85bc4efd943f9441c798128354edc68bf6a8d9b76f094853ca34889c99998b18a1eb7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc42922328842551914677d8018117a64ca32203e0e55926e69e195de395f187c38a87efb5227f8094f5548fd6b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aba60c2dd46dd346d2641ba7aa1e72baee27fddaf1281debcec95d916a848d5bfe19c3a3a4d21713b48e375607;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93fc9bf385d04cfb868143f1587c8639c0c506111bc3a322802d532d1a7756c6a5fc2ca6bde4b8771e8f20b3cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcdfcf9fa0c935c1222b166ca4ff69e6519d1ee949a0796e9fcffd0d0d789b3e1e607b50390f342938b078e1788;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1236549349f7e1d9bea69204f19c85894487e347e13289c9e960643ae3fe91a4d7569fb88d98b418e02ae142f08;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d959effc50af512f471bccfc4a0b736dc85364c8bb1a2e50a8e691768d5de63ccee6b1b2f4a15ab38d96be8a2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6991fb2b268bac82e9d7145325b3528f5184922aff691f3bbc3e5266130f0339b8136f1d67d1e004c6dedb4896;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcc02df965fb70ddb9ce0ebaae73b8f65e1fa14bda747f01eab707c2536b4d39f74160ae99ad97a98badceb3fd1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7481ef15f3dc3cb3a3ceec8457fc0c93cf84b4fe8f898c92b8e7f99d3d07a99d363a5236f61fb0d900d8e403e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd5fba55db64cf50e204ba757d7ea0030a93fba5a3249c92e610040e38a885f2c1b5146e47f1d75fb304cd836a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc2e0fe320e1ce80d6b7f5388b5ef760a2b1ae7cc8a42a5cd039d4b4ca7322ea62556f4f7aa52d586476df74c68;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13fae871bc312402749fe377303d896cb8656fefca5de4e9c33d379b78353bcd9b0833bf5b872df4c6d5b0b65ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1601406f9098694afe6bec169f5a126898181838efc5f441a112c2d00bb66cde44fc3266c2fb8852662ca48c5d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117ede155359a6d9442aa588e1a6468d084de37e4b473634749b0e1f30990d21942877969f04a767523618b5816;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h188d987eb240e481c5fbf4ff040c4c34da8db6782bc1ada1ab97bc2c0d2f22f7821310ef4579786c8099e724790;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18db79bcb56444771139e686767a190d8e3f4467c8f3f06904671dca8d6a4e9db2cfb1eba0e04210628cdcc5f67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h20567e5e3d8195ae6bd00db1b121e3cda3cf64b776b69f40a4fa50b6cae8414d6d237cede36275a0efd18a67e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7ee46284622742ce5fba4e748d62df33c137c299f5b67cc45682dea2b52aa56c6dfa9d7eecc96a015690a7d5f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h148099091f54d0ff360654544a622a3a2ec01a213af9d70630cad49f49e3084b64df0ad7f2ab34eae322738924c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha993873afa6050e1d25a745c48a40626c752da535c8e83c9c7f16bee2553cea270f0afcca4cfdd88ad8581b7df;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25532df7b576c1befd61b787a21788f4a71863d52bf7ea1b01eef651e58691ef85402dd101ddf0da057d10fa67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h109f13cce7cd77aabf55018113ac272af42a313da6dbe22d4e238ec3f90a9051370b6854064b81282d2f906c51f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a856af03ab13c8fcda3f2acee829b77755a9eae3b98b4f06a4a987ec458823f8e6711a536c4dbf4560575048b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118a562dfeb120bd208231361fdfb512bf41a8f66383798aca79b562ef3b3cec71a47b3ee42149397edc1324f7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14aee4c6c068146ce59ffff98872296959c638e09620ddf6bba439d5518ad48eadf55c664cb2cfc677d174f51a8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9afd2f23f44fe9e45d19e19a6edf9e39af6a4c842eb145aabcf63c03c76a28b32384fbe90bf0817ba177b0713;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h151b6e8ba6f0eb078a165c0809904d7d7d21c1267ffd8f26826441335593960a273b229079dd03c7632703cabe5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124eb71250b33d3e746e51bcfbbf53faaea628cdfbf486d40b193e7926cfa53d20a4f1b695942bee136b9249736;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb227f3db4c32baa5aebc08b31678936dc09d3ce0ad0674f87c8089ed8524cb3db2d7af3ff1cd0071961c7d95fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a5a13ee972b4e22dc3e4d0961e6229de4bbcee374f33315217736566511daa3b843bf633b55e8d425d34359b1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf261f89023bab2dd1ec52eeda207edadd5d2bbbc8394df319fa489f01e66d782e1022682df70e1302354625aa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e33d9c1919cc8f4233b4b7f738fc93a25e851f615e1e9f73e780aa9df0ea9cb52a2e91dfb32b5afbe8ae36d6a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ed822145dd1ed22bdf89cb39a91f12bcf094dc666b57615c719fe96202772fba9ea5c9129abba83c678baecee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7cd745b6f59a3fa2b64bf0ac756dca62332d2153ba65b68c88cbb4961de54f09af12d0914c035945fb8f797a43;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h892023b00a06b86f320920e5c51a5fe7617c2c50c623b127fbdc6dbd1fab6c84c3064a43d000cf3b3f2eb477b1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e56e7d7870216319b000591a10a1eda951779c60a5681bc47ce5382ab5844afb3b31e3ad8eaeaf9a511515589b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e8a1dc9a0334194740e52b3f1d02a75a46346d751c9c2ecd893cc5a67db5affae9f1b2e6852b74f6b8b841a3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha939ad4f2df734c1d8ef79f3358c79c77d7cd2195a1a04dff2ed1b8e6bd7aededf88f10c0d49ed5373f43b4094;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba43d34fe43e61730cd656f28f2f4b6decf4308ab5aa299a987955654ac75a78ff66a924c8303534e35538ce76;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47ce4514cf8b679425c4fa8a02e9515eb2589e26eb640a530395b6c57d7860cc084ecabfd1bbc1c630087a8342;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12edb50f2272881c9450ab5161a67deef2ac50dcce34961a1cdbf5fd24ddb110206f348255c011275180ce0f35;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ac10aed1d2f5f78e88877a9776b9fd192059823ac7c224e562c4f03fab483021b88772d9b9a07c5f8b1ebb705;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17473f496b2d679d8db9f2f101d23f80933cc3f220e1701f48dfe4dec99017305c4da981998b9e82f8fe7d0e1b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cec5d0d338acef07ca511d1543ce82a556732e8a2f66249474e96520bff45d66141d5d9469af703cab4b9e2210;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168837dea57b1b8c6e58ec8078dd874cedc26899ba2ac57760ecea62629dc4356c28d1e46bbf87fe9a9d965fe7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a8450b800aeed0f5834c8981fa58270bb65c50fa78d844f514add7cf309ac6073974d39241f7d1be6077d0615;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3c3267c2905fea27ce0dcf388472f153662c0d2f43c692a792864d5fd556d788f7a6ffca71bd6315c28d32b2e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26e0d0fec2bf89fa0a9babecddb0737018952b4fe1a66009cf0a1515f46c2b33dcbfa08f25466d9cfcd3cdd1b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5d71e166cb422eb8b7b04434fb10f87c1af716f4d149d8e61b99258468a1fc2e8d4bda28c68b3d21ef2acd486;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h228237a536f37f47e4ae687b431a451cbe86adfd0ed1dd1c7ba3462cff6c215667f42eb0403268904a930da225;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1697e00818cb41b1fc894da5a7153ecdddaf7c18dd3bea8cb9b5de957dfc6824da387463850ededb49850ae6c2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bcfc24c11d58b53319140ebda4212f087b081a03e3349968107eed7dc77850959ee7747e7ca91af85133111f39;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12853356a96950f081576f1252a5d7091bd8542484e46a9caa588369c43254a1d82442d2d2e12eb92257557c9d0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c1aabd00697abda4a3546c93aca6ef19d89024f005a55794a67bb8ffd6a0141bebb87245d1f1469fae98f4ac8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d50a26e67820a8a6434ce0d3956ee53f006429e53c77167912b3a29bd558f573466c8dd2f7106c529859f3721;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed2d5c0f7f27216ff7b59ca1b168d6aab4fe5350044c3f64eee1a428b018fb243828f93c023df7bbc555701e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfaeb9277a3541d7b37dc640cfdacc942b26646c933c6aa42f750d7a0effa7799768cb2db966f17424e43f452ae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb9f1782b84d16b4fc03c9443b5fd35e5c221b96e90b1178c12fd8d2c4ede2da8b2fd013de0df033cb20a9f80e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h196cfe8eb17c2aade31b866c65dbaf81bd54b791125482834d395e4fe88f8ce43167506e429840ac7bb96befd61;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcc20bde7ddf4b2b25476ba6bb29917e266db2c7adbde75917db1c5e707ef95e3340eb5faae67d44bc1ee9298f6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89911ce2dfcbbee151c86ae5554a152f9488a2102e844127f5b74a1fa4c5f63c04a55b6ebb7df4b994e5f94680;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb0dea7a0af4d0e10e61a67ad68eb9ba3fc44fe1808d55b0fedd8eb2a29acd03c2a06c9eafebedb772ba5aafa6d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36c456eb66f6095512764b2033366dda59f4c655bf997347dc5d28e117be3e9028aa4feee550498501ea72832d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16233f3bc37fc0a30641470b8ee8d496401598387b520d9627b5288bf9a4b83e7441ccb699a7ab98f64d106aac6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181459922618f237e6d223ed78569fdf9f613983287b7aa42b552c5d2f9eb8081f4950516b5c238caa2bc480af9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c33aaf3303da2d2ce1eee88247222534b3772de5da5464d2480a07b6af5b3b04fe5530dd7c98d439558d45f1ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e7df166648cdf79f42138a5ed8029e7607a9dff2cd1587efeb2c80cea7b3027a8b8e9267e0b678b3bd4076ab7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ec7e66cd8f8e220177ebedf06f38bc97a465988b0d2e9eb3cf0817200ce1042320bd6bb85c364823f36538760;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c6563373915549e981aca518378ccba9f25ca8e8637fa854c0cba3b365018a68b4d62e41c1a65e94c522ec66a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4adb8e6d822a5cba909a5a7662879de686f621eea3ea1a5047aa8106f39881d59309b05eb69679f7a2746d8cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h776d726558865931845dcf3af2cc4eb65898d0cc2ebe8216f43b93ba16698ea2eb4d11eabf2b8c439fe0157ec9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc52873ae4b489eedd81cab289eaa8b6361a33f80cc4c4096005307ad259fb953113750116c140866b6aa26fee6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb6da21736931968513b4091fe69956a5bb96a9238e38a5733c3b3fde054a45cd390cd602884fdcd1ece507e701;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f8b1ddddf9e30566a05a18221189f1dc6c4a6c360269cbeadacfed17b3772914e3d76c1026b29af26183e52f9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec3633443916f66faf91ea1a5ef8d7ae78cba06420e8837f00ad18057352d4e16c80f987944c13a3e1dd00f0bc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha63e8c6b1427c1c654909645a433c6e92331d16b9bc7492015375a22e78e9c1a37ddbf59bf33ca9f32285450f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h130ed639096a1ca472b5f9cf0c1d233cbf24cbbe5820f0cca39306a8cbb0c8b79734e353daaaadff8c494409790;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4e32939b0319d201fe3edff4e61555e928489a70fd951ad610cb7358a0e4128877830e2dac8125a33d3f90cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c241002859c05af678498971e36f874062c0c81c33e1c151876d064fd6f0db0e4d329363d32edffe4719d02ba3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a66fa0bd2b9d1af5654035157b499facdabd702411d66d91f17e37251cb4673bef2f57e3cf77f7442e6924ff3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h301a6415f111578c96acde90bd577c8162ec000da2cb4ebc4f3d1cba5be05ba0ed850852a99b44196148416a12;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1788a0f75e3504f40b1f0785fa721bc65bb91ba111773fd0ca28dc71858bdafd48b94f3194cf8c2af643649ac78;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12bba337f5c9d394e55660e9e41498c6517f0174c04135c5d2464dfc24c7025927bd046b9cfc16d61febd417cf3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc9e5cf262aec0c97f1853fef816f12f64ff5276aa60b1d9f7ded50a27f066b1db553cab578f7183196f926cec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122169843d41b4a2014297fa27dbf920dc61cff05bf446ef3307c96a2f9de856dedc5b3744b14933bed276cbcd0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5a9c040232c96c58623936e622af1157b59ee44b031af82cdf2102196a59403b6c9cb6ed058d7a079d6a5d111;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26857a2bf24fdee202e3242d605b990ca5836d7249ea3f67cf8b41a1e8057c2419737a9037a8db840df588a27a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha82639ada8b35c28f3c828ad61a89b524ed27b73949100f24eb56e23b1cc8e90288e4567b24cec922152c3e3cd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d09b5d90962d0932ce95183ae94887658d6412ca749bbf6528256f19fb478c1ef75005dba85767ef42abcc6225;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3d694b89f37800fc2cdeacf8a048d55417cb519ad66e0e5c81a41feff9128768fed0182d6c78001d3d3f39a988;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h147504ac91eb04364ae36007317fc373554e095475949a500b43791a508fc67d632ccf6c0cd9d9d8d50a854c858;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h902eda7c2f94a16786de55ee67a9c22e9ccc53710a9f36fd3bfb4acb679f9c5369cc61f813b53146ae58dd2315;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1972c27b873bc12ea612bca8f4639a477b768a08d349f220a3285637e7ebc38c5d5585d4242857832d1faaf3182;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc423e81657f289e771ca17130c0bbb0c94e030123c5e20db9bb51fe529a5eb8d81e99f2f53b511043c48bfea84;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ed79acf0c24ad1ed7f9511f797ff48ebd923726f632a5dc53b4fb87a3150752f18bb3f4459d4abfcd4d4a3e36;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fac4cf61daeec95d82764c4ea5e6eba788010178327a0e6d9680978dbee913ce121e54e6891bec118058a732f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h543fd03e5487d4fd38762999d502a73ef5bf9cdc13430edd6fb9fd096c4ed56e879c6e992d75e1032f3474921e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1762b4db2100eb6bf2cf483b8e3b945d4efa316730b665b2e0530495ba5804d641cd164c7b8aefe0fce3c3abc6f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b605f558cb7c6049c9091b8b0d3aea32eb593803a7451a5553ad98df119d59fc2aad26beddba7212e6f536296;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f05b40cdd84bed0c82122a74959a15d049d483c0c14a6a98cc3cc3bc5f325c2825189fb4a067daa68541033b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d3a71b1bfb93f86d65ff5624bb9e1028f6b5151bcc8e4d10009f6f61cecac0f4b532c1047a7220a2f76177df48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f0ab3664d4e5449c9e15d06937a718b936169968f0eeac66a7aa4d671b91d3720a49ae261d3b157803f918fa0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7e16ea2124c0ed2d3c3a18afbcb57b9f2dc93d7f2f65abfb7e7508441adfc3750b5cf4b135c6809256937911;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8257128f88e7d1ae27efd53360e20cedd95dcedf5940ecca4ea3f58397ecdbabca6ac18d7ba2ed9b422f33716;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181eac42522a8c373cd5767355f934d39c2f02731cfa336c8a76a37cc2a1a2ffbdc0cf223f8162f82bb1c157e78;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h425241259c77bb21f59c6751c9275de3bd1b3363600eefb69caa7c64fd072ef758ce3cf315aec077f5fc6b9339;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he572879f73fe43baba5bfd28a7989dc78e16ceb95c47f9d30daff4dcda7607ae0430d6e68e49dc71917b8fea51;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16824fe8a40af415e2c7d1e7aaeb7089da3ae60c9ba95f28f644ab62953c7ba93b538ac6c2a18f9aacc082178bb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e638fea0b64ab9808ce0917ece54524ba1c2943290f4775ddc0a8239f2cdf1a581481690a1c0e6193485c5e88;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17816b9b17e07db817919f51502be775bde56ebd74ce2f7807ae7cce75b833758f16dfcfa8dbde216e24c1db18e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff452499afffec7d9582219b7c738d332c4b693cc593361611fe5ea34bc97c018e3d9a3af40e4e7fe3d6c5b75;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd0d6a0ca502178697f6fad20c43603e234da0f242b61fda6d51ee6586c327d711576bef95fbbd7bed2e9f7ca0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3b973e93d7460cbb9477c42f8ac86f04066ed6feb182f668a020fe656b9bec708acb2fb215ec4d4871305440d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha058f38a68c68f3d184c2d07e57d804a555c23fe5bbb13950018778dd670665315d5bf66c7be6387cac5ca9205;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b041a2983da33ec914b536e9046faa6429ee36af30fe330de1dee3251899c5c1e79d7c394951f2a6ee1890944;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1962ee3d1995a27418a988669a2a356d93c2d0297c7790ec5d1a3967c7965127680d15ff14676faeffed809488e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133f28f3f4e44ff0f2a347dd00e360e5bcc612f577e8d80905067a3f1d45c6b2b61ba079833d13185b28418d5ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e37d02599fdef5955d3cf3feddd4f76b8e4fbd9774a9c57b911c0aa34c68bcc64198fca8719b393db19bc43716;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2883479c882eb466b8f08d62e226c33ee107598c65f8a9801c6dbbf7cc13ebbd15b742a206b898e3d12685ce9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h40f8e5c778d85f7a8800b457d1b8896770f8928d960c4aa68b907f1d56c6765ac955df0ca215610a37cfb3c0f5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1598c1968951e5dbfe27ee753db1e3a400eac709b1a4f883de45fdc1089ef58266c53be21843ffd8c45ecfb2cdd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h39cb2e38c1eea6ca1c15fbaf97c268e0eb8942b7acd5697d9128eaa6c77ba511f89a73f1e817d6af0ca7e1473b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c86f239c481ab3ff85456877b0acc98e8e9b13b068b162b0fb830e1284dd65fbd6d41295a30a37b1e28fc1fcdf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ced46809cd2d99932a306c70fd9b5926ef4b99cf8e2ec230463a1790776a252b2028c9b57cf691059610283d4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cac68e96e84de7bf1d01b084199c62f0ee52dd26dd723cbc9c09233ffa8f7074c499517c592b7598df3d3bb026;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5624ac29120d8976e70a5f5e0ee774e800d13c49e07898f0a04e8c2df317e01345d030507d4ac527813aa682c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c019d3df0fe06f18cb67f23318b2a2e44febc636f2a4fd4210c7b8d45c8c1a2bb3c4c722144e77c4783e074be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127a67fbb99bee3c357b4c0b7feb6f9a7741abef35b72064a30123c4387aa5edeb59a610f85f55aa77b85f8d2b7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f12c86e4cba39c4a8964cea85be6f5fdb0978b78fc786b58e83d17587a434f58569a20fb83d0d04f15e954b804;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h46c5059857c8122bffacfcbfd9ed2648829309ee0c1a3aa66781aac37ba325f4a6b880d8ce32ee673306a72dd7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5f17fda22fdfff2ae62ed64f9f77c040cd24d983d747bd632a86f0cf402bc97483a1860ab89eb1c9ad84428bf6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad6e1d7be350f82be4c51a2a9728091e6e9f203d0ab76f242f3a07a6c039f63dd174d1e4012d97a54a6548080c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ddee43d1ecb8fbf34cde4cba7c8d4a8fefc6de2025d43a8043752880a6f7d1ee3d216673e78a9f8b92d8ba8c3b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6b3932640d3430dc22096d8cb0489fee26d316e4ccc53b85d4da42c23d8959485ef892cd01a1f7e50eca8cf85e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7109c2f79fe17b4649909abca72e9e0582219481825c1ce95553e279b71cda63b67497a714db597b031a1ffe60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe6ba66edb18ed988c909bb6367ecb7a04867cad311e983cae4df86d5bdf7c92aef5b430e7a263beb9c3302f99;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be0970cf4ccef971f9ca65da66cce6335bd14264f84f97a0c2d6c191c2a8e7590b880434769c89c8104c9de929;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h171dcec6989c195d1471e638c0ec6022c36368cf25ff8a32509b0316f479e9b765e51ed7d471cb11912983cec58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc00f9bc15901e914a2dbc5c14ab688c0e6cdeaef715b8e08bd8c1cb900b3d270d8d548ee3f3ceb4114a02ca830;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h536020b786460ad00182b3ba1c94df72550c5d58f7a042008c71fb412a5a184a237353880f9628f4b6b19ff123;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14798543e7910be808118279c3db03b6b7ddafe45f30507c8d3faaf375afe6898f6a0bdef090a3f50c5f4dca45f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1948ddf97e94a25dab03c0c2465caec6665d72fb4bc071ecc26355e0ddab0e1dbc7d7d69372cfa80359bfdc57db;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed45e5e3c05fc8a6a98ac336d153fefc0ec2aceef727e71ea97cc3c8c9dcf8ce6f22a16a569aacdc6cf7d27113;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d502920d9f25e43559cf4898926a291ef3d9297e87aa24da098012e2c1c66a394c47f562ff5ee1a96e2e391cdd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcfc335c19608ebebd042f8cc940274a27528a80582049f0e865bc1d75ea6446794e582fe30ee500a35a67ec627;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea6cf0f8cb39608e0b9022cb5fb0c35f66630c338972a2a88177c71b782e20559bd078785e249cc70a8190e16e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c771de3e50cf6d552f74c6a49daee7be52d8fcf77e453d3f9f49713bb93e8d42c02ec804e7a86afea2a9c8c222;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b229ad327a7cf0d36317ba56948f50e76c5d67df66a66d487834a596c12cc37d734e4f4d2217b754e14b8d6333;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175ae7290f6e534e444aebd77e058434ca75742e04fea97f0c7d5de8f193938703b3bc53b21c10fa0fc59db452d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c751f268b31d0281448be2bcd958ecc22c7b53ccccb09c1901d4473ba8a1c8476e1ae720f56da550c579eb7072;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h284567ea4283560a0538b7e31021d566eda39812bfb596755d886f2996654a401bfae6e70c7998bfabf82f3e8f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa0f354efc5c978c889c1523d148d0cb049103b5d4f00928d7e9e8c1009c9841251dfe84cb94077ca4b92075ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h140c9f951d80aa29203ab5fb89ecc50c3cd732aa44068b7cbd46be635b70ee4803cf12ee5d9b9ba5d975ba429a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd0bd4e5eb9389b4fe3ed661c78c8cf2bb06fb679fee6fcaae394392f59f9950e397fccd835e0f526b1c4434864;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f16a9ac1ee50509443922d988dc462fef7ad46dcc8dce196d37ca185a6544b960f2e000d8a5a953fcf47210778;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d2574884f98fc99beaa300516ad1240bf3e9bcd173cdcbed71facdbd167b44151a417f3e6d09e389e5d448fc7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h83e3476d80bda913c612d23684cfd2b83a6eb9de9383323cadd3d9336f558307fd8af855cf7c1838b07113a3f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6599b4fe08b8152972f8b318f4b0825a39b2809833291951120e62adb960ae2bdc3e7ffb5f95bebb30d21519ec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3fd0a714759eacc24042bd1088f091878fc2041675a8ff9e26536d262daf23011d4ed2f61d67c7aab80713af8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2dd5f059872e4cbebb8f9cb8a80aee256a0b2d7fbb203ee3f095e1f98a718a80a8a08f4b9acdb574a446a36a28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5dcc648e8697e11684dfd4dcf184a233fdf1ebb8a3340ca5eafe50dce2fc384f13ecc1f5d5ef422add29d5104;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1df7fe601443ebc4deb1d08b458a64df8bafb8b24945686ba73d2d8bf9afb39d6a22b84c9e0268484502bfad3c2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f905348369b51fe0c4806ede08ada8976d7c2bf45bb547127e96385b7c980dc57c9d772ff101487503dcdef28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f16dd2adebf5bf1c59b6d91141f79be244cf949fc8929c54450b31fe368bc50fbdbf913a690d008995ff96563d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9b6389e580e6815d77e65a8e4d46e911f01b5c964d15cd66f66b0c481f9ed903102e97783a1e53914491aedc0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a0caa6afab2aeb2eb88992a3c78863434b6c5ac8ef3af725db28b2efad4e5dac7ac28b8004c7fbeeb743f2684;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9516c2aaed235f53b851abc6cea87f88c3c74475a160cad94f2046309cb0b61f43fc4526090b15e8db7a461b85;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94e08d0a740e206008bd12ec2a8553cfa9230bf523513cba29291586fbf6b372ddeb4bd015363b013fb83f5833;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34154e33e0b02c7f1d6f33b16577b7254ec86ca687de40d938b04b6c076eaba1036de0d14fad2adfb7c69e71a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2edf004433fa200ba63518e4d9203f89e9406810522646d476203e7974e2105f9a2da90bc94fd0cf53da33a65;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1715558e696391aacdc922a40b8a90298169de9ee2b20a8edc9c6101123e7439e3cc7881059aefdf05a48d2f397;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3890486336eb9af769891a0ccbca2e6e96ed08603e34992b20605f1b04adb8800162db03c99dbf5e34cceeda90;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb008e0e3e8999b70f7c9f859b455fe849e137564c3911f1a9462602ad2003633cfaf5934151a9a8f00b429f24e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f55cba3ecf265c4131445b45e955230e673373352209bd832c9df9bd19662be427f0f495b867b3ee3a3f021241;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha80de3cbc656d23bae855224ffa301cfea6648ba2ae40c93cf67112b65646af0b5171c255118a31c4a086388f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6af9499126d2ef694e3cf53e8ff662891cb96288c9249b538e499badb13fbad784a802ce5940caecfff6e4960a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h113d11b80ec2396d83a23f15123aa43e72e335e10fafbe54f28f726a5379fda6eb08d5a203fa7a88e97d9908f60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112f65cb655fa022193fe0360979a283ed61f5bd93afcc8fb3b0c9f775a69edd38abc8eba22fd2da132e0ef179;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10894ac51427bad0e38ecd1ad50cb3ae8da90ffb62928656c558534e5280cb8e46d046f88f1c2f873dee78da65d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a04b576790c021415a9d7f7bc63aabf73bad3c23452874c477813e201030e8dbaa41f91880bdcb8f7f25f3f0f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e9087b68d5e870a518000018297ce5484ae488aa4a181edc4663be4fb46901606ce480e6d4826afa1e7caf995;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd2efdd6fa89e6cd27cdef56930ccf1c786d555c9d35285c8260045fae57681c38a24b2d9d58bb0b63c04da1827;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a935b6477977ee464c9222861268e65ee14f8c64cb089514e1371cda9c40778de9e6fd508fb7b580657141824;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h863a716f3ddc5265e41c8b46f6d93c979b4049a5595e588dbbd5a98cb04a5d796975b25b320825a1a6186dd384;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bda71aa592bb7d95bbb2f7fcc35209cc1624389db7904cc87600bf5b72a0ca2c461d50aa630013575aa633c90c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd66ee7568487fbd95f822877ac6b3d3d7d5dcbb0296ea2cf4e74c3bc837dc632c252d6e846d0babd53a6cd0130;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c610b4a3198b52dbd4e670997e884755822672033dce7ce5cf69609d3ba89c69891a5c73bcdb573adda0c71e58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h77f9304d14d78963a39a23e34dfb1d7d4739f77a13dbc08f848f10dc2a1902f022e1b1de397ec71bc11e6b5cbb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b79c2a194396cc6875e8efd1c9e070d58680e839a5027be1c5dbc3ebe838400bc82f7e3bfea7342d944044592c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hddfcafa75f2d380fc53f33bafa0cadb4b638ee35c8e576907a698eb13788661601117e2c7b8d3d66dff286119f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c7be1fe2f593a35a83beaeb394e8a8f6a25ef4e20dbdbb8435639e6b133cce06a334ec7269687a76ba485b0bcb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25d3c9dc04dda73eab2d43f0688de440a5b92589b09919b3b6a3a6cd0f2e1f61ca571d403e712c489682df2b48;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd3d502267485a21016847b4ba41fdb8e89a0a501502f0886f630fb811c184c75832d7ca146cdfcaa24e7e5cf0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16df75b5db6f9f6df37ccfa62f4eee55b32d2c98bbba07cd3ea2657465b47674066e77ee523c20c010a8e770b5e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbd7e940b1f651d3bad275e50ff9c16f532f5e7234411503206484d967b403eb95295350f00fe10dc3b84abb82;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha1a455ce282f1ca8a6b0e13385f20f617e25e0da2a4ea67efb405a64d88038b62a6c31cb6497ce84ea50f7baac;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h312e7d9b6e8b93214f2baee6cf962ba18ef07c918f8631c041f4d9d91b67ab2aad0f1a265e72a656669d6bce97;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd0782035d3bcad73dc4305c66808c73f5fcf57be36dff53d1b460cbb53a4cf61246cc8079fbd989613b7cc50fc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81ad7e4983308b2efd6363469337397960ca80642f5cd03377e366bde4306b401236ae35648712f167d83072ad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd3b47a6247e08e3e7f81ac922a0632441045bd653fc35194243cb90f2d400c2aa7802e70bae24e65a4ece832e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he77e90d1fd9b1d3eebdda7f686aaa0210befd7d6194dd4adb0ceaee5e365bd3a472e2342a9f594b8fb715efb16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3bd243cbed43d78a91e8e8600f10e23ed1b6cb7729bf7f14fd9e6e7836de5a0feb375bbf948245d8393bdf2882;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6639d91521361a57076b16208b0f60ea89214f61591e2fb65811a59bc1cdc5d812f19aaef94118dcff6f440a42;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af1d9ff27407f7a41f2817b41a039323770205f5ffe2dbe1fadfa6fcf96739006a4d64e85f4589b61e71068f46;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab1f3a0f787b68580eebc886c2d902d6793692df14eb52d978ead414192eeacc98138e1538a0293ffcecb1560d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4515972361a307bd1fdbbd653ffc9295636f6b22764db4dbb29643b4d04fe675cd3d6a4869495677ac6ea5e67;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ad486a04fe973d79854d3b74d6bef56c67933c108589acab88bf13e8422ebfac61dd8a731c34da6f31934874b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h49d7333c2ae33ebe54349c13620745c5aef8ee234609ad665f870c9bafbb399b9636cc63b8da386fa9e36ebcae;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ef9bcaa41949c5438fd437107dc88f880f8f91c5afbd0ef61e70c1b0f20dd68e308a2f7af633e85903068da825;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1475cd77a09645e8afcc8ec874bccac62edc2b383233b062de3c7ae315dbfb18fe02d203f03544283a05118462;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd6f4cb2b1504eea0df6a380b211ab365b7fd7505b451618bed9118b0ec5bc4a8bb03ac01bf7f73a3a47b6e9a8e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h101703400780b354d47845d9fcae6cdd6f6b36fb6599b88c7d96ee05fd10beaaee8a5ac296743fc9bba8dc4e47a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb016f5b2bdfd10bc73f91b3ec0caea74811b8166df8b91b315947abb96ae9189d1dee38b699e065136e53f11e7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ad699f9f8a9d9476f23342cdcedf44affe3c1087b1e6345fa3cbf2500cffd51c1e97f7285842d782f10a272c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc81b8105852901fe802bcc840c68bfbd574962cedf793f9ee48855fc60c267c6c28ef477e8c10722cac3164800;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a8aa1a0af58e955c52d60afb81e5955c7436bc7480044a2b9a69df7554c0413a69f9535a3f574248802233bfe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f1072589b1d7553910fa9c7af6deb41c86a15156e38e0bb00b19850dd7002bfb4588ca2e5547ba1d27f9043a36;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe37daf3ce1ad657134a8f461a93be6590fb9b60466428f9e4f110248ec69307a1501d609f6d68ae840e8aa651;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7698b737623b79ae6863162b6c50f86320e0621155fd7e545644b45aa4d749a87a436fd8d1fd4f6d0c9c7d7ce0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9326a71bdda7eb1f1df3c917ed586cdd48afa630812d33f0215188f8dea058f931e645c70cf2e5209a10cb527;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h113cc7fa70131d381994609cf3a0d4c0ff2ce7c4caac2ec643aa582c26cd651bddb241e2b334b548023ded621e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h722787d09f92d9ab644bd7f84a8ac7d390dedc80f107305f2bf2ec2788605cf879d7fcc717e5c3d51afe4a146b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1223c9c7037667041a6456f1ab006a6c6ac1854b0a06ea0b512c17d1b878baf69ac27c23f4c993869827fde6729;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1565a70bd54a5af41885d52991e3e5befb0abb9d74540cad79305be669731c8fb734eba44355b0e9fc73e25ba7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167a95933d23062d9d3a909ce681a06fbb1c519e7dda1f3ee833954de5b9f27f496a0d648f6415f3d7f3866910e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f584c486829dc9836c8d83f0d6a9120b44a01b63bf3f875e13218b3839252bdee71f3297c729f54693a62616f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d3f6255d9f1fb5d8c8114c0fb0774efdda904bc015bedae3e3c024cfb595bd5e57f844528b41ba871b7f0c411;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c325b28e05970a9f8e7e52cb3903704717ad55cea413472b7d2d0fe03de67f42aa1d249b75f51471978ac5a4f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc6715519863acf6818e143f9c5955ac65cb178dfadb808ea0037cf1b344433e5b4fedb20640fa2f78a724f26b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h109ebe8f25a372e4f4f230beba60ce473921a3e8864de10902819c043006985270ac912e7f8d643f94369a3fea4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h113fa3839bbda6f78a5064396062321dacdbc426c4f853d620b4e7746cf9d6f30cd798a34f7b784b3fe9b962520;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5e4fe5f851f9de08503a55238a02c85cccaea306147d85f9e8cb0db4d3b2e252b2eeaa6b6a96a542438ac7cdcd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdc0db39c49a30117380edd6b1abdc3f8d145e067234950a2c909b66f5036ff075a60158086b6fbc92452e98ddb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4702eab05b86b54b1a0543478510c5426997d2942ca9cccaf993eb6bced6a34d5e6bab952435f9e60c1a99f360;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc834ad8156092d45faa4d08f0c15cbd5d790b7f743e15118a0b4d834d5917dccbbb88b2308ef63865deee09f90;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1411a00bf0df11e870c9447bde46fb788e9ce648904d95d74db9d6b2627944b6c183b0718aa2c89f41b75bb4b0d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16269e5875be268a760eb639f71c31513c0bfe790891d7f8fdd5eb83d28639ef8836f67077757e71f51070bf70d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4692679389dae7b01c3a9698f3a5987d3b1c3d27770145c73a0e83e3c0b39b51cde0efb42dcd09072bf646af60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4617f37758a3049eb414ecc7c25548d6bfc0186b7f99c46ab56029ff797b72952be4917142a9df9399aa40a2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5f9f0089b40758377f5a3fb761a06223a3fe888f031282cfdbf437301b0fbf0f5c9c2081392e0c1557aaf83f77;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h48ae4891ee6902bf8b6a3de882e76f119ae192bff776ae833806c37969e823879dab155db5cf0e9291a8d5fc1e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7813850747b7940c36981a6fbde65a4d016abb90eaf85d30843e43202c59fbfffb0e537dd42e4c64a2fd169181;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a8ad07bcbb7ff6d23f2a094dd0d6f5274898c34e92673851a924073d101fb24f4a875eccde8610c6d592170c4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb832946bfbd031eda586c719ced9561fce31dfd358aaae8050f0bad1135a5a30386d45dfe4e67e715e73f5467;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7e7949775ee18e264c168b0dbc8784ad4175be2a60ade3a91e6d22a5b386be0b0211aca2dc6f22fc2f87261c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14146ed498557d5af66974587c647ab2988a22c3dae0a67e2bee801af16d8bcf5ac148801199f27c8db973020f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ae51149ea2300e8d8c62a0a7e3c471ee37a89ca50518758eeef7e0d3d104a6eb40be3a91e6fe60da6a5a34997;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9d55752df4b5f09c70f1895e43e248ccaf7aab96e945d21eab32d504bae347a29a90bfb7d6092afa6123859ea6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19810a09690a4f14d311087dab84be18a094e03c20590c98af511f57f5bd61d54cd445587912c2d6d31a87b3ec7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc894616cc9fd6d9689db4d0ff784ebdeea602c65fe089577f3881950594cacdedfb137130768d4b3e8d9d2d0ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c4e2d299e173f115f6f7b5e1d476bfdc1d35fd1db99338308e122eaac67266cce1f5ff035fc90c9ba79bbc0da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16bd7cf08cbc6b473ea7ce8971a9cd15e68ea117232f173228e9fa965e56e538944bacec7cddfcfadd745e968e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hafd91f4c9db79a2f2ae8e163302468a4614f35a691d10bb588940e1d90d036c98038c4b5e20a0eb3d055299637;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfaa105cb2d44557c7a9cbd3b5d2a4d797edfb59e439650bbf522e012ba2c7fe6024e03e66ff534a8c424c4cd32;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha191d759a2ad9042e1c0d9c26e85f9c6139145d28c1171521ce21c3209e4686aa2cf35ad1686e410c1d2003c2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b5ae9d484fb13455ca9663aefaa80bdf380c961cabe764779eec470cd0df7d948337032f70f7638448237d23;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42f6553d32e12b6544f15dc185268489d8bfb9769112fdc666a78c3735da971dfdc0a6086f2c2d8232da0e392;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d85f2b45e8d9363912293f2f5b68e1bdd6757139d210101cbe687d27a0ec1a4c8b1dc91a8248b0ad2a20fd8a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a0bffcde9152cbb0fb8f0ee8920716a316baeec00004a8fe2ddad6eb9b939b19a29e2909aa9e9a1fb6b85fbc6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c83e31116f6b450247dcdd715a14ec0833d4485ab6f4ac5c96a1fe82c05a1d5b823790dc7dc64fb281f000a38;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7471a9c2f3ac51407195b693c4c7366406fae5bc769fb465b1ecdbb252cb0d898a138326461ca3f4048343150;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88873ec8603fcf2594bc32f86b40a98025c6b5fd94b5b228776022e586e98f51a20cca3cb6d15f7f46abeebe81;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1906b29ffae30341dc216dc7c17f393d2c9be0828b2f444f7e4bfb2c34e99d9855daca1d8f1f528bdb62f5ddcb3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143b3b66d9eae7699e01bd3e623d1ac1dbf8bc6f74a1e4fe9378969d01fa668d339126db11166b164697a7341d2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f21801bf1de5efdbdf1b8ba93aa788a784712eb23b3401abcd24d64608805f3cdbcfce3f9bb38e18294fdd18e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17468730f51b2addcb60ef026205d3e4b4b65125d183a019196fce1ef76cd33fbd7e3d63f95a5a9ed30369c7637;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h174bbc2802a056ac1d7f0eb51ea94c56f20c3d7b02fcf7a9579a1413f8c99f8fe042804cbaeaee3f8d261b932c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h149a37e0c38eb182ac33bb5c25c2dc63d16482c5e9ea4c27b6e0ad4a81eb9aecde5a5598b7ada679061a8afd8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0db64f5ae4aa4f86ef0c0883ec030805fadec361b69341afe3d8aba0f1757e89c4265184e94892e9d050dedc0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd08b75623a8f4e42c94794cefcb4b6fc97bed54c0c30271b85e10a7d18a53dfaf6deea6ff0f6b65a95d39cff8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1efc1177ebc92bf28116c835798c5b49c69ed363c46137e42cbc88ba809d596e224fe8f7fbcd5d3d1986dcb154f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13290eac8a7d38e6cd6edb51922495927ee55b4cac54cffd324ed05ff1fe4c84764013c231468f2ffe34f44df37;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16f2245ae6492a7631220146c0a53899d061a58d8845969e3ec066c1677a714721d993596c8be3e81ea64c07019;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f6ab3371f6c12965e70ad2fbbbfe95e988e47055e20a589d8c976bdc1082581ca22c48d439497927ea64ff0fa;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154a65ddbd3d09e6d3a792a9bac6a5ea995e79cfbdbd223674673fab0c049c06ca7321bd8993b3e5e03161e66f1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha5cb602440e1605d911fd0ceadcf031c7b17516141114caf594ef48026c9577a6373b7c5bf5f92ec784ad30a2a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2288cfe9ac76c16b9e79b6a962c9fc2be4b318aea4a5f7f05ce1af55db6027625dd56aada20406006d9ce56b03;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14b9b4aa6ee9ee8196eb4bff0c3eae8981f958d20c6db68ceb9894bfbc3e1f76e9eabf2398d57b55f70ac5ff280;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1904ccfafb47903bb9293db8883b144588ce2611f6a0b1e3eab6f4133adeefe8553d286a63c3acc40489a325395;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13b4e5ea56bf383e216d17c2fd11809a75ba4ca9d368fc4f8e4cb332a1f5093f5ff9656858362a93b2024401228;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1b871f2425b48e2f5769b8bd26172260df363adb989c89c26e829a75aa69c3eb643fd1242905d28a955c72777;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c37fd9ed2e087bdc98c3988a9a97434926ac19b8b6f82fdea2a0aad2e6e9f9d21a428bce1548c2e2658e42023a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd9cc77977fa340860774e83f5e6f5c42edf07b1c8fce5899bdc2c9fcc7c49df21fa36f2385cd02bbaab4e56836;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170a3862d461623df4b82046133ccc9e5c2267d9389cb6d5a32fe24e7d884ab2f2d2d421256753ea8dfbf11f860;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bf052eb3d5139816598edf59b306cef4d9d2d72499325b59d17d3b20a4cf2b764616039fb2d045a1ea253697d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h867acf93f753ee47db76fc7bce51e2a6b4ee724e74267df414acb95775ebfb78af5535b4f69c59d1f3abc52934;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf04f954a9c7e68da775db1e38c2cc2ff9aa05b65fabc33c39fe3370a3817a4953260cfab19338d229ae2299b50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb1625b4db3cfd707b4bbb8cfd810ad8eda99b1dba48e98415a1821c4c0e654ee0bd3d1424718bf13ef036188;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e85983fe23706b7d9b8468326d6a29390bae80b0fbdb9b02612a4a5f520e6487b97525b3820dfa3531322ad23e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he97bb12fbf923ac6e15ca41b644cc811600e5b32756c57192eacca91c11573165884e35cd6da110e3a56aac61a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36402d808045ca187e1f6e5d71d114d94b3201cfcfdc25c1f8325bffee49de038429912916ce949a9179416e26;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18971232551a8f02f75167d781f6e801439957cda7862cfa1300017fe4f2232bf669dfdf3bc28e386910d64b20e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1046e14fcd237d92a4ea6a4d5899adec70d61e9dc601a7fa0d0cb38d3d8e7b78853bc440dc4770991861bfdfcec;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72604ff4d2888f221cc32953136bc29dd895a80c8f8ca306380cdc24eaeb402e066871d90044a7553ed6505c16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e69e64f188962d5016e0cde6eca272df4058f6fde87ac7cd413d3f7d5eaef0ddcf378a7e301cd7ffe3ac93be30;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143a9d77b0e0defcea26933a1d6a9aec9f68ced9973a9952fbbee09a34b45bed73019d57782aca85f43ebb208b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121ec012c3f6fe33300c8c3ec9cba3aac7ece309da69de935a90cf4eb676ed65833e0d7c928298d9fbc54daeebf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcc01224307ebbdfd93dce11d44f1518a088283ca84a5a29e7642ab0ef41300d89fae62bcf55358c211ab5f8a71;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb586c95effbd40eeea799d53d0060f4ad45a00535139bb196e5ebe78810ae741238a8343b1ccde07f56eca349;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd26ee2bd622bd32f42d495c6ba37f1124b4c3dd61dfb451f0d055fe94208bbf18e66d464200b85d15272c8c9a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb01a6d2b64aabbdabd1578a9ebd301a32c83a707474658fa2a36e7ff710b22662fb90b62c518532317778ede24;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9db60cfbce6f7d09ee149f01c79f949ce02caf31c1fc166da3ed8fe7f15206d0019754da96543fc8f627640a7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c462d64ed695c63e397744c99871d4584b83db27d48688c004f0c49f9eacbd96012d4f5e6edcd4c199999afcf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15e57b3bec1dfbf292e22af7f1f0c93594f754a66d221d9f3ac98adea62e7973d0e07e21d0eb06698ce3b31080e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f6143b5f4b921841c0da74ad8cae8ea00717dd07184056c12125e055fde3a56e8381c870bc5450e648c118624;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h91e318aa3ccc8d0b5054f48a28d39a2fefdfc2bb54e53af527ea2d3d5d355d3d494eaaf9b75b658aa4eac3b7a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8155f1abf01436d54adeef9adb4dc10dff79eeb65a870a89e3594d9a12d62146d3fc6f5eb871be08a3b9f6115;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1236c6e212cd43cd9ccf8e9897c46ad07172e44003f01f7f38a87bd73833648b79646a319a4b6716d4e09b3f251;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dabdc13c234fffbddc33f1a891b1e04b6402eab9d917e2db885cc54cda53c52f91eb9f247c68d354186cfe06ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc32e399d2090359a7c32c78865c6c22513131d235d3aabf20279edc98f2b4b7ec12a67700ea57cbb63d2c6542;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16907aa9740b5be480180922e071a4026e22d46b2de840e21463d4bca9407a1691343d20a26b9dce09d9e4cc36e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98ab390a03dae9932011e69332c73b4fb388bc14b9ee2cad46e7308016ed32e54c395db12862ccadbcf315e0d3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a75456b8bcb53a8c8692ba00156d4c0920a6d221073605d5470e66a7ff3fc7d06eec734a42b02e00fa8e3732;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e11780f4c98604f5dc133bfd1b7ce103905d4084f8a43d7d3b121fad8bbd375dc74b7e312295b91b616691048;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h66eb4ef692c00b9bd8eae69f7433b5a49e1725de20049898fa47c570453986480eb7fa002b02aff8882c1a26a4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a924644863ac2479d9a462cfebd78d702c260aaa68827551e82004acdeb44b47b664023a5de02727189f18563;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53487515bc2ba7c62335939fbc58196789877f006af889db64b3be4c8a6875fbd25ef3689f1c5e2c6ec92bf16d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h162fc5bd7db421b8f94a45d2a17be7f6269b817ddc1c8c923b8e6b705003c5c7346beb595bf8f0df3a40e6a5d87;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12b451a4ccf115883691d73f979f415da9ec7ec1c5cc3014cf8e08836b5932eff1c9cbe8a6102de135101d44b1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10005499e7dfc896f7f1af881a2b533c4c4964a922607769173ec1bbf65c69d25fdccf646ebe35d8955071b94f3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad60d60fe3e7c9d93e1968ded3e7ea9669344fe3fbfcd941e38044da962281834e2ea7c3f935ea3fbca4178935;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha29f62817c97385e02145bff29c4f8bf2a781a123c2b361385a6a589e5d5575661eb394f6804879554e79a51d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c5f1ba6c85649bf5e40ea5cf614c1f874c25da22cf09d967d34f7e829e28080effe30b4712c9d6a22130bae0c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1646e3adb3581da113c52f5f9d7cc1583d9216e8f68d0cc474368d230afed41d89559a0d774a9ce1269534b4fe7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197d9ba5271041d1a63d07ab3e925fbe701de227f791e7e11e988fd0420fc4ead635200c968d2cc4c1f418d27cb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5cadb244301148d134d0e0be45bd99fe1603f54f48998d17f2fa6990a295c526726dcf43c5bca9c82d729d492;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h99dfbc945ba8216ad150a9c7176567e8c0fa86f7bfe032b656e5755c1ddf6274532061609a3ddb6def30e8d576;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d131b5d973691bac685d16141fdb21866eeb5f9faa6a27d5bd6ee151af6b8e40b5cf5d415d15dac4979f80a8f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b56813f299036719c98207a4c2c0c0068ca658dd93f6f04687f2706a92a2600790a8959fda75f1050dc2a16544;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7820a6f3ee627b4e97157820f3e9bf269722719a0631a0c030db981d70d538ee0c77e840d3cabb4799cbcb3c2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1f96cd76a7caa0e72beb657fbd40eb6b94efd04a6054bfe719d2ecd930fa737a007b24aa196eabed58f888215;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h54ed5c977d088e3ff1c0402bc2983c201345670242a9765c56508314687fcac05c70a93a5f45168e9d5b3480c1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15e889be3902b0a7a5d0cae45c32d203ebfcdc52921948ab658d581f05010776f08e3a1b9f0797ebc31d71bd9ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c5f1951de978a15e9435b929fe673ce730787005187f050af612d901db5632aaa3f1a9582812960f080b874e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80b2868c39f9057088906a667637c8b99d6a0d01fe723c49bfe36c6d67c0d1351d5ab780a32975c53237c3031a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15893b33d9d0be170ab334069cff5202fb142801141cd3a074f0c4ed151d1317caaf2f72daef8ed918d8cece69b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15653571b485681cfd8a2423e9f6ab48c77641ed6f4b6a28f025ef97aa38c29de718a2d349066a7992bcae87e75;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b9f7306ecf3871991ca37a5ee3adc4fa33ea29cf527a074a79c2aea22cec05d72ce8ca73e065d8d825c9a6ee0b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195c92068d0a640c79c270ec7553d17c356353c78995526c74c72e9dbe08a930d541d57668ba540916a0d0608ce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he5dd5ac7fc80e9d7d2a4b3ee91837c70ac55736fe11c7818d44f7e4fdfefef0d18715b5c713f9e46b2d1cc13a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b5d5bc6dad577865922f756f6f07232faf153dc5224c110b0e3d197947cd64a64846a85c6bf433ba8aed69d3a0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b682f6c0f4ffb74215df00f68dc2f2f50d3e3a44be556573369fa1becab8bbfadb4510938d338ce77dfadb406;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82fc4c280e05b9b2432c026ee38db0fb4b3874e987a7c8fefed14c49a20a7d79ce32e58c67437d91ef46274dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14d9fbeb7cab7a6f723d2b236836c375cf74493e741aa59ee3ff6bae173b41fb99d797032a63bdd9ee31e1ceadb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71465b66edb230c179277f653374e67927ac50cfd4fb87d666add276b938c24478c0b62464552c4df5b1948b20;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45720c26d310e64b16a554c1c754fa18d94f212b094190f2cbff2069e7fd6697f544eb27ae3996d18f6afa731d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5bbd9ba89f25aef473bf7c65bf188cc55c01be62decef2b5a059816bff615c8c30f101905f926b0e58f7b2c4b7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha49394fd84755cd753abd18cdbe73b8ddc80975ec5b1d4c979bdb06f70c9f7c2399b36a707114a80773200c958;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heebff238acf6816079a623466bd2019cd512a38973a26b324892213f9d67e94d93fb03071c34aabb6d67d13d0e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ec1c06c88be081fd230bcb808d08741b9d622719aadf4d6d899fb36214c5d1a76f4606a72c5755c0d4026d2a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f72967f1bc10aa56e754ae753eedee36a26475cfaacc0b301d3f708b9b80f23c4f29fb33fb02d2231e43689ca;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ad6f8e3f575e54b5cfb1df1e1d7fa1dc40c3573e6507ee0f56fcef3da22cf22bebb309196bbcfe5e1c74d29a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1935f44fe2817eba126adfdaa7f332663cabdf8b3e058df9c4db22a55fa9b3ea0de3c6b85402940c1ff832de9fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb687604031142ccb5c533e1594890dcc822ef482ea2ab64b66df66abb7774cdb5511a9e32a48997f384acc02f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8822d5fb40cea594669ee7b5a61d996c0ebad1f9e58081d62d40a931214ebfa811fb97c87e4a4415907b2c44e6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d6f52cee7ca44bc8046857710fe7dddac1d8fd1013834070083fe6f1dfd6912dc95bb874e27df8e23f22b6626;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc2efc94fe3da0bc143c53722ce9447316132b6f95e1a4bd19fd248942534311a4fc2b2e72dffb15d9e368f3377;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c7e98643c8d5882ccdbfba2bfd9266d9c00cd8e990fcce315687f1f31fe30f08a8f7dda8b081fe5cb86d618cf9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d17dc613d7c6ba15cc4c3f47a36843b559a7ef2de40779d1414a1e9ff2c8bbbe34f378198a74bbe372825da3c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a2aa9bf219d7029f247804c1c4dc4b2df07a0ebdeccee6094a55fa0d4307ae06947629ff229cdb4113b4f443;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14205dc399dc8897e49bba9a95f78fd849e9f5f3016627ebc63a9a80aab7b7d364da5ecde76342c4971ac42c19d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3df842005cfbba2e5935a1216b06d0b5143c1f2c70a5edb13f932afb1b11b6a191d65ab8b6fbf196a4ad64a36;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f347d2e62d9a13ec952262165d9833ca423bc054f898c9e94df39f889de3d96c1832e90307fa24a02c9e71b21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heff6b4a546dec57c97bb8ddce77de51d4e0d28b87d46400f38552a0b7140fe528b097f572c795369fff48562d1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10be82490b082f003af23eed022672b0db1aa6586e8fbe04df9504a614bb2e10cd8ab54688e241d3ef81a86ae7d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h32ed88bfb1aaf126f7525c38d400ad62d2b0dbd9f16b6439150dc0bdf754c24a8090d7abcfc214e33cf664b225;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h437e99bce3b6f7933d1d9b2b815acb5fd13baaa16d1efcaff9d4f5584075f98024d4afff831d6d452d2d46f0d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1907d4ab7e628c9b17ff5ea2724dfb898ed16cac383e90242c277cfe7a2efcd408a411c72b1356c968bf83cf65;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c3d84a9deed02ae67da1424b55f59a6af6d411cd39f8e33c0487f84e031648f78db436ecf79caf851ed8614d3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a1a2780e9ac5aa9fe64166608405e9ea8993404014af514acd206bece79a95ae2b9de68cb5e5aaec42f39ebe1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f093eadad31e2f3648c8eb09ca45599795e1d42706d994faf2215cce58b7f3a0611820d312fee054a0eab4135;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h103e216bcb2cb7eaa864b0174fd1ba14a0688b23ec7536ec33b462bf14d3e5117e80a1084e0c38a7f51523445ea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1605ed339090e8fde8081664db0c226ec11994e5812dc78aaedb316544596bced1a399b666f858837924e36142;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f4196258e9ebb8d2298c8909d6d65dc324b5b405c5d02790036362c466dc94ebc498643235c0cc54e455fba389;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a40b7a23c45bf3d2e86c54f90a18982703ac5df838c8663bad8f99b2eb8ee160309e80e7a4253ba5f2b73387c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h98657b0bcf0aee9b8cdf037d96dd7de113babfb09155a9ccb9119a5844235dca7428653d7e86c1916e6f7c4181;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1379db087f1f7420fa68c638ff5499e8b0bae1a665fe469bd98eb0c6c0e1ca5c09fed7043c719f2baf28519c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff56e242210b5c1302705e3bfb0d237e3a7dfa6ed047ae9efcb12314b904b688bd84cd6268e542f7b3e689a2e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1775c6d813daa64cd4ee53a3a75df937df8386c6af631de53ce0caa9465362e2ba38e2dfa39d828cf343c9c5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h712c459c4070de2d9db8777aa11df55dc34f65e0c4e4924aea011dde48fbeb7248c1a8069b96430741c46a9212;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he052a1e5765e004705d88557ecd157a50b52588237485d4009b39d1931a121751962314fa8796f7548a2fa253;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1caf909605b656605292be70428a747425a4e3d9528ec8cf9b8cd15e7731406f87e713ad550f46c8267881bb0da;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb177e6fceda842092cf3fed157bb49e726886422b92166e5f09b6969c46a49687936b08d2fa170073febc264a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d64cb56060a65d4fc0665fc5f30a9d3c4a28cf90a96116471de2b4a80df602cf4736c9911e9beaf4d1e8cef1c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f2269e7199f08d7e8d5389e075c6cef62ff4662c0bab17e274aa8a1f849fbfd1f2d5dc48bf50a85594607ecdc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2deb3a869fc3383159b3d65933931fd123e8e57908910c7098910c11ab5fd419dfeeb35754e1a5e8f38b4e656;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c97e2a530d0d6b2e0e823381d2d070af1e80b65f025a443f327bb0e6aa0d9cbf08fcb7693d00e31f017ac62c3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf315177da94523af663b65978e74f80290561cd99bb74faece76b2c7194e18d9879f91665cb0636644a31d845b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e8aa6648b7723de6e52d7704a8f971d9f87f7a3271653ef745aba397e42bd886e9847eec475cd9da0dcae445c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d624d297cfaf07b8c2a942bd2ba1a3183dd337d5097d1b7db1f60d41d25eb4791120c329708075e4542bd3cff;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3bae8e03c941b9ab4e0e59f7bf7d0dc7ac5dffb41ca0a0cbb217ccf948407508afb238d60316d6e3345f561577;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h85cc12457ad7a1e04483dd04ba7db3968c0a8ee0091a0aa02ee00014ca7da645134e5f94e6e5934d6b0c7f2991;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16fe7d12941b9cea255b795274c3a87d1c6c46217c808c8d775056b0a463131484244eaed2e7b7a163de39176c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa95fe211cb9555572c12cd7325ca66698f86d60c614c50bb3b5355b6a8484bacc46eae374a2a19c45aa61a17;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1871328c62cce2105664c440a9a60c7f2c68964d46125e61745453ca41fb99ea2e0065d0de6a9836b07fb65135f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1475172c38620e00bf1d4ad3b45b3af0ee9100343e966f2dfffc269515dbdba65c07e2c120d6cbd6e72358351;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb0e84c0a3ef5cbcddd082a831119fb04b0002246849fad51d8c8d9d2e20142afe7be4ba8253cfe62639aec7dcf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0c12a93e067203a1df0223b709903ee4584ec43c72d85a70b9bb1805e6776a31aec157e60dff5bff7a6ab09b7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a9fd7313785b49db0302b00f90e4ee8b5b5dcfcf97f667bbea9eb1db210f171f4ed3af4d5184fda83c59e8e8c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3481330ca91b99264b0a3448b175ace1deace01bf9f43be6c4085aec6bd3321da13471fbc5befa8c75b25e8b24;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf9f149836a73e03dc6307db15cf2a442d9caac62158e52d7ff86a057e6b318e02f35257ca67013b55a9a9cb128;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18fb303d9d235250abebf8138563328ab2f1c7a27755da4320d5f616c11731ab5bc7a739959702dab90d63a9f9b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h759e11f0f77cfa70344638a4f0e47c3544107822cd6ccf8e5881af0585dbd1f2b656b06fe17c8575b4c6bf4e80;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1585eaff7ce33f41146f4e4b3c73d1b4e990c33c15415469d010eb3a54690c4aabe35a1a26b29c7a0d0368f61cc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he01fd13317655d5a637e00bbddfd63311006af5ad35b12ea6d1b43820447173aa86b3c83275c047c8b8c770297;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5560caa377e930104b06067e65529186beecc63ce731614771fb0d5c96a951384a76a4235ace5c9b745d245df5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h223060e443ef9724ea9d6aa03fe2c75c6d27dbbbe49636f62947e0a6a86ba7f57349b5c61a96d4d31c0d5662cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e61d8bc1bc57c5887d688e166910c981d66db5471e50a0f2ab097b44c16bddf916e5a79f67bf0871187d10704c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15fd3451bf5eea957000afeadabe31f4f9e5c158ac8dafd3d0795b3b2006b28f53766497799b1f011dd0656a7e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf1169e12995e2384da013159f8cb0b185319ca44ac436f158024f2fe4d105bc9df2c9d31d07ba2f03db92ef642;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0cacba69880de9144479b91a2f64f2e2c30571a5b8564662c52301db88b16f12ce0601114afd7d283d5ba3593;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b198302fb366a2a6ea0301e1cbf5f4811dbbdb5e3ad5b069a554497b561891271c0ad7ce7ab7df59e0a5860560;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd98c449288007bd98a114f2f795ef4c2fd163bcb433006fcc735803540353dbad6ddd23df618d83187c1d143e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdcd00edac600d6a6ad3858ed83949e93a2e7821b568dcf6c6445b8642cd0e4751342431fda313fbdaed5bbb5b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf0d0ae7af1184eb8f157710a079d48cd1575c47e5d68bf9b013e2be8bb7e4d80b800d4cc36a2ea52e789b2ee28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d4f5bf4e075bf9e8db1a91fcb72ae9d126ce480446315dc3cc13264609873afe1f8d74fe1be0af1cdac7f3858;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbbc22af044dcfbd72bbbc541eb7b23997730ac5ba12043fadefcbe7be7ecbe99d6a04971eb8eb626455dbb3be8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e5b278c984da2798c70ea03c7081b54d654889f5a58894370b75818964cd58fe03419aa510452a1fb5f766d3e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4a70e473d3d483981668913e5bc11572b0498f467be61a06f7d86a213ccbef775a0269d63a85f11e74b3ba462e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb42db7464b9c97a4ca8a13976da47037c0e5f2ad29aa0941343eeb96592149f5e0456766ed114af11141ebbb3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a2085cc29d535d80617e21c73d15b6c8b61ea4b75619fad75bbffd99a7a465d8c17934af3889ffc0c9c7aef28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd6b10d0ee544b5e228e3e6b9709cabef9ab07263d91a209a4e067dc67c8f8383994290c2bb2ca0d79e5022e593;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb839a2244d69e202c6ac03291f1ef5c0dcda13e7e3f17f2d4da5be7f32e2e05a5dfcebf62ea2177608bb0a1dd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b2acb62903f41a3c8487ef5381829ec5822876733ab2e691fd8b2b3fee79c0b62fe13e956a2da0f0b6710148d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19958cc760b59563d47e2653caa9a36a3cf36cf0a6d2ed32295635e1eca3b8098e3723a6abed876b4a0b53b3480;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ea1966be10881979d1019a6547d8379025c9d198ac70c70aad1cbd4370a4f23701d9cfbc276686417737c947c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6dcd6f8192458cc0216fa5efd251e0f5fe8e666e8daa90200ff1aaa55a4131f811cabb5d5bee32ab339fec3e75;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8dcd4cd44c5ee69ee41c61b297e265eac3cd40aae675a357ee381b4eeec3d174e0c5dc5955d28025c0120b282c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1149d3fa068ba5a0ace6e5daf4827c8251de5866503cb659054155a1bb66edac352ad216ae99f36c771c6080e60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h22f1f0d1b451665e022b8274fa97fa249dfa4b32bf7231cc656cf86a215905012ef43e4bed273ec84aa9292fdd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17c3459f7b7c92814a8e96619626ed00fd5cfb8e1a77c90e481963f2541095795f50d139f77790d655e9bfed8e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ed782020cc160b65ccc049fd694aa0de5747ad00c1598ecbc6804ab77ab36118cd76e27bc85d895ff030fe608;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4fc49e155219a153be9b3e1e9e8545e10ca4ad5b2aac2876d8ed6225418817c84bfdd07bdd2bb2933d6ac8b429;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a34b645a92605bdb1df6569b4844fc494dbc24b0cfe528b65bea5fe6033e16a34d12b5622697d0bdb3c52a5e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14e559bfbad455fc77718917ddea615b1251e4de69feb0b3caf9701b1323c803584905a96b89cbcd9389f8df833;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c88cef3ad7e029f8b41c4f677920e9b2bc01d54acc1f79f3e0768a97a6cece5feff4426592b583739cc442bcf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c7800bb688b870c7e2ba001c269daab41bb388978462ad5f8b0e5cdffd895093760752cdcd603add2fe1030f0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14115fffe2ed0bf55b591f4f2e54aade6fdc80d01f315f5b4f451322e4cde52cd74524914330697089a8b3882d3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb72b20ff848406bee0c414a5f71d8f42771608ded5ee345b228dcaebfad3d64e41a1f5cb2c73d0d1dd5e1ab6c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3f8ad2bdd449cb37e104c0a26c54be22a0aab8e3d02795fb628f415d77de2679efc65e828aa1c7c24a530e36;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1625ea4fe907f13cf41793b53c2bd403eef08a9922e734d4cd3037d7026ed65738ffa739146e6ddaf5c9f49a2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114210860ac45cfabbe314e18cd421958785b8f3f468eb7772c9569c38f18fb06d41532fd4656a42c0de6536941;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b95e454fe0a9bbcb956b06cd2bdf2a2d80ec8e397bc0f93d2b9dca34268e7b9c513c50ca27df32462844515c6e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17644a631aa0d873c35b2be4c62e02a4996c4653c148d6b2ae0d4b192a6d48643bdf6453d5a3741fa412ef14c6a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172aad84c25f2c0cde097b8da75615a1d1c07ca508d245cd0e501c8cc71168223da729b17c3661981f8d098cf21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he951eddbd7c4af5382429ab07fe64ec5d97d34afb8fd5a7f61f06ec21c3a3936b6a6ae0d46cead01815bfbf00;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h154d14c9542dfe33413c0d87bbe0171b157f2a6e20f4f9aeb3d24f2b04862c02cffbeb69b091b6120382523a0cf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106ce8c5092d42014cf4fe6a7d9f1e12d82e9e1e7bd5fa29163330a37f8e50bf14edb9dd6b7c4af1450959b1ef8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112b05e2e2bbd0f8085959c496673f502fc8f2f38f1831873a97150d8cd110df9028ff1d1f95a26276cfc4c672a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ff62ae3483c460f27d9c0610b03880aa8d6d3cf3bb324deb5344be4ac0600acaca55d860663d1dc2b2be79084;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h181407d23ab9211d6c37bae069633c41b7ba56af98655681f5d0446898e6d89f6aaae9fa3d5abd1c5035aebcbb9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5ed68edfe20e302b13a0771b7d946697a5c33679df3c2c3b93e13ad35264c6d45cb7004755ae66766af1c3d1b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c417a6c62e4c1d7c40238120f9546311f166330a1ebe4f57431415f92c4231d6bc689cfb5d1b5b50ed4ad49666;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128e0905127bcb5624708685927bbd1dbb1c7e33fd6e52b1bfdf821921af109445d2851be0f32db48a13fe71d57;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h174e5704236024030a8ae0da883fff651ec03913823fddb51f2aae2c838ec98bb9c06b67c7bddf6f320f52fa259;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h38f6528362431b27e279349d787cf00289cb2c53b8068f6abfd632f05d44779cd970eca46bc43787e9b62c6c7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150a0fb96e335ab1bc411e590d94e0acee8a7584833a96dd6f42518f1f0b39590aa11c95ddd0ed887e16e12b229;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1614f67a958e766066b8470ff313431c32c594c539f34882e37b79dc15f874ec62b89af1d51a73f42d2afa934e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12f49fefec8deac63bae42c64315b60414328bc3d6f734a18297855be95d6c1051b6ab98ad14660eefae37cc9ee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a74dee92052b68a558e018ca80856b43baf4b04744c246cb4570126fb8a8969b6210ee4a2c541fd1a0c06934d6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd36a5c8a64dad4a57383b857a2733230b8ebc868e6ca62507e9e5c80528d89d6e8b9401b1d41b79ea03f0b9eee;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13cea17e6d729f4b24c13303caa8edae3f259a906418db01bf68831073307b30d508253e7a1f428f777bc7cdca9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e85b8c08f25c4e9c65289a4faf019925c81a3fb071374312d5e865a5a46626f7a26540697b85eec83adc7155c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e4a9329fa85a3c2fd96927360474c6c3256385ef2ab0171bce6d9189758b6ee4cf6e8a15a60d91e24cd40072e1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf53c89ac2c6a8dfecc12ea986b0350b336c6234e9ad0b5074ff18eb9419f0abfcc3cd5a67c9b2ae180a88d6e92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e341d230c2a7d1f4bf282d6119272db4087dd827677bdd5635cc7097b62ab1bb3cd9ed5ca60e1cebb1567591c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82737ad5b28b8d86ecc3ed3a4ff3e05e5872a9837b4a89f53223dd926c42f68f7a6fb3cde25a5355cd49301dcc;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d8cbdc3c6e1d5476475ff4b1d8c28cc4b5a6fe93503ccbee451b731670458a34aa0f6c16a51bcdd3cba6ba3dea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h195ea66727f91badda234f82b995f4c26e5df748c26c162d711f5083c298b9299f080db1d849b1a1cf20ad1ca9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1bf54338c5f30140817335ec2a77c2fa01c3c628d17fa66aac055454cc3f0122256050d50a87a997a2e37d02;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a972a3bce298c804b302d28070f570e98f2b08b7964a3d1e3a5c3a719e8e6e6854fc24b5e906054f93cc17e4a9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1603af92fb868c4bf5781d6b2b371ab9d9d716a6b017f922a96e2e864703109fd8e1389ab43f1a8b1d9fd379a09;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haea33031e94c84a8160cb2dc29cdb9d215595ebac35003b135085b39f9a1493b8dbe72a6f243f9dabf4a360b85;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f36cbabae8de82a933c12cecc3c4df37e09557bbe3008fac988126e20d741d64ca3bb0bcc16764412d3e0837a1;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ebae5d44b0227bfd87aceb6ff90e9d0ae574fddbc9ba38da4ba68dfca904989ec792777388df4c5570da1efabe;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcc97640bc2fee1a553eea7624cda8f017b22f97ed02f91b38e85047f1b301bd84b309c626a16eaa89db8a98e8a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d7a4102cd9110e7619ddb5685ed974c09cdae8d1e85822f90e0c32a7cffc8b5843f6a1764d9f1819f06f92551;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e84d2aa91834730ea67d11b981721193c269f110eea67b11ccedb511872fe3561fe522eb3266a07d686e12353;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c3aca03427a28f0e13af59730fbf24af71a5b4d04370613f2fd1a1f37f6a9a46817dfed16c3f1598d231ee30c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3931ab202507e2bfab6f14498142b663781706fe776afc0cb861a19af3e697f0fd04b4da74f130071b776210b5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18520ca9290161ee79f4c13b4819f9980700286466ecdad32376be9cce25fbfac674c255f2d2e2b4737651cef33;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a6373017fb2e5a66188fc87c3ea91d399c05b37586d2388f5aa45fc92b4daeccdcaa432ce1c455e9532622ceea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3756d4bf817e50db67fa31614a31025148cb35f21b3d6bc9065f56f865ccdfa033af9aebbf1804ff4787322e56;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71da5a90804d5046576b32e16ae913b17328d564a7b534bf7368438358234133f86662f4ec686c6433c378dd42;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa15c759aa62c11b1ff7b926acd958b4e835f5dac38215aeaf305222def27b9413f5f15f7a21385dcd15036669;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he69f823e3c776e3553c68230cd121f148b9691be19e2e9dcab26f15d4acbc2774b18f6485ed314cf6a8d9fd948;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hebeafe19d0654e67972c088312dce3129337ec8158eabf55588b51ae89aaf395151ec80c1ac43238aa67e444ed;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4fee7f7110d78779af4690393b43a25a7156cb302eb36239d5f93f3c4790514ffb0ea8a5bf3e62afa9a7c86499;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19ccad86c7b215addb4271aaa2e3b8db842aee0aeff8bf16e3094fece2a91537f88f41f1e340fcd9434b58cab28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1511dd42419974a82d2ceefa0254d9b192f4b2c75c45158461b32d0c64be45a1171341f6ba6a38d8f511dc474d8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc502b7f331958f20d2ceecbe17671c8bdafc9f28d0b78752cdf14b9fa443bd055a8b935b28f23c8b51830e0a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha2c622e72316cbe209dc907892190729b3aac5ed20d2d4a7c014bff7db309716949e1feb6c464e9f859609f4e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c6059d7e2eaaa85b6667d97028588565ce5b0527edb5902ea1d5602c8c53935e69aedea080570466d769a134eb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he65365e411af0157cebb5b360533780371fd3876768c361eb3dccab9b0003f90ce8e946f78f92c6d1f875dda51;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdea3bde1cb57b69d3609bf10cd5199214f64b632f2615aaf0a4eb04de41acc5c65e5bf5d712c77e19f54ea82e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2dc07c18790c42fbe0ec0e0ad7db2fdc64da12f38fc1efa6006432178185c50f0a473e8364a3ebdfedc23d11c8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185009d600a64a3a161d66035cf026d83885ee99bbe825ad22fe2cc6583b1bd299eaa607f6bff5a1a83c7d44c28;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a1eb48d3d4bc8cbda85f1f99fad3478401437a378ae4028020bc3ce257e4d21f513e11a56bb1d3a421c8674db4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b87b7d62f2a00e14fe4ffefb8d3f73b1adc735eca5e3f48df85b9d00a5063ff6ee462cf0cc3d6d19a81a9c082a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed93b892abd1346aea9555f0a9911b88f273201e963d4f56da555e01590ed9a2f9de73c14218be456437d88ada;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ff64b20f57472d181bbb15e0ed97ca58b566bf647d1e11c7727452b6cad178a44884830e326f0b7f07113fcb3e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19232d7b331f87cf00eb448bd0c3f036395506e8378091df4ae4dd643dd836839e777b3e2e794fb1463d4d337a5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha61e55ed25f2cb3a0e3b18d83321b93d115c9d19413c3a773ac1583c29129baa3acc3d94193260d4040d472314;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h605e2965c1516651bdd5d0d0794196898e6ce13530ca62f59140c1d06557a3bf3f247020c66ab25439cf91796d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42f80d607b048808ed7715604b2dada16c59273e559de771d4a9e0afdf26d8ff41f8db85070e9ef57ab4d80c2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8c3fcead5ec0a011cb1fc7a0887a78468a6fbecfc41ad350a68495194c45e4e8820bb60ddea50ecbfe655997f2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h115362f8425da8192a449c004190239c7a0540221ba2028402c8cf4b70fc5114ca922a5bc9c6572ecaff68223a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0a0ccbd8ac6448050ed7ee9f2f01272ee8201dde735fdbcbff4849ada04cd95cff9562335401826d3ea6924e5;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43489a1aab2713469c5442098ded1e53a5b0212c0a682939e9b3c10dd680f1c1a4deefdd06034c766ef4d9149e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8982bb1af0f2760898d41a7152715710001da1fd375817f68a199e0eaeab116ec701b82bfce36fab70af77cdb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa158051a755ff9d5ebd8250d1b0435ce89c635c90dd687421557726ca28f914d2294f1335502fad181c7d9300;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7de03b3d26c07e82e38baa49d43ca505c70a3a8b8c206f82077039b73e8e45094b2f2b77ebb175a04c688e02be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71209b777dad377d49e3e103421b0d8191099f22c7d340a950c4ba540ddba47fa93192216324b956c3adafa440;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8d01c97cc4a9d841ce840ea9d78aa505d4593075a1ecb57d47df773a23fdd965289658554b13363268649a0b74;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f2e3e4ce1a702fd5698ae32e6a39a02ae677fffb0f39c01e21f763dc61d1fcebb9c02843be779b6d866588e60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a06e81dae4ca9e1ec051f444eefc3a78ad6704206c1e03a5bf79d33bc289ac1b9de7d8c0e882d788f7f3a6811;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d7c7c27d3ad6da801320857bf913c3b3112f4ba6937c9bff55a426cab512bf678b1e2d23aa74b207820e63b58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b545ab1573e5fe10e6cdf83af0ff8bd728a561b5ab88eb85d82f8e99ba480a47e28e4c147ce987428151d87aad;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h562d6406f3365741f00984fd4d23cd8eb3ab02e6fa0715b894042df7b25e79daba21a3ddb09f3dd061f72e83e0;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h174e53fbbfd45dc219098c4384e2b7d4e570c793b9c084495051c4cd949a8b5b52f40e0ab0ec071ac113aea0cea;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1679f9d1f5606a12ea4eb12f88e17e79f8fdda9ccd59a67386f7e7e8913dc690c7df65cf40c491c53f756c5bd64;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111b1c802c1ee3aa72d66b3fb43afc1cce809943c8a2e76cdc0248c3907825fa188f166fa955ba5e9e893a4e150;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3e42b2d1ad2b1ca01a25b20eaef6fea5e61a6b90a2b26933bcde74fc9d638f2e166a497f3233cdefcc78f6f7b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e7474a1251c3f2e1806a7baea692fb51c87fc51ed39d7ea0ce4d4f2cfaa2ac334c862d3f529a9a80575e463de;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10051bd01b5a4df447f1f1611a7bcd2208726981302bcc9f8c0590c8cfbcc0df4cac64f010b8de4ff04f6c71a7c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1482bda59828cd3a2b42fa0ed41d0f64d2d438c405d71296fa40db21ccabc6cd3713d1c5582094297755e34c871;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bc699bd1a43bbeceeb414cd10b7fcde2c19d8d56b2a69924eee27b5c54d153354c8e94f8ddfaad040935ebe7b4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1335cd74d1cd3ab7db0fb1e957c6ea7d5a8765fb5f9945495bbd85122687517dacc0d9b675bac73d91d91fa5948;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b32b4d4d6a0e8608605a3a437a59232de8cf133c5cbd40492abbfb0d963aab130d4b9e7a3ec7d0061ef4d1aa3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1523cb7701440501bb57ec7b214f38af2afd5ea5cfc1b7bd5df666ab849cdea845cdbe12b89029bd45942e5454a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17958e4b9d17dd295ebe38401d539b75f184108093f8fdebac84864dc38d3ee2118d2feca3371f753cebf1d6291;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9bc7e32d875b48d0dd9a62963981af8356ca3922c8d6fba869c72f4ed9d702a045c676012ac26e56b3bfc5fda6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h105db238e5411880d15ccc1708c5f0a111d57ffd3a8a428e669ef8045a7f992a0ccc443626eaf551e66f4aff63f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a6ba45673e2a008eb0cd75f9725e0d6346a19ddb25d876cc318e7cf2224f41a913483f0b730b2a6c411fb7882f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha040c24fb7184057cbfd4a018de4c025456e842b5f4e6e18bf9a1db0422aedc8c681b96f52d93edae5d4956c2c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c6e1895503403dfbd468f15db9be14ba1adcab3a723a407039c5815f31c3bd479c0e66fe160ec89abe7ebb38d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cde53ad3e80019cf44d1202cb433f0b3d6adc377eef7fa464154eb050c7e1c1cb69590af35b53305932c55db4d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ae58e5c2bddd9e04328520d3b5ae09b3100756f86b472aa62b8fc58120b20dbc0181c1e617e59dd6d9f4ae549;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1433e52aa86ecc44f0218da103df457873d1a8d1a5383b61626d6461e0850fa060047e753991ad9824fc6ae6916;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17ba91edc2fd5ba025162b77b254b7c0f96df820059eaa793492067736824154145caf25ad313597a63dc8ccc17;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdcb8aa50d1d7e5098ed97f19ece874a4be2f9eebd36faabe0cc4352ec951c2ff22587e11bc9f5a350f83748a2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d55a722f093f7d2d82a12e0d086fedf77d023dd263af97a28cb8300fe1edefc5ff2c99002592ba8c0353e1b50e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2e30cb863c83b9c4aae2cd53837d664429f2af123e85b1497290a19e2e56e02f256ed44ede97326e2ac0d41ac9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121137dba11c8b4954eb077a0291d0c543d75feb82bb1d183e6354f386c09258a4759052c5601b47b7fd926177f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12f774071f8b4fb4f6d0ef5713acb05a28ca6b72b07368cd7ea03cc97b1168103846ea02c48badc0bb97dcb717b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d608a3c0ac4f7b1310e90de29256bad505c9c93bce22697562bb01e4c2ad00f5ef535f9ad1f5444b027c1064c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146f780b32bfb86703fe9e6f760f8cc522b7b579ae1aed4a80e87a3c5544ab4f2c5a2dbdcebad49a82092dc3329;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc375b087ae7e7b4524736a7f63cbec23510cef06771b7eac6f8e170cb77e2e5eacaa68e25d91b1142db700bc4b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a5ac001f4a3d5d491fe4e2cb3a265e71651cf3b3b772cb63608ad1df724077e69190c093abf16cc7a1b240f2d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a60f4b4a4bb6c00c716fd0fd5cd2fc783a9dc0ba8a45c88709e31d6abda33148d52ed2dfea2b42f47249b1bcdf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11209f623f090cce4c79555d9cc84a55ea7027d391a7167acaf74ed11541751d60ea235aa1981586a1c63cd1f4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50edace8c4c4e6193455751e0325bdc4ffd2a71128beb3999da1978b03f937fb7ba6ff1efddd0c7fc4f7531674;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he7f0dd2177df4ec0ddca04b7f93973b5362437114e28b0ff1cdff9cf4963f5ff50ab2021a9aed0952b71eba53d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9e6816c91c12bed06e44fe888a0fc580674fb4b6e9ff534160c8f3dba5dff0d52a803d1e4e369ecf9a41bd184;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb2498e688b870e7a9028487b8fc399b6702f1aa39bfff338d9931528f1a00c20e86072c20b224c87a11bcd01c;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1039b4de6cfd091dd63f034372479096184d6b3741594e077ac713fa313746d95ab9a83ba5e2a58083be183ac87;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfdbe7e65ee16dc45e17ae8eddee174be7a7aefe011f639eb05cf33a04269ac849f774c40de107d37e7233fef16;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16137318716381c3024050cbde97460a72186d24331d4ea58cafde629c34484d797d547a48ff79ad8ae8315875b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175782ece64684bcf759cbac445a0259ac78ef46d3d20ea7b2854e7350aa0fc42c3238bd745ca3de2e9e1c6b193;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d176fcae87b15da5de4df88c3efa6b75b850bb8abbe4680d35e3935b3a5c3e7cc028cb091f57d1597b38e38e3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1040b5901d3516884ff712a90ca9c07e01b5583722bfcb4814baf918cfdebc94c2d3dfd853a2440e236d4187ebb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13307421450580d966e4cac2ea4a95b0911c547094a2d734fdabdd9b4e81d80d388aedfb2a54b20c1e82764e940;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de0270a7bd25303acb6be685721b61521a740904ac1daec8989b47ae112f591b0f00f71192ba4215a6f051066a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbb22b83b9f7e8fb69c66d757bd869b7c5387847a549b97c53730464f5b8a7d59503385aaf902b3717ff384ad14;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h577ee81451eeb1c6c6532d83b5cc6a02740984b98467deb637f5ac41b6112707f8d0010c4b1fbc3968fc3db656;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec577177107471d75b40e8955a1390cbb2a4120feced6bfd7ad3897ecc7e4bbbf2381fcb5afad31db788b3f577;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc924b44cb5377954728a47c6f32777a66e96aeae44c82b80f2a30341b61797cbbd6bc769304d1485fdfe96246d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9ec22534ca7afbddec2249bf001e51c30ea495cc98a00d7f34f498cde7fee272d06b6be0c8734e943db29e4970;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182b9538c26b0d992af56034ad051db764409de25dd542955d68b935f137b61ae40d97e9b6696f155e4a96a9397;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8346693d1940a8da0b9f73d7f779847b2c4e77425e188907f959ae69536339602c5f6709fc46ef5e31676e2b49;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb822786839270919b5b1e0a01dbe599877fbf0c8da773dd1e8d9b1753f3f3e10898dbf312a92095c28256fbe76;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb6fef9ee3bea3474c199c5fb83bf84fbbfd01fef380a58eec2e6f6ce247958711881d33662310d394351ae373;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19171e693e28811c929a6039c09ea32e347d0deecc199d2112212e88b65637ab054f5e536149f86bbda521c050d;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ad082f885f536d9823b2c58700aa9ee6ca51ccadffab43c241f9d272d5d4a522ecee93fd7cf68632e45b21b1a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fbbcb86cfbaa27c9b5f82862e83f0585ae42afb220e6f2d7ba5968868801baf43d6fb4d41b6071ebbf93df2e2;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hffecf78d7e6ddc991271ae42fd87feae80e70bd938dd2dc2617b5b7c1bb8b9dbeab6073202815693048493a1b6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1292a12a17909594784d96ba6d89a2e6abae58234c2fbe37aaeb31155b5e3ba3f4f590149ec3f5e9727a3c04eb7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165c7071b8c1c7f79efca2e0b66680964e2ffe2b724b78b0fc6f00c629d5751fc260de88ab2c689383ece472582;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1902132ada759a29e88cca64f44bd5f171380b11e6eb5980f077b803e287e58cb6b15fc089a7405879988286e92;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14dca94dac4ee4f453e5c607e3749c0e6733658c9059a0653ffa02e0db35538f614a4b5aed04175515e73065579;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb8f6f43227f028427c5a45ca6d7bdfddab34a370f6b59910db7a9eb6402aefa2b9fee20ca0f7938be657f3ab63;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88ead2ecc48eccfbdb1429352226ad83c23cf12afe7b2043f7d0abb1307be134facd7b9bf1df7b3a5deef0c774;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e4b53a026903b68a5cc5bea60b55a3632df722dbe818e682a660252eae0bb3e36a493a5abbd26563c4b4c6bc3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108463b3fc15019637ea1ca25fe4bd5bd27c762db46f1bc65489869f697337aac27aa660ef323ba2dc3aba3e8be;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a01d3d3201129f9e5387e038478d3f7f99bd4e35bc8e921ab75067d4e27a66742b387885f236588f44c3f9d814;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12fff7ede103e2f0cd95b49809aa63118978385317b72dac78cff75fe93f08cee82e68273eeed024ffd5411fba6;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16fd0e0f43ab51d3945d6583745351d678d0e4e722a46100d4d77d301d94951e6929100e0185ada47b9345592b9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185af38112cb76aace19a9bf3d61ad79dc4c4d7da2085e638fe366ac63390608d6e7ed3eee0ea833636a5b0fa40;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1823c7f103ca9a2edd82393d3b2b91c960a2ec27fa4b0298967a448b4c1fd08faf2c3d4f28970e35d329e2fe403;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e74e4b8bd7d2ac19433396d5a29011bed2644e692f8c043183ad0aa9a7138715032dc8fb7bf91ac489b8aa33a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2a34fd4ab184989db41590e9b6310cea255ac27a54c07680c45da771a9e726a04c4dbacd89ef659c94b96fb58;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he0c5285ad15dd0cb1cb2b7999f156692095b996650c2f552f5abfd7cca9901d9904588d71d50adb1e0c91d8cd7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3e982fc5f2035b3ef5e0590f4c803f82b0bcb90511acbd4061647f24323ae4b08c17d62f511683737cf6780fdb;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c8339469a93cdf71b3421ed758e009845c9f749adadb814cf851459ff6b1c4517555eaec4092db3738d6bf8504;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h123dc8ece35fc6a0d5b5c7be14c4b75c782a4c286459b8ef9d206119845a9627fc800dd73b7e8a3e192e7e3cb21;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h74d3c6742770f376f61f03c00cfeb6305195207baa4edf7fef2bf8f01f9e807f99303929a4e88bd704e5da78f8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dbc8c9206de7986431444e39c5d87bd512fed1110c37bcc087b542e135b9101da95bbb7f82dbb2ee17244bd44f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8e2fa53ae43358840a8c6cf3f2a2beeceba0a510a2fc04ac74d5f80c55ea6423f57ad6108469f39dcc108bbdf;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5ecf6af9a52ce3f6a4d71f05762ba64a80b3789b0568a70e5c0a98bac906f623130b3c410a5ee9fe58d1dc0e0a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4c7165da5cfddf0f80b368a193ad996e19049a7b48471d41700ab8781d6e03bbac8a96760ea76d77ad6e7066b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h166d31110ca722cff542417bba1eadce127ea47fa7ac02aec5e6e06b3c58e99a41e4647d211c18f14c394e64c50;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd7ae4b2d43d17aba92257f3758502c7043319d96f5619506212167bfe028ea455867bfc97753569d3e7ef4fe4;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h288a81e8acf6027ba3a20bc4ec58bb2f7ee10729c495b1d727e17d425622f31b7ca1d5cf1a812bd79ba16f4355;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd83f76e6dba70522967fc3914eaacd0275f7becf675c6a9cf341cd1559c8050257287ebc6ef725feb3e7cc1e8;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ff58c9830aa9dbcf7467938b7b5fade67e3d91dd377411845c0831fed636bdf3332e13196aba5bd9d2057081f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9bd55f81076ed0e970a8f1ce804e9329f1a48ea20ba45e64fc2c23a03ceccf8817d3211746805c22caa6d53e53;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3d2c60a486585c305180932ff438c9e005114edf56eff53761c05f4dd57b80abfdd75edde70c3c1bf5b5720b3;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he085b935f679b9bdc9e051ed294174a41f902e472c95551c3a70903e75dfccbf1d44a8c5e694f35a582fc71788;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfa4a5dc7f3189bccc8086f499289352cedc2f82ab5f6fe4c3cb2180eb84c24a7e830061a64e9ece727b297a4fd;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee301fa11b2759d70407afbba69571dcb3da055867ae7182e92db47e35e6a7b01d6dbe4a1aa6bde9fa416f296;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c794ffb323ae307238fb13f122c5dd759b5ccc2a9132a377721e5333ae3248e125f1c5de04dcd79f43b35e7a6a;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd579860a1472d9783e41a1153fe58b648d72e62f801ed611067e42aad9149954f8ad84a0300698ae3a76a1e4b;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b70cdeb756ef17668d0402046fa47e1623021f1757cf63252c8fcf3aea8eedc0d39725a5d8edf829a4fdda66c7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1135e0611bb66bb8313875f8d87aebe894bce0c77818e229aaa310a30e6c8f647bbfe3eab365e4346a5aed5741f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc699ec83d1af09e95ee66c0fd26fc7af9daeff5785c451814ebc4f490368a8c17edf21eff8b61601207017cf44;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf2d033d4660244ee5d61b94c2bc62b050161a9dc675943b8dee12f677a209f6c732d84e20b0e979b14c555de3e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h578289f55eb961e6e97b28667c15027169ef9694030fc9350f67bf025758a820027dcf60ab25ae81fc6cf33607;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b17017b66074eceab35a0b51f3f2c77276868f1e6a9b2dfcb385761c5d92146613d4c04fcd7d006cc8801e27f;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14fdc9984fc990edb4a30442ab88139c0df15bf433e9bb1b540a444bd803a57fc87bc3e985acb94f354dc9a3b4e;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1164c996119e60f5adc8e714ffd288c093dffb02a3da057f305eb6ded6fc2977580138f308c0a5baded5099ddce;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16f969ee91a9b706fceeb099675dab3c72f8b9e4df432261601b229ff43083ff5a1b9ac91cc12ac91735d3ad6d9;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11a1af11344b02edfa06906ebc7ef6dd06e5592f54eabf0e3527467da9c86a8e85aa67e7d406d1c944d8d621026;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4071c93be92977222dbb25e1aef7fb42f9a379cf149c47c905fa5f73076643abcc3857bd6a7b1e1f47a0f9d639;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h32f9dd7733ac1c28b92b0a2a5e5ac68263e109a2519ff7145443b385968f025aee6a87e1346cee8dc6b8ed1ee7;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128c9bd0f7f7019b1505f263f7d44b0dad04eac9a19e027b7e36f40d634be57ea4eae278c17fd076af4823ef621;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14587fb88a5be2cf4b1ef0e8d605f065ad02179aab9f9dbaecb682b7cd700f889afeb3ffc3744b6326dad209368;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d30f760db1c4c9a0f37b0daad49a800d316718a48622379599e8c85eb8d2618c122c5d5fe90628e6098dc94e60;
        #1
        {src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142b7f6890ecbb9e84d2b6143f5995e29e196572763ec8ff40e0a42716d9fde65890054e15edb3606b8d052a57b;
        #1
        $finish();
    end
endmodule
