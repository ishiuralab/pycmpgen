module testbench();
    reg [27:0] src0;
    reg [27:0] src1;
    reg [27:0] src2;
    reg [27:0] src3;
    reg [27:0] src4;
    reg [27:0] src5;
    reg [27:0] src6;
    reg [27:0] src7;
    reg [27:0] src8;
    reg [27:0] src9;
    reg [27:0] src10;
    reg [27:0] src11;
    reg [27:0] src12;
    reg [27:0] src13;
    reg [27:0] src14;
    reg [27:0] src15;
    reg [27:0] src16;
    reg [27:0] src17;
    reg [27:0] src18;
    reg [27:0] src19;
    reg [27:0] src20;
    reg [27:0] src21;
    reg [27:0] src22;
    reg [27:0] src23;
    reg [27:0] src24;
    reg [27:0] src25;
    reg [27:0] src26;
    reg [27:0] src27;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [32:0] srcsum;
    wire [32:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d75b9f44c2f81a33ba6212527e77a3522040801865da15127bafa55b00b052077f4d0d08f4b06c1f0f3561982e9ffd01216af55ded22ebd5262aca104e9e47a126ed4ea9c48bfa136717507980e5c3fc7962d1c7f64cc6dc5b2ebdced3ab80e5fa0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f6c97f283db0cbdbe63d3d88ac88a5ba7e4a57813ffcd6430356b0383bcb4402a3fa5a2beb048b64af846f610a1055147f2c35e0229aa92e3dfaae9a40058a968f8a17c91df75c9eeea20fb74d0c27e96367917c19ea2f9c3fbcf5d7c6ed14fd5be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3520225a0fdb34aab8238b97c4220f86a137a74026a6f651eded0a1f035a734cc1fdfa5cbaebf820c2ecd64e5c19998b5ee23d2664bcd5e22e367865aba4a14308797044b4317dd0f2c3fd071f14ee63e8e70d0569411df5d3b71e736eddc977747b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbfe5eabc54e390cf6c04cd3b906ac5c35984c9e8ed71147ed37d5d29b360c7fd400e1a319983988d791a65a437ab9e94dd42ec8bbeb1b563ab4f292972d9a59bcdbf377c6a6cab18152dc43ccd283c72f48f5967d8c9ff18f9f082b4bc66984b39b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4840df95ee574467ee13c6b27202a731c1f8686a5ef61323c60650e7b2b00bf36aa4f71b55b575044fc521c76deea9ccec59694821483a60c10557e39a34c7141142bbd2dc9785eb95fb7b2ce2eef5519f4f3aabcf8d1551921556264ae4f647716b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0f0cc5cedb03dfde795229e147252cff50019add46bf56f3ab14320060c7aee34307dfbc2a79ccdc6decd5a3b18ac8c1c469b9fa7efb1184c73e3652aa593600012b28550c3a596eb77aa163221790f9b18b1e9d7cfb8c338f02aa65efcdd8229e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h479c0a32c6bb55e72a689e672acb8c0e519ed044455e18d75f47f3523769c85f673e01ea433f23df4a2988963af4c87390bf4fd2ad1fface3306a5c56e9406d3d80134c5e29f2ff573eb9437d1278e9c752e39d71d6ff437becfa3aea343edcd7687;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha42c3841765899591de96506e5fd889e3f2c54310dea7d0464dc7b49ed124ad54d5e3d7bde5acd4e91924397800c792cfbec179bf68e5b501dc78b13a72bebad0a2c9c9e685a1409b25918136f8994b15caa14d0d129a721d3dbcf0646b14ccf6292;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd7cb80f9d86d471a9e0965485bba9fa6cca8959fdc95aac8a6d429e525c1126e1e25ce958aec49424ca0b3ace3df462211a5ee403091ed4c06b6c046e4de05d2e619d3e91026b86a7245125d267fe4d855b16dcb0d07ebd2720483c252300147e2b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f37d0f88c54bfc8218ff57ac00163a4a947bd41cb59bed20f5c2a19138b48728228b203418287195a4f06aaa7cb5be9b9d97aa91e42d230c9cecbdeeac0d34d1f5b996edd25700f27c460227f1abb059ddc646042cd28860b8dfe986b2d474b22a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9849f17fa0dc4c18160681b3dac4f1301e22d76cc5d2bd1b1299f54e40d8bf175ceeaec46adce89e1a763fcb575d2582cc59940f3a0e2364a5d8369e0b00378eb3e5bbff3a914ce5c20cad11894ce5c96138d9cbb759b9be1ef0ef4a81f8e3cb6250;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb93149ba2f928933e56599fc0e7f4b701413345149f8d291ee1a0df8d3535987a5c7cd5f1a3846aee14f011356d6ba2bbcbcf25968c6197ac279cc09b6ce628c680123a0025314750db31c73e703997b9d1ae064bb864ea46a274c5b9e0ea88f4602;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2790e463d684fd3517d9bf5c13c09e4ef28f39f6362012ff6a78232aaab5c0aed721b910ace1f3198cadd031539fd5778b71f9746a391cdc0ff50041b71dc762f47c874e1b89a43fa81555bab33d9ab755f46467125da927a3037dc240dd8598c7e1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17be6079b6f515dcb202877ad4b267a61d77f072d0f43653177994c3aa738ab7bdbed3f16fc27e5197bd7e1bb8d6a0ada889c24b5ddf3578fd3707dc8c0fa087d3495f2be33b79d2a0e2d7155324c5c1c7ddf3d103219cddf0bf60f7938219152995;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd8e814dd02dc0e9ed1a5ad1574cab2c15b82e7a2389d74a4148ee20944f8b89e0e74535fd0da876759d8464100d652532b715208f3b0f7fc27e6e9b82fa214e5290bbf316fd1a7fc56fea77735a9d1ad1445325059a05da6e8c91ef08fba00c8e64f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1aa6ffd97074bcfe87e20be731b62fc402fa09d07cae6aa1cb660dd514a12a6b6da73fbac500f73740ce303450d908255c7f94c020ccb01d98ca6344ad36fa1d0571994c63fe18dac037ab43f3d6cfb6af6d2b64d374528e98b710ca4ef7d249aaa5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23429b1f6b44ece0e363c664bb4324f96e0e04c52e25fa4906c9b75a79ab8eba8e005e720bc40cfbac5041dde5dff11f7d2559f7801d274f3d061aa536382142c11804ac9db70af3d11f5bf07e5eb8568346974bcd46b4e3f9c721141b1c543a3250;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h322f840176da9569edb390bf5a4e3a9ba5b98f76200c5fee7b405d59372398d0c77fa4d9f39549d6d2923c1e8123d847284b8e253a09a28ad586237799734fe7c396014b163e85e6daf544714c0b4f9829cef90cf4b86da8ac1b0e2539352ee25f21;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf9b0837ab41e6d18faee4007ac71495761cf5e2dc8d9bc4a73ea09594a1d8c958b46a29543a59b6a60221eded0c88634ba7ec59e5eec1c72595cbc68cf0ea32eb108e5631a0a467cb47edb6a46a07e388e064a6272b5905f225ba29121a149f6ecd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d7e729c00a8cda75f25805cde942760671377fa97349a5b6df8d226e51189f05ad1ee58610f4b4aec88bc8ba227f321550e33c59b509014a12f97a63949f3f5d87256b6af04f15db154326594c5e664bac4b377314af795561f9b839b68f61d0b29;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2fdb7f7764560232c6f601d8144b71c6ffdaca4d975946af85f2eb29868ef630b06e110fefe9ee0fb36e05971746f887229410d4c8c1f89db55e2686943de26879f97355721fb66a56b22b28949720d12795ccedf1a299c75fa03196165a643003b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f190ea97d971714c0cbec38e916b0f3aba5cfab28f64120f4bdc79b5f3e273f1b926d8387a2180ee57c00667a15993977bd6838174bf46d85d14a1afa7bbd42d03c9e5f8e40ec82d330a76a3a741999c77db91401272df0b2a6eccabfa6905a31c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd02918127168c556f0beab50f38837d918e766c607a38ddfb2f34e1c897f8e2081d96d93b4a821e166e7f882f12eab995b0df2aae22625e102ca5c685d606f22ce8b45225bf6a12363fbcd6ebc4c49d2f136127651d9afb0e4417527a0ab8ecca1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he32f9aa15c03cbcf11639e85927a34c7613e15d478337c66d50016eb3f27c5644b74ccaec3ff712f46858f8c373e5feafef12404afd16d3e7d4f5c01839745e56b635da32c4b673d1ce708afc3af9b67dd49d3a7e7ea2503384e821501a837dcc8f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3da249d65dea4b9810c68e94e4db6ed45699aa8fe87541bc8166117e32cd56523e5cdb62bfa87b529901ce0f98875829b194397d0c606ac943a5d0ad92c2ce014c4ee21b35d116186a8bcdbb6f147792883c3ee83d44cb999baa99b942954d91c318;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8acf7d02999756b1714b067769b865a12fc34fb95f37901b30ee0be07c23a8949d4b96fc569cebfcb8f9c3e19969502e4d9a243181437cf0ad5f757929fb4f8b58789d3d8c5ef176b59ea0c76d48f8c44171c115abb5eec7e37486ff03e09b77fcc2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h195aaf4cf3746705705bf1576b7d9303e3ba5df36588202502f7593622cc05460e6290b01afd2b6c284754adca3640218b71c7738a949e8ee227c9721180b6d532b4d2137bb3660ef3ed491442391f4742655600523166f25ed81f84c658d97634a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ee8e8ab119be6693260d529faf68d186031f5847bfed1f7bab7abd66647e8ad0c6a229f0a42a75d38a3686ab9ababa0a606ff22755b4ce44e4424c71b0272bcb8b13d3c6f5b2f59c945bbec01c30ce470ba1868a73ef6ef1c69b7cea69ab9f6dfba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9a18a194844a6932b60a04df4350aba045c884bed2b1ba06489b545780c162c28b9cce1429aecb532e0484cd81582dacd4d6a694bb496cf553c5ad759164fc97ca46da47a1267085a6b7699894e332ce44ab03ab1b17e95fae7c8b41bf9d64bbcee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d5ad2d1aea4d04d8aa071a88e53952fbe868f076570dc831c7d6f916a67e0667ba280567453d1b1d0780f478ab6fc7cd2b6a33e015df2c7ba60b6a626cbdf42ab2fc87dc46c19914b3bea5e2c3325c091da4d9159dc38ce5ec3f3914a54e512a8dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd61f18deb4dc1eb908ca54b29470384db4ed6d8c4635b84a1a7a7d64d2af5dcfe4d8f8d45e64d3b9553cf4c72092279d0041fbe26f4836bf07b72649994c3dc51352187ac1b300f5239cc49f5a78eb05652e6b3050a8d4d1e9a47d9e2540745031e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b6a1e45952df25fff2ccb28fcfc4caa256eed00477cae38fcb9b7421798142a1ff57963b330354d505bbcbb9cdccc99d5f04263392c781511019f9b754d34aed14bf10da05554167d36591ce1ab823e19d3015f3e457ecd883bb52d7e6636ce6779;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb16156e6dfa0217931ed5c50b83d7d326e26f20c37b315e02d6c9812eef70654469cec05cff8c1b2520379fe82ef41e9cd4d4e85691df0e1e2fdff8b2a30a294da507d953088a4fb26c2074d270f88856ef1746f277c4698be4b9df95fa1b07d636;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc56be9fe2326ba1a7ec419e6be17938cc0c01d7fe2ee46c07df7aa2927286143ac63066c222a6aa271c74548b16c9c2035c5ab02b9df57576bcaab54881e22c91a6ac6d0d12fc14cfea1b253943c9b0fabc645b41b427d90907a4b6dc1c0f4433d9d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8c227026568b29c5822b0c409ec12f493a4c84e6e2ac6b67cb974f0523ed5d11b6a17c0f59da597123ce935898b3de96d409e80185c955afcfa1e57e4f9a94131553c749a7af9834311c47328c3fad775acd1246574282191a242fac95a5ae0718c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfa737efc00fa1d92249a58e5c940992758f4bd5bd9bbdff08a997983a093b4281ff41b1a63091e1ccb8d39738dfc3e337885fd65483a88da0a1d15a2fb500febf0e495499d409d344f4c71588af9c147ebb3a77398b3c21327b43ad3a293670ab3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h421626b5eeb85e9db4052d18411d4bbcb659624943aa72acba9b42dc3c0e59d8f607e14449a1fde7086d464567263e21c53a080163fd23d9b29194c2cf4516da17fb5dcb0a5a8942fa28df18a48895da5c7d31c0c88ab029b0fae705feea414bb981;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2acc3079db11fe3970accb64bcc19877832fbaa67a3d9bd5ed101bb50ec7213969556619d7e2c03593e970de2ecd430eace5550600947a17ec6b99ba8177e04fc91dae7eb7a9bfab866a35ee4b151410abdbc130553d857f9e08cddf6b61787a8835;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2c5bbd0629687b7522ba57c6723482dad5a2bbb609c70160be04863d16b2d6701971bf98fd5bc20acc24831240fda36693c64f113a1afa57df7666fab6f5b41018d35a7a6e802459f7023d8d7726950d92d6864cff71e567c4c1751e8d0cf9b724d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf90f3e6e57918662a1e8ca45d85d365f87e22baf5ba42517457eb9e67caa7fe8c66b7a13c540b6fcafa743da9739c052ef4f7c171ca2a7eb336dbe275ae81718d28fade3a04a9fe48896bef7d7b5bfcde42955d9377c8c8cccc66642ee4d97ccdd46;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b38ff04b64fd7a329aeda6c1b6fa417f5ea81a6cc2a18c6c1b0581e4155a4229c004aae1b2b2a074dde20e8c7907bc3eee87771ecf9957dec031878d42c34f4d644b4a6212d5722f9bc77d602b98b003b0cc2a0c3c370dd87dc91240c8f84070524;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6084bedcdcfcd65299a1186a9d90838d81d29489b12284f932e40aa179d5cdc750da0bce84b44d5c34265aa410e7aaa7858452f25c89fb4577685f5b4887cf8d4433126bff01230c49b0d8550028514c503a17f1a2d068c8f3becfc3a398a496dba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3702ee1e9af9b7e91bcf6e0096c9f88707a1597ba554d3d8c040870971a056f83c8fc273cf9ff3a93cc52f47942e2be1adf627b549aa854bc67851da737d50c723e86ebf8bd84a66eedc991ed125f6b9619de4e57e41acac3289b251094293eebff3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2189458ae8495f6e5dc4d0e4be0e07bb81f6ec2dc3227115a63e2cea886e79d68aaa68fe355499cceddcd35d9ababc206ad47f2bfb35dea1fe167e6955d8948dad193c457b857ae8a23812e9ba685195cffe58342431935c3b883fe86b6bd128c9d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b082cf38279cc21b9f56e75b82fa51087611f295d62ca2300b7dc7833c29735d90b793c1022899a2d6b8fcce88c68e3cffa8968da2f5a90a0f18e6bd37503ab8d8812e86d43b81f3faad6fa105cdf82d0f2b1330df477e781633dcd0a453e48dee7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74ecdaf43e007f8e5735920211847a4edd61cfc26a577da6d2d27ed0be48d52690dfd86b186e4cd264636c7e84aab21527fa95ed18e743dbab31c9e8eb21e5f10136e9c3ed028dd2611fff50b0177649f1785139e2f2f12a240ac725ce75d2b52d28;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2919f268e586d4d3cb21935271f3896da1338692bf0df675f585a2d5282be80ce35056a5ad9799d127932e05a33a61fbe7d2d25281211c3f970e645a79d1437aa220080633bdafa165c33208753f4bdcb7c46193f13d64dda11c8c085bd70b4d15f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d69f056c507701255f3c2b604c965c7c83c839a31a2acfd94c806b3649b6d2cb73f7d6b546594d29254d4b9e127a749f6a6abb9a0414aa42f6bdf71a4a3d86ebe2c718737e2cb8fe954c921b03f4545a8357fae82fb233ce568bfdbc44e1a120ca4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbf4a300e09e69e44509179bfeaeb4abde1f0681995efda4204a3a277611a8d2b17fc202dd079aa9ef878936de621d96a0210d9b92c9c62d522a1193f502392f90aeff50fe8cd1c018f51b41fa1c0ec19e508083bf193e10193a41a397a655452195;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcd212e188a4673ff7ca284f44243beb04f99bb8b6fa9ad142e4e4eae0764c6fdb09a7cbd76d7a900093685f405a1479c89816044423fac7c4c3eabdea0e82bf6a757b4eb31bbc7bb7fea1c5c4aedb4fa265310d5f6f1ba3c84fd2beddab64bb7d1b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f65a788f212a388552b72a339e39e649a81fbebba8777873809f0d8920f8b6d29c71c75dc8977adcbe3beb4258c579661fc706494d6d4b004d5552a3a38cf4fc5e95b5f32c6ae0cbe817dfd52da0ae93a823e611d264a0408bb3e2813645e1e976a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0ba37cbefffcefa91dcc9c4cb995c162332583c73d3f340847d8fbce20b3a2005285a7c3a9ee0f07349fbdffc1065d66751d1d39bdd60511442095cb8803ea682c7ef0c2182127d4defc20911331d94a001bfdd182eb465a60bd2a2d2b0290431ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48a281ef547a3afe1c070d8bb7016fb97525cd176080f312205f9b095724df6da2f8ffa57d3a25c31ae37bc1c5734414cce48f99caa617bf486be9734bb25a9073654d4ffc65b854e10062f7bc27d168b7ac2407b879cd82cc00c6a4b7e38d964a10;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h82704f4c2ae5ca6c7621c091444021fbb9e7013c5c7c0552953dd512e5dfc82f443f2f0a662b5ff5c45c09a1cd8f55f8dedfbe207218ad36c6acfda8599bc6ccd9946fb39b8584f55312b300abac2554b02c113248ca10c5f944211d1dbbf52c7f53;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66262105f0f589fac17791d88708498d7dedec6e10cd0a26d8f8b53a94b7ce90b914b1f3bfab9e8b9493505082c7172942783854e38a8d05219bd4138bc502d8d27e34da86c1ba8b3bd2ed0ad2317e5ceda4fd38f1444a37532ea8a2dce734044ae3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6e793e8c13c547378f7289a18d1b2dcd5cd054eae64c88caeef0e4ffaf59720d795eb68b2ad95f2cb07d5eba24f4e10406008570b36df9ee4e76bf5089096132f01d3d25fe5a7965445213ba8399980dde625dc58ee869d3f5547b79f7986b5bff6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd055924aa8716f1dc70f43995ca1ce090b3fbe9c1c9e59932d0d849fce8e6327ba750198a872c2d477abfed8f7e3f9b0be86e4a6f31d786acd19ff14c0d79f0d2b3af2333a6f38760684e92b44d8ec7759f4fae7a67e4e750b07924f52a68efe41b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h223f7ced5899f0c45a3e9e63b8a5686e5830f965b1503c97099924fb29ddaa1e8a47176ff79ab33907e6f71a9ad91729caf07e93307a4124aa643d461220ff68ac4c414e772f6ded33ef3590b24f3bf5d2b126a8fff999568396495c21b6df6e0006;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f8c6ee9d827a6324a752155bdc62bc43f87e17ab07a6f0d74636e319a0642894d84848417ae32e4ea4082b44658ef032aea1b2d8d645289c89f5dd215e811b6880237ea516d60fec84838bea5c04dfee82fc4452c126d582bcc2e47522d98e8904f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h691c5fe4cab302bf37a448cec39487562c5a93ffb7db9613c2d66ddc15a14399ae111e29c61d2ee792b5fb1efa35ee433baf187a74445cf686634cec8f8212dc54bef6adff0b9c58318af988cb6ff4c73ee06c212fef1a594b2a20abf7aa2263a577;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5f93a9c3f3f978fc69fdcf9018c8927cbaac278a957f24cb06c0e6df655daf95205fae4247768b6eb451b748d1a755696fc92c0813507b1aebe70a00839d4f744d56833ce5f679da098f9ce1750579ec820552ee8120c8792b104187e2d1a7a143a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd695215e9826074915d07158a73da93aee704018a2a77260046e1d9261a50589cc3cf7afd7c6f90a18c9e61edcd162ad788beafb60264fcace46c23279a74589bfe70f3d056641f6909cd4d7f1fe5e89c793c34c7081db0c22564d20b8b089cbc92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a8e4e20e4aaa1ffee4089528ab24412fb6bea75975a014702bb93611c44e61fc1703c41c481ccdd7aeb63d67f6dc76d76891111314baab20797a6015994930e2c73cc391d7efc16b65770acaad3dc1c7ed794d9a50d0b0663eaca4caec182c4fe34;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h638091ea356947f9a14281924812dda95c4e2e0542f91302ba8e6549c3264f606789010d8a6086730d7f392b2211b11c020a367efa5a9b8644b447804113dc5ed8270494463fe470493fd31dc088bbf02afc23d37be19abf4e66d69906a11119ba25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b47f2732f22562368103ec9e4f16c281394cda7c9403af784fb527793bb28827871809bfa805772d1ca4fe7b0e217583061ece34c738694c1be2d5ae3a68435e76055cf5f097df3b0622c85c26ed7893452b3badefb01e4ea3d14c77b47170273b0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haabd6c0e1719982b095ed9cc5f5c2fe2d2c1615f5179939242e4eb6cf116fcf835394cab099bc1bbea9293dab24cc22d07677dc64fd504a7d82ac80f8c489a36ab5b4a31dab9336379b88d65c3f9112f534b24feb5cdcfd47e3628c508ca10fe1129;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bfecae8f627072cb499a82abec91cdf0770fa02732b2de9ae1004e4838b97ec539c9b1b9c95651efca1952db2e5a369c0f397ba75529d1294fd57108076f005f2ef572f25f525ee6e94fda5951dc89f248f63d15409a717647c563cf76f3971aa7e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2571724393ffdf092a870660573678c1b0daeb0d959849ddb32412f701e5752bb5a02669981c390c181c8f64572ba86828b042800e91a456ea365aeb9c5797d2449068971e4721126d4e02be46d050db00f740edbf045280a8e620a8e9163f99421b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd71c5a5d9c75f1d6f03ac8467e483296712cff044a521096748a60f917454e2f36fc27b339cc06cff3ba034d47ae6adde7dcfdcfd9e6a7bea6573e3283b6e09928110e57b554d97f87d144381ffe2daa3a21d40e60aaa2a4c4d77ed37df08c70edf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha51aeacac3bea4b3765c5c7d97329669edd72e5fd3be86261d119ac1a32e8ffaa5932581c82c688894dd130bef41ecfad4d97664f873a5361d448e97fe3ed3027bdde42ac1861df19bc79031afd2867f4479b76b6b43b075ad3fb5b4672382ba9203;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6cb4c348397e87de92c8623c59a77a68151aac0b7df16f6b5d26157427710ec58def27dc47e2ab9b06907ca3c8cc1a25250b91ec02da58c5d957188c0a68be63fec82f9331b9ff98fcf7b88bd8c19bc650eb055485def785b12bc6c7592772a2861;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h670723f28396b27922e6386c3e0341c5a5822122a54b179851edf894f7ff8febafeba18bcaa60d4b50d20e688733e9236916e06bb7d4c83f3aeafadd6b084fb7ad832959f6e0e3ef574e726e4d113c5e0ad64d1d455df31d437b587821468df70312;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5be9bde0827103b9c9416f425b5fc352f1de552a328f668ad8549621ac313d1dcbb8d93b2d2a24ef94b007bf40cb18e8ad39a3efc2563c514b5a675567653246ea5fd5a8a5daf00965cd04938a99834f5b6bd1f5060580ba59f1096dae80a88399;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4520dfd0e54a49688a761755912560355a64ef4198f93bb328acab2602fd1612093f12c2b30a3b66c9e96bfc990183acf11324f2b6a26cc2e33c3e03fbd0a649dc72a4e7d191e7b18c26e802c56ce317951a0f47a0f4ded50995bb5213955558286;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bee35cb90fcdf6f5f351321899cbcd2847c67a0903e49246678e86194e3d9809e0231d7e3c0170658a0b5927347eb740e64a5511725ef9cb536586b84247574d14283f5174b5d78b02d2fdff5ef682a953032f954641259d9d33696f602db89311c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h580f8160874d2d6551ae1dc8b56443a9f77d57dca912299533a80e8fc5a8ca76423c3bed8a0128d349f66e9c83733d7d1451f1159e147ec5e6b31be2f34fd2a8a4e62ec9d23905260ae96840f4127b772543cab25d662e1a4facf017fc4e6a59490e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29d07d41b50ad5f97df76627d7cdb972105de8dd67fc0a0206f153bf284db6205a80bf5bf182dfc350e9b47e10f4e4f707d464dfc8a25f83098fc7f5cbf62901b900325cb6cc88ca6a81c6de8b17e78614d1503ac8837b4424b8e45dfca9cdf6932e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b1439205390c728dc715703dfa3dc6b89f82fa4b77efefdfbaeeda5c365bb75f8c0faaa994dd8a01dc930cfb9c83a669a23d65e11b408826a39709fa2252a41b908ecf17412aa4770c15fe63151463e9d4facbba292bda7675adfbd479f3c6af251;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0b2ec16815f121dd466400aa877b749359f826f28b980d7851d94488935fab525a29591a482d08dffcf3c3cc11f0f1dfa7d01b078372d659d1a5aa1b135eb76301d89c3e696b970ba7647aed646517ce8c35bd73c529d35c683ec7a1c8ca51fcc7f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h695d2318bc08277133e6bc43885335220aadb131bb985fccc712e4830991919eba66f86c9f88c2bc7c190aebb0e0131e4bb404ceecb36101f99971e1f9c3577a6e949c4e2fef18836538f85489b05ab7a1dce43a6ea8690fca0276304400b3b99628;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfcd230a4cb4fefcff094ee99ec7def02fdef98dee2ebcedb79ab6f153c527d41f8fb27fc92ced73ac235c6783a8c928936060b3cf18187e49860489fe8f4b4e52fc889b6105928908d41b139d935434326ff15120eb9b00b30f365ae922e6fcb81dd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfdc611997ff4977e438cdc492c4a98ac6348a26e84095ee581dd471d73743c1dca44255c3d9fa6457fd8faadaeb61161d9260c24c876f3b1b442468787284a91b15d3b09771ef963e6595d2b7f8042f1d9633fed62cb311c7d68d4a73e5f8aa071f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h126059e9b45f6c7cc09f897791733f4bef099ea2d48429b7c14ee19142c6dff7b50973592b1e87d32413807a275d241050f7ca7ba7d122db2364b373181cf9f79196a3bce34bf398ecf1cfad1b2be9c269b355eff4ba43df92ac0d2a6bda26345b8c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf786683d2dec2a4245e09d8407fbcf48145401726b5eb2db9c74836fdf34d43fcf744889f206f140ffd81ee1eff362a257aff10a452143ed4907902ec3ae5931a9ba62c640c81bf28af221e33cb699537edd555809bcec856335293d516b439af3c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50ea7c36ea5bde821d7b28e7a06bcc94c5355a84cf462a1694ab5676a5131c1971fca4de3c2249522751eb3766ebb595434aed29beb9d4dc604ed53c37c6be17a390a05ee0f601b1f5d3daac3c4ba1b13ab0847fc8fc816751ec912ae3f87e2194dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6981de58133a754418689399ecd638bb2005796ab59f622733eec46d0f4a8487b6f4e7d317367957084ae02e0f70545bf574e7c3d6ef81058ee5e2a0e9f9cfce9024a9d9a11d55975c89f820848c3665556c7280c702b58c1a05d352bdec4e07b162;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc5592ae718690649db01a55f10abc06a6f851baae81a48cf1a11bea65ecb1831cca4351e86e8ebcdcd51717090f5ff799460ad74e30481a8808d55cce6be92f800a59200d0b20fb4923beb290d484232ea0a1fa40227251307623feeb8fd75be29cd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h468bb5aa26c62b458aed90a63f8fb1c6a169e5e219882e3897f1f47bb96577d58deba943eebc2c4177af67dfe243a8adc60ea4af6fe3376287a384646f78daba203f7498472ad2c93ab1265a225f7215e953efa6be718718983cc49ae563b47bdaa0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5761afd5cb5fd9c42933e3e4277bfc117f9f97ea6a5279a999c036b554623e1cbf6a6a91dcd96f0eaeca5fa025bcf6a1af61d7ee2a9415a70da553dbebfd38b8da81a6c718f14722f7ff8288fe62f58a6ed54199ed55eb086f614246342a32ad71e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4378839ed8eb47da9c8a6009f72fa6db072338603754d590f5954d33416b102429e3c40f7ba973819796fa8345ae78559a0dfc6d44f851ea54686177e09d94a96c94131fec75c5cc7a8923494d34754601346c70ab2f14f2a36e5b99a6c89a06a3fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c3c33850e24d0b4e74abb7601a238be1ef0cfa8bdf18a95e0db5c68f2408d5fedc354ca458651e91fa7a42eb6af7dcc3661941a3229d96a7e7039d8b198f8fead19f46138fb8de34cb35cb668893348398da63f327109ad3839ad575d2330fa0209;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff1b332e7633a08a3132e94faf32483a5d694498a66a4820c5ea959cfe2fe20480a48d0574d86456d113d64829b2994852da0bc3fbd00945e328603d13ab60009f4f33e03938bfda1621904ab1641df567d0933a8d375d6dd212daf03986f17cced6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4fd9821d14d9259aeb5acb2b4938a83bccd12f6033ac10fbdcb40850b8877e18e0383c103b40816ecd70e250a8fb73553b3075dfb0edc11376e92de06537d4bd8f263ecb7b5dd15ddf179e27432898375e85cd7d7abf3757a423c68098db0154988;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cf2043e9d54a1d6b9a7c1a6a57f678c9460187755708048206d12bd565269f0fcad34c733c4ea166664ab84dea213678a5cf8e87e173386a4d9dc16ea8f13cbe4b2b928f18064ef011e3543f01c59cdb8ce93cbe762188d07b7fe057ea254e54175;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bf679e531638988fd3322a194b2c518b504180f45d434de26b6e085d0c157eff13f9ba103faffb9cc412a62949a28a6386788c2b01a98c7d27fe53a513517bdb9840926388add0c358254667382de3b5cedc5065bc56f6fb2c98de915ba97cd6ac1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd2e4612cbd8cee173f960df648e1e55e49f2b8653afd2d51caea19f16741ac8c28af999b1f6b7c00013dd377ca1dc75da74e8a35b20ad60c87811b03f57a00613fea292316b7e6d4f63faef4d07670f7c06c4410ec91668633ebd56f3279d598da4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba6624ced36d27121b524063bcf0f3b9bc4f40217f21ec0bbf046600aa4dcf5ab79aee6c6889d5655e8d1dcc2b7b7ccf5413fe280a49ba62ed877650a0795e65b3d395f691dbb04bf0d24dec3b4daa0fc8ba922237c7187ec13457c9a36bc642ec0e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h289c48aa468850e4db57342135e35be4c54e96158cf54e204d297cf6f1d11cd57695d44ce590a76ce70fde7b2b617bdb2c8876aa174d52c4cbabf1a7c361c414affe2f82968d292534e62312b4417437b940df644a39bd1aeb52ace20c602333bebd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ecbe4cf1339a921d9ebbfdc8d1bf85ad30bb778b4f34b01aa9ce49ee89e0216eebfd51d078f21557dea1406be1082a73b5c428813b4386bf24ccd915bfd2ee4ba140f6d2b8d3dde98ab3f90d552062369aa57df9b874c01729336997c8167a52faa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3c1a0ddb9e630e7c14b78b8857cf70fac6f864f7ce0e75f008ec6b23f7b486a2b01c231b266b133f4b64bb9acc99769bd4302f10c0c17ad63f8202e9ac972e85882e009e68fe0264bbbcaba888405147eec03823e3a50bafcab78322b5349975505;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h696ef4df87974ff30f7154f5d105c75b451004ecd9db4a61eec533dae6b8e5bd14f4d2e8e905aea9b1cb5c8f1ae5ff07aeff0c6601fa281e712c8e6cd6aa13d7b65079e19801c56b40e3ff0be35b3277ef0b695ea0ef411f25ea2ed32f5ee41871ba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99f635565e2f841d465e2a8ef26a7f4f1a7604abdf83ed62f55ae3454a3aa202bc8d6dd198dbcf0adf54f95c653dad878a5c60e79f7aafef11d5fe0bc4edfa9579716b4e4dac9a4e80f62b27e73e3e8493a01e9e5495271b0877fb9df7822957486e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb44c71b4f402b481140192fe1ded658c82f8ae0d7a595e677b96f7e68eb7fe530dffafa4c472536431a4486a1da792172b31112bdd90c6b4ff5f38c12443c142226ae33a7775813e5158b1ab5ef28b1101f52a1a7b0ccdc2ea6ef3dbd96898c9a08c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42a20ab032020cbfd98c6bf0b36029de043722467ea35bc6cc2927ec24a650a8ff29dd574fa00707c4aa78b9b38ff2c66e5d2df96a673f85413f450e328619206566f5ad6ca6b308ae494bf3abed90c377c44e23414d3ba029bf83d97185d4999569;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdba3e6890ebd158f0b39cc8c9f180c8d05f9aa3982c0e51d98376d878b97ae22700f8bc92c75400e54fb2a8010a0bf88b3eaa3f912ee9a1fba5f54963c2090c2fb8e95cc3f1ab70faa2c0ff2aba3b64bf930d8e5e247652aa2f729a92048566890e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb977e3749bb350cef446c997f7622e50f79c8b1d806c5c9c4d10648987f43f101ac9573df0c03b9daba8c89afd6a32f6be92565afb4cfbf2355bd5b2e140b4201a45ad2f814e34b78f535df1b5ec4546585eebd36c01a9aaff12b46c2680644b1a27;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h24ea778e2ce91b83036259258c7659f882169e893930236a315b7821538ab90fdf54850ba117402066ca830baee9369148c6e185bc6859c6867d1b1192525e464e8a00e41b4c38a7b3eefb4be00a0bcd7856729f9524de0a835ef406d57d98365a46;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5bcc9b35ea52c61a2da448606f91ab423e4be51b76b0e16f5d727756340b81ba359b060b0781245cb5750cafa44aec16a192c4a15cf52be617c20dd2c3c867954f832e587c6f90f795740e9f11bc15e4267056cbdfe16d39e1112d9a007cae7b9a05;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2076d59c0fe08f088b3d98d8b87f9d897ebca580abce538ced7a9df14ee4019438a65a32e440aee6f49f7f2dc5c50d9e870c1cba1ed35b37d379d605a2dd970c9e0dde2bba2b31cfac398db1917eb98264d1530770dba8b983d3257817ae1190fd3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4a2f86fb6d53677b77612d8570221affbc27c62ebeb906ce0895ee3bc122f0cb2d4a5cc8c14283fe7f958465cd00ce921f6b964d4317c658e68ffed2b101c30a89c3afa98b48bee71deef00b30945484bfbce7f1f11a48b75a244b79380741e1b0df;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89373afaf709a6b9d3f735c4478a744dedf91df5ba2a3bd2e6718145ea86ef20199e68b177c655fe1e1e918dd53f67c8b37633e3e324445fefbd519ede6dc24d063b546a71f4f7dd4050fd376148b5512a18a13c5f6fb18a3d491ea94f5097caef01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he42a88892a38f47bb25e36cc7ee8c250d6d2b07f69b6f366d4d9fc9acec9b6184fa741a293a2a9cab1f7fb5af1ba6e0c8c31f749a4aa770dbaa0d4d97e0b23fcb46c58751203cae36a847a43053dfd19e9cb0e0c594fb941692b9abd2b783061b524;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5ef7fe16627b36c603d24fa56222d5b578cd0072f2e533982bf570dd2c2bb4487d4575d33b3670a54d6bc51c8c64e3ec985d33cf875550c22380273bfa051b199242ef8ba86b2b6fed25dfb87ee09be31077e37f35ecf436a845b8d1328546647d4d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haaff4cc3ae366b217e1ba4497d521a517799148add0752dd69a4780fd7a3ca1b0ec8cfd183d8bcc0829e5665dea22735eb9071b8e3756376d674be62b4873c0f60882cd0d51cea4e2f3d6150fb2a7f9a5d1a35cdebc6b95352f74942d6689dceab7e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49d482e75abc392bd567db29f9e5541d9ba82586cf6972dd9a0a19335ab3ac3acb271afdc8acef586823b911bb4153082e8a08f9b86f2d912c70588b4bacff9c9b8eba90f7a41c1acac1a1cee9fab8e65511bc84a2687d779f443c80f002f3f2fcee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h78ba7aa81dbd951b1b6beeb9f2794c0e068dd3066c1fe0a0008d1b96fe9629ed2146ef51a789b5a25fc0c245e685c152cb6e9f248d250bc4eb98d885cf5c398dcc5a63ce3a49b666984d2a14f48b23766e66c1f98aec06295595bb6f44059575adfc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h62a6a239390801614fed8e1f86b191bdc7c5306b1e01b1099b67be144ea8408ea8451cfea068ec901108d3736c92210a14eb50986c0daaff602ba30e8b5144ad6412501c1f5d2a8ab604a7f29b9bc6e3a87e96e821bded78e51c0373dcec016286f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b2c0b159fd4bc2c985c26fcd040ca065376dded7dbad0e506ca9c3311a0210fd5b9529d8936ed912288b5482077c0f6ccb84be6397bfa683153617112ddf9fe23eddd680b969fdac66f0c14ee0bd7783aa193408cc7cb819ce53dd18b86a7be6a01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h853f27c54926fab0f11e7fde3cc8986a9a8f882e4e3bb0edc15d9f8066d0d5476c159d4bb76db9031502dcdf99db66500590fbc7934ceca86b02c0f08ac6531542d158de03652c361ecbad1348aee0e3a530775e46baa196bf98feb89dd1d37f5f9d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27e99b7529807acb52a88cece0d839caa8ebc0695d417074eb8b68aba361ac3b22a59947ea7a8975a57ce8285823c6454961184475daa3775fba3841f4ab5aae6dc391267762a93be9b68b6d5355c32c010d0e56d45a5a8009bf1d9cbae952073b2d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hed1048b7493738b41417506a76329f555a403bbbdb6f59655fc9068e4ed1790bbaa3b5721c3f84c3e41c071a3cee6710d08ee2f695769b198ecf5c078ff6f4a916c5f411ee3a4fed8f1ac98ce303e007ce67abeb1d60df24e93e9e52be607c20c290;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf22c76c7bdf78474b04dc62bc47dfda7b705b8bbd5e3d979c7a12df348bd1e3d53700cdeda44bb80d39013298d3954456ded12f2093834c3c24c0d67add79fd2c9a172f2bba89f47146ee65bbc19012702a7d4231231e864fcb0a37f07f113e89138;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8561528f786c2afc890bdaeb1f38bd968161885a38a0afff14838bf08e2658481a2ef19c724d9e9f116545aaf406955a107e3f19389fa05630f27d1f12f3b2d82b2060cabf842a3fe56750fa261f4d2bfd0abb64516f34df60c8ef39fac9cda513f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39a46cad7373d1c63d2b2f5f8d292243abb8872c869cb1fb464fdc40b6064bc475dd1bee7394f771e97d3248f7b1dc13672c94fb8b988806703df3ba96ca4930f975ffc147b5830de8aeadae9575fc5e6f9f794237eac4afa37d9a0db889b0ab21d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5807eff9341650d756e661397c80ae957cf309502efc781c933e5530896d023ff2ffcbac37c8cf1411d796a42c72fa6f1bf93da4fdf320f2f74eb448914b3d6653f2f3024449ca4d1231067941b3bbb28b12cc35e5555d174bb01f9fe22d9f6238a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h118e91ed6ac7e31af4482b262a8f8a2ea6422be190a689464b6f94f1da2c32c09a284da9477772a32225bd5328245e66c16139ff4fbb50c42b220706038f3af3b66b3a01e79211edba7ef481f5300e8f8df548161b405b61f7f9e3921c05087a561;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb877925bc10483a2f4c56b3f847c2442351e0a6afc459dc1b3277a5d14003be0acd0beef40b71fd2b78b1f70c1a8f92773a6b9b9cf3e45da88bd4896b17557702be6dcbdcfd5a1752c1ab04b39808dead236edd3c16e9ef238b336d67cd956269441;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ce039b95cd50739d311c343af1f16eea9109888a79b0db5e723ac1792518bc831f5d2d1841038c9a8722ccc3034f41976cd7a2e3b0abf5222609d2a1e6cc6175bc64616544b6d5c31a6d8618de9acc0151c66954d5409f68e12d785b4517c49295b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haee160327bd365cc1125a698243932079d92b2699cb3cf3239db2b22ca8726f88def5f7f8be3e152fa01352cfc2c06f5a677629a0819b3d0b8cf0857da58d013abcd9c341c135cc0f8b8e95ae9c34c4960815fe36bbc9fdf853827e9a10904254f70;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h202fd9e4f83803f57ca305912ad218e7fbe62665f8b2933dfb01c4c18e906c1532b9e76f3e4aa7b7afca2b5059a99629f7a9029e90633dd821385a63ce9cd4676540f324f59b5a6cf5cb159c6d8b9b71de90c9e608a6b8acc3e73261e94f82e35e5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d7d374702cf301f1e03cd3ceebcc76452a7e5cb31858b7de097cf55d8a9c249673eb87c025d255c8eebc332a18f913372ee5d94a99c746aba25ad49b5b4a4222e7fc1d8cc66bbc211b4fc36804005c33dcc98ee1f88ff4bd9c8291509f73b4a4134;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habd3dfa16c9ff19c9de517a0fc8b104c9e8dbf2afccfb8d26d1f94c1761e7d42593f1e03c039a9d4532acf26225cc1e883a1e3a58657289f366638a6fc192fa93a5ccb83e41bebcf7cf064d8cd40c10917cdeb30de363f85cf5b8ab19dae0a36fcba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba305d558256c664dc761f022ddee6e3f7cbd4a7bf714a04dc31ab56c4ca59c6540d610089d49d6370e4f1bd2477fe51446041ae5e7fd7c57c5e0ffdf4d34245495d80fc71e9309e036bf29eb0b771a3af4a1f766ed732ea584e3b5d9021173b65ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95b3a64bef6ca6a57ce62f09aa29ceb15c5d6cd9691011bdc14be14e0a78cba48908721fbab6bbcb9637b4a6694b4cb751c4efcae274a41b9f6d0984ee3ff30f6f73e8e8059638104fc03588d7c3cb187d883c548147818eec3d27fc7e25dedfd396;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h692fc7661432aa2d5e8083a50f258586944ac419b9e85c6e7ec14ca6dc92090c6acf3970e0535e6479b8c63cecead080b6429c0a8ebea4cb0ef3cf05c1e1878b11356bd0a711739a1ca8fa43b1dc4f28e6729fd9a09e445b00dcbd142a9638f6f966;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69211359ee2676b1ff4ce51f4e027d52e668ef86d1c7a9b484911915c3d294a180926a2d1bb14e2ccb0c5465a4f27ce6b927c13f01826688f618bc042fbf484d5db51b2ee6c1470e86a57db0a3ef017908edbbd662b08c6cde1677d8868e74e75491;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h999286671917ce08279ed013e8ddbc8a7a1c16b408b4f5a58b0546715c0fc55ab2f0e54cc6ce2fc6346186a2a5e0b88419251e6c1cc1994dc1ca477faaebf37fda8a47b6cf1c39fee4e8aa4c81757579638be65ca074330038c276a74d0583d44cb5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b197ab98fd1eba1ef89cbb525e326b06374d89dbbb313c3be25ff3e7bf4037886281dc9691f1dce357546fa5edd2605005673a9bb7571163a0ff73138718904d6bacd423970bb8110d50981d524ac39b66135062f1630347690f7789b2e4868e429;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd2f5cb1a39cfcdf47f2377abd97f81be2d6f23bb39f6c6e9d6a4fa5f5f5fbdd3344e05df1a5ba2810280de762936917623d827a8ff4e20cf3e9a8ecb1380e41791579dc68578e89bd1705903adb78ef6f9846e24ede064b89ba216040bf3887be85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e874b1a363917fb9db4f86ab0130315bf9244a942fb12c1d80ae829cb64aa62d2d4228a3de777aecd9dff2fcd18588cadf3ef6cef5f2b6fe618bf86ca740d9af2ddc8a78685e96d7805a214e986a49116a48b7f4064d628546258fd4e3ef4d70d30;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5fe66c24f8d91077349cb6e958361cc81283da8873fc55abc40be26d4714ec2677862791b506665c7ea606efbc224512853c638d7ff45efe29d09612bea656f1edbbd1ce37ed1ef4201194fc2db7a53a97931d9cb9b57ede8aaa48d71f881ed3d8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c66af74495db4a0db70586afcd19d512a178426647d94c066454233b9901d573a40bf3526142f22d29b2449d63ce40aa6707a6bc4b3f3fd42a453379ea8db0fa4af386ad49df8cb7f130b465fc29cc452787807681dab56fcc89c52037caa92f34c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a78d67390f880719796d3832f1dee8981bb20c46eb7fb618fa62cf1858a3855c4bdf468e9e04c790c564a5ccd549eae2b5b4691df3627b1ec7bd584735aaae6f098a22f6802a243700b65de724859fffc864c7580560e58261f6a520171502335d2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc19a9ee78c9b0ac9b17601fa60a3ddcc3ad26215f97942ea1e43879713f325c1ea1d0af5dff2f33a7e95d959e81fca8508c0da849a9377dda55e0598a46a7c608e29495188e27f39afc4a0dd459802ab6b879ccbf598744e6aba45be378a39297c9c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff7a69412206f9d9be6b8799153a1a8691b03ac33c7bdbecca39fbce6b16b43af8e44b3c685167ed6a8a2253ea9d78fca97ef7940827da33eafb7f7bf03424a9eeaa0967f813a13c5bd700b3247db69eb2589e896e4ec287eacacb1b762a1c9d458c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2d9abc2091cdb8f8f17d426c07b2329bce3c0ecf1eadde6ea44fdc26c93003234b9f9d7c3ad2eff40ffc6c7c7ee09e481e6d945c1b5707475fe0898ed7845fb5777ea7fd1c67af73119ae532f913a5e1c58ea10fe63e71eac21a1565ec6e09e0b642;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf637654bd416785ded5a9b8961ef81f3713dd2a799369eca41ab9a900b78192ee9fbec7c78d85971e717523bbcdbb6f5db69fd87bc734f151755b646cb90bdd0671157ecc6e157be78fdd2e5f76d398c81be302af3e64cd94dca8100823fb748b160;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8458b531f8edb0b7c8cad4344d0aed2be211ea9e3f869821a4113d637f68f7e3b9bef3ab0cf85ad3f5365f36ad9387bde0bfd27c0e470fcfe88c8174800078f6abbbf31d94ed8666d5aec70750f87a02e8daada000d803b71645f182a331a3563ac4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2072776211690939cb2e12d5ccc2a4897ee39e0d8ad8eb9537aa6873ea18d465591c2a4d4ed916c8c91f18cfc48e1e7b48b9451aeb2f4731cc5f8be47848c3a75cd568609de13bec4786898cccb0a1c15b36ef66828dea10c61c0d393fe9195793ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c9bb1023db62a1b404c89ac6cbc9ea9e95513d0a832b164206445a1e954e460db4d35822db6133bafcad2e6d2a9f1b600e5a00a199adc98bfb1a84f31fcf3c9326717595e953fffc0c70d48f7a7b87a83cbf2b7e2abacc661d2174ddb34a69a8cff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb76dd7c2a55d1bba97c7fcbb2edcdd207c222e9e3d937db14b0ada6271b9b3f5b9a99a813bd994dd039452a8ecc8677d54718029a8489a46a9bc6d6e31e89ff7a6404ed4c1d393489ed30de95405cc9787a3464ee9de2f8b84050c10a178c9e59204;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9a30e3a8abab8ab4b3345b35bfafdbb3a8cb6aff345ad45c2b07b2ae1c5e08b99bf5bb29b32d566a2500cadc7ac814714d8a4e091fa1b888e20c52a014f14036e69c4fc31ed64d72a845f0d6c02f196f11c0fe0a9c810c66f062357209ff2fd78da;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64253cdc1ff0a01c982bd07566e02c8bb0597c5580f7654ccdd55765cc8def8380bb359f34faf31df57d43ec7e06338a1d5f0f536606b35bcf348df64f389d775760ce0ed84c3440f4526ba25e1414506d25f1e2c23660faede217d3f944570155b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c37239ea68c9706158204143f0ab0ba12d8922bb2d770a08d1745d7af30c6777ae4d59ba697c1c8c3942ca36878412179a8399533f70237156b16223f25dd90e55e7ba926bdfdf26f88ec6e133f1936cf7e535d78b670f08d5e751776e33ec6fbf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc42e0963a31790829da0a0c78a118dd599c94e888c73f8db7bede014866ab8c0c8efd1563d37257792af76c42008a9375b668a0d292be388596fb15bb40e94dbae85e6bbcdf0929d9f67727fc56c0ead3cb19ffd50881e3a64fcf31912a68c8b005a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8904e3f85de8007edb62bd310f4dbf9cb008e0aed8a60ea893a76a780d5d57a7b6ccff73989f077f5c3ee966d079fbd625f6750cdee4b2e796d540ea0f9f0c85d824cdc26ef05ae44a37cc7ef43f6cf1c0ab04cbad27a55fdec3d2890b16bb82aa09;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d4c710b3d6b5e41df0e0ee90bf91e9063ff0b4bfa10de7f8e3a8aed4e967aff7bfe49346d036d9a89f6fe228b7aec3ca699f624b4308395aefe9da449eac7ffd8f3e170c15c5241b56b3f4eaa867159b6a368a465f8494fb96c7ce00152ebae9cac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8e54e9be7c6672a637245871be657b8bb9e3bcb1d8a8ad0d6738a7cda5b971867a2e9bde1c101b02a837aa298cdb34fb5dbb733d66a53166d1c29335b86f8a9bac225879f51c57bb6bf40db1a3316b905fed5d6a9f2c1934a87756372df86087732b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1708216e0770be33b14e18b18131fbccc0e0bf30f42c8f1a4b972a1de6cc27ada6f71d8a20f50d8a440127b6319a6848179d227594277ce40b73faa116e23ddd01270f4ed785be1836831ebb074cac1d72b56aedee1d96a49b0f928427012dda55ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb56189d011345288071ea987eb4b17b3fb728ded98e341b20fffd85d2db6d535fec9df7435f658807f162975570879bea046a82f8d72053ab085c2bd07382b18060d726e1ffca1eb87798c5af4655be5dd0610aea75d77ead7be725123bbb50504e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5409009892c765db4acf75ae14477dbe390d428745f4b9b56d36dfdd74860f6c834f63933b8be1fb6b0b6c2ccff5d2270e594c8a4ca433704c19ced6d9547098121dbd7f5a6181e8bc611c2c7ff561cc78ee801e07bb7095bcf39d27b2da19f0c5b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1adcae0514313880c886e9a9c77ecf37ff7469ad4802652169926f2c41c848e0ad88da289436f422d19fc646329d066d2e7b3d5d655c353eec660eb4b309b5ac1124220aef48f6ca410f2b9263b946e4b8e8158fabfa86f9679aa9a50f654d830669;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7a2584e932215d149be21af484d310ac8dfa397b3209bff985073dd605699e39fc35156d1ea56e25ee504edde3b3abe5b517f9f622f04e441d78156465e999a2b7ddf3ac4d300e48d0b2a7f7aad74a214524048bc8dfbd192196837caf022d0022e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2a78e41ffc937898db645b0681c509897c49a4cd71bebde0d8637ca95fcfc394868490c4b65f1c737141564056a2d4d8e58ee4a8e3ec33f8a371fd12f87e0877c12883447817fb77d1c209ef55d9e72cee1331c06f2c52f006f68cc0cbac2420084;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31c5182a5504ba719a951270c5962947bc97a3e34ab9a13900a639513b21c372d01ae395a7cbcc6f43286bd4b78f0ee90da7ca6769804cda0713089e76f101e767fde475587a702d2441109a86601a940e7af6967e491af5ebfcaf1b62a649ce20aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71c25dd67113a187425ef1459e5281dc268bbedb956607ab4140f04e79fb202d7812fe49b525c1259562831477ec574357d96f849a630d8cc57d8e18b645a5e82568ec443693cad896ac766afbcc082d9c89eb850c243306c3d025bd4af7efb65439;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha004a10541a86005b3f1208b10bbbae09206c8a5427d5ee844801c679f342349d242c21e9e02c7dc3a21cf276bda560ac92c7359d176984f27e9dd1721f0a4b8f9e674e83efd31377db111d5f49b54d1c8508b225382f41b04cb72f0f4ba832f8ef3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h729b0a8fc5d3ac009341bd7a7c9478d1ecf29bd5dbf2e62b8d9233c224d04935a527b6afa3f057b0fd7c610b0e8f3a3a42c6a5d87c155521e97357e35867f36f9a1ce748823a2a136f3b98c8b78ec5a9dac0d5d4dd25456d8944429426c3b16c37a0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d663b039b5f6c9d6a0809db83c35a6dffbf183f54a910f5fefeb35f6fde327cc2b41d990ca3ab97221d4e12346e58bca42aa698c9470ee62bb23c5182175e7d520d9db8acf8588d6f4aebe86ded86e9a4e837eeaab558d40ff376e2be16d1606544;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ce311a015b3497fd9b447cbe1196961dfc5c0c691e8256aa2785ec448d2d2a667a470d13fa2b31496c7925062ba9322d67738982ed4cbff2c7e2e709b59fdb0b71f608bbddce3d56e34c3f2becf2bcf838ed866f0f100c4c0edc3e1577199a43f84;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf45ac68cd9e104f76427fc19aef998a0875ba01e191481434e70f82e44a97e96d669c931ef0a87e7c32203086ff6ad13f30214aa007f2421554c098525104bf4fb710cc766cd0fb40ad22c5d330da5defd00b36b66e78e9f0b98a2e140fd4473e3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9d066d42e282cf3f46a5465b3406087cad49efe82a70aa3beb10cd0e23a4e1c82ac83abae5c449f1a27fc55f6063a9e90af36a8293e50e3b8bb60b34b175c5a4ce70c1d153806073aa733f119febf8778e80982da41397037e9a6668428121e75f2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha89db61593bd315ad1fc027b03086d33d15a129cdf71496bd7c0bfc02e96339e043b8ef8d9ac1a17d1ca8a17ff5a1696f954fc9d309263d8f40c1e16c250e39ba5e49a191ca178f3b0b33f138adc70c9ba70f9939c35872c9090796804451f0ff011;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc9ba5e7b3ac167799e2adf2797dc1fc04c7efb80a4e8a344ed5e0985f8d3e7fec39718c578ca6db3d98b406a4e480ae9868434515db2023bac2cff0d68eff7da483672633e1344aab88d03424c9671eea0560af3e4cf67fd1d3eb6d3e7b02f9ea7a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd51d07bac1f6a5878b524c92d7995704ae429780cfc2e2fd8cea67bbf2d856d1e52b02cbaff1a8b6568cba3bddf7d63e89d915fb4727e21a56e801b7ff212af2290472265d08c320c69f95a5dd0c5fc28e6a251519154a8566f48d0f7ede5864650;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55831640740babbf4f238d17468dace5e604869f9d0d8fe7ac6d2d8aa506f22ddc2cd3ec757b4b8dc2ed627f343ff4429f9899ad0f66ca9b349b11a6e33c5e3b0723b4cb860b9b666bca137ca4133ce1e79e6818c32a3c2527fe0ea380447caf9ef1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c44535e7acd4d7e70d88165ab9926bef61a0dde4bead304c2e49674e2c006abdc3d9b8159e39ca9293f1441dbd22b8a23c682f7dc06d77fec189278fc459e1c05567f9a1921d39c01a3672d086d8d6410f5441add673a1ef2862bc1ff5513832d52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0561750d4a7cc79f9d0ec5ab80932eed3fb9ca9a0a1ad5d853c414fd8a6d18f12509c01d6ff1557a3a5e28a52d6533908bc0c42bd602d339ed680d4d0e9431e754f7b5f364c26683e2dd81347b9c6723eabdb9004e0c9424dc5c7133e6fe569bfe4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4729d6a2c3319dcc920ab81de05dc738c5498142b63a30a4d1f197e052361a714f2ef489ee33302bfd4c7f2ed25a505ec9c100e573d6d1542e4d5f23c8e862f9d8abeb703039a0a4d9624868877574e872b22a3abdcc92b521a8f2a514225d30aabc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81e42076fca6a9e767187974b5a987001d0f73d12e9de63323de9285c97eecff3d603ac7ba16cefb55470c2b3e37f3a9fbaf36487cb143da3ce057aff48d534fce29699417ef753d4fbd4e3aab0e5bf92a6c92003e6d2554720f4afe538c5800449c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87df3dd4610f14bc625efbca5c4fe6b1e65fdf36643e38b057f9027609e617c0b76c75f06494fad28c10a0dd4b34f01cf613567cd4b1450b74495900e10e8f5329265aa3ee29db80a512765ac6e89b5fd28561513512118324e91387c6f4aac85b44;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h63e1d88f869b3ef31582a915f1e330381f508be5dff06cb54fd9a4710906fa0885631b35ee8172749d609e576dae00441d43b03a230cc15a2141cbf0e3d78335987a3fb5f23bb1d45bbbe69771975d0f06bf8d8b9259b5a6c76085fa15009d130503;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had879f9e27184d6310aebad72fd2a0eef8651d017b95f99ac2eacaf4e2ff5dcdbe19b548937a68cd0dc97f3f0f9cf76c79a9fb5900c6f3bd3b693c2abfca9a2cb0e5d2def805e067a9e45d60196a1070c88d21200040e2af7eb7fccdbfe7ba381a4c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hffea9b7bd098d25732d1121a9450c6a67be5e604a129659090284facc39b3c0247252fe342fc2631bef8cc443ff6686f4a00c8ce45e5c2ff9837c2352c96692a7d33e07e922dff8f85f235fabff397bb92cef7dc0b735b040193086d3d09c6346d33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bd509ff590d52c31a62220bf9c689d4d9ce62b601237a7e6921ccecb2d1a6576c5de2c3b20cae1ab58f171e4de91d62b09f24047cb46716ca830d92ef95320b2667d6dc1251be74999cbbdfa9a47264499e630b83706996440556632d6794d95511;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h48755322675efa816d0e718d49c5e848b0dba7b6c4dd8831a55212f1653fefa30f013febe083746ce661da7e8e38cc7619388f43baf8f8198385a855cd4706bd0de952c4f865b5e7826323069154a139de40eba27e71fa5b598844182c613b03035f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4901b69a7f19902c6466fb00742870afc9353c1eca1e8434e3f97f03762ba5bd7c265c5e12f4ca134ffa8ec4b11514cfb9b3a3946ca6e7627499da257b4d182633466eeac66591604efff4b2b5ae474f4cf835255578ea5ac6efaa20ef1ad22c48a3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf64c85db3380dd01a5f05914f97ab23bae60b5cf31374deee5201292d28afaf2537f045b2a1e9f2628ae6542bc9003d8ebe9567718aa0755cb3b677c1739d4feaa56bfdd00e269a8d69b1ae29382b888b619a7b78e1377ecc354e29728e7e509aca7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89640e319b7c1d9c5fe8288ddf0a4acf1bc56a5da0436c79380dc98123fa60f2a7a25cd8fed79ffbf521374cfecc5b404836571075e76c9d676d101b7088c3722c1b60d55eed3d70946f40e0e2887915edf63d2e94ffd0b4f7cf8db178a313170d48;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c8f7898d149dfa3f0689d8add8150e4451940b29cef13165e2710f655dd4d8a2133dc0bf1c8aabf397c496a364ee5c50c4291813a0877c958e85dc1627f2887fa4669728e7cdaf563f988a662c9175ded77a5febecbc3b417ae2cb6a95ecf940c0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bfbb0112ab044ca9695ca535f70ff7ebcff5dbc6a9e2fa100aa98a6aa4c2eb8134f76d2c16670a91501e03b5543ad62b45c4a99ff6ecb6e2f901c881df7e2b97aa2961977b40a34ad72cf688d77b5f3622a7e0363b45be563b68a164c0a6b8bcdc6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h98b501e13c53ef6b3d575e38f5a66f818e88e7936d4d6db51a0a1937e6ac341c442b0ca1fd6597564124d3e3285ce6e8bf395033b6440f2dabad275ad2d1b62f273154a196957ea772628cb883b0c356614cb56d47b78e59882dd63308e4de2056ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36d16a355ad1ea882a66b14a7ab17f4b1a98a44074e37729824246ea97f69c75d484eb8bd321d90953e006f47520f526f4709590eb7aece89b3ac752577d8032344ed66d3fdad25135f150126c9bbef1099d8a66e66c6da79e0d0fe3bd3555a2a356;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51a825cec990a81d3603447075e6e40c44bd71d7973344c82d15e3bde054ec54eafa1cb2461069d00ff7594638b6badc2c6c7cbcdb1bc1d02c2df62daf460c618a6c51ae4f4bf9888d826296ab60e94481711194bd19396746b6d8610bd70490bf99;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7aca09849233977d7b8a9e253e89ac97038fefb3d7c54f8e7693b420659d5fbb89d163c69d88f5ead573fd2559b026c30f8fba91a9f4fa1865ea91b132e5015a88ee9ece7c30b7ebdafdf896c3d419d98524b73e0a40cf0a55cf949acb00f2274752;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ead356fca6b0d08eb009d7c4ee9c3838ec57a8914b61d65001afbe4c0aa5d450821a1377be618d5f281075e2910fb920ac12b14de5602b1107502bb37ef8993f2ebbb3a105e97a5dadbcc73e05d0fa68728c18f9c3bf8666dc26daa51ea75c5599f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f86d805e879ca7944d0ddf64d0218c85cb542016199d3e8d408da121aff280249dc1360124a1157d46a37ddf4d4166f768692ee4ea81a8650bf6899369c71f297bf9f562b619f75c5869b8bf5ed796d2df47c7a95b89aebd3441b3321a1fcfb9d1b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4149ef84ee3c129eca4abfc7345d80b2b8271721c673015df7d3d538954f8ea87af345ff3367ef7fbee926f47c55525d89b68e68d1611b936d12bf99894f02a1a4d96e4521484fcd2c5aaf3d5900f40a16d70c6dd282e70563795c715b1707df973;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a1d638dae333364c25a73d22d4109a543563d54aabcdb69dcce9eea414b8c4dfc416e53b1096048af6e2523f3b361617c417f562238fb188595a45cc744d844f9497463d1859d35a2d4ba9e2ac89a45b1945ac2534496bdd7dccb005d40e3e38bec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb19df6388618d16139e7804368637d93ec7ba9696e22f75bc2d91059dac90116067043faf02f11576b5aa1d689851affbc7b9f4a039c25fd4ce552e8612cb0006ef0d2b709174628a4899ba3c10fb9c0c14a2abbbad3ac2fe30041398516fd48702;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa2beaa596280ff6f5f967aad7aa207e2b79ac1fbbd86d34193c328705c2e2e0528ed91e6ab4f000821cca1389d0a297e9b46198fbc95c964cbd353ca8c5cd5c22682dc0fb2546f7219cf4497ba6d15b61018abc7b829d205befad5e36287af0de3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4afa5cc17b32c61f89bd0861cac0267a94e396b75b56854293a8b9c7cd555f6b9757b6852b846bb9780b74b92e176d2af07606e8bc6963c280e93b3d5beaa97929e13cee57c5422b3b1580c5f33071765b926d7f0d0e1227c4c0f10aa7d78696881;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3679dfcb4e8b5986cba83491b3cbdf6e0089aa01ce8c271e3b092353c45d7ccea46a1fee4dab33195ec293b325fb27f96754548a00831e8712281e49071071d3eaf8cd290bb1a4fc4f4398e9ade1fd33c3e669a883be69ff3e4c1184c9285703af4a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee8ca888d10a9d80e3943555131905db84874adb244e4f171f89b353511d3b9eff4567b42a430be3370bf3b4ad6e3b0ae15429565a7c399cde79acb11efc64d3d98aaf5a0fbdb4759b1aea406cd0128477e1e0a3c5d11d46eb24d0a91ea5221860d6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd98dd01216e0a6c92fb2c2bd4fb40d855517a938994bd5e7b4276d905e7a0c8827849fb1553750992a5d8a4cd14e21ba919ed419d1dadf51be268e4989536fd3475e2d61c14bee70211337721ccdddf24e219808e4a4693aec168403413b554bb768;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b4ac172794b4170a869c3101535bed6c1ef8e4dcc0898124b5e344823d8fb862f394c502f2f2e2ea25f8d18b18122ed5c3b10ec4bf64661087b8fe0646b90349165b6cf855a9f8a6814c50f0847ce11b6d13737fc747b906535400ca508ae86d62d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f2c8d6b0193b656e1510cc3d527c6c658d53cc85ffd0e97fcf27b60c699c51355f0b95ca4b0023e56421faaf9a9fa2bac4339fbf19f8502599f3ead813e124b4d0e3b1b9fd0b808d3c40605483d5569a5e7cdd2926f74e97e3104671300eded2a4d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h614e92eba63180b2b50321defb67f224f619870d1d1321a977ea569a60898a787f3eef9e5c41c5c1fc83d1690a966ce5eb22d84bf1c629bc8e71ab6e67c10924ac1a1d417a43c14d00fca261f002a4425d8d255e4757d9c2d050fce93d541a224650;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfdb3200b6550b7cc2540cb45159e8884f7e5c9410028d686ac02358d1310e40dcba0aa2098681b139be3d00d3a0a3566c42d6eaf75bbc44a067a979c2fceaab7a75e4dcc85bd351eb1bc5ed20880d839bb71cd1c751742f55bd57a4a8db91958b820;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8409e4220e7cbae01c21ba22491fd98b5c800cb23fe7bc970fed459cebe5e530b0a6f484073d2fe4ce897d045fe653b1b0eec5b5937a9c0a712cbd49a2a4b1eee7cfd1aaa95345e9b80cf9bf673b8f36e10bc42b23e493b19611fec6972455fa10f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58e845cb9c489430b7f83cc5b59ad0c764ce67bf85de34d849faeef7503a31616a837cedb655b6ab650d39507e581a90b5ebaed64a2f643fb4cb6afcc3d88866c7cc51a0989a0d6e821dd332e9bf9f0b2e66fa5054657d07053527fda55220789463;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha130d84321bb15e36ab0cc7cd252c23f8c22e3bcfa04d743ed68c7f557dd48d097b497aef59fed0f8a43af03982001514a760379b47fbbf357d4ca9d7913ca17de8b63109cd62b3670a26290e86a79858dabee8c7e99eedb50311355d1430b4c9d6e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe1aae53837c342f024c35637be2506d94a2a8cb27c51c0c4f349bcfa591bd863555f275e8233f101caa303fdc27cb4c8fd335bec2e2b7f9b8ac8435749be59eea2eac37d86cc05a958a3859511eb93f88a906d44ea285ad350384d4a18cfdc2f118;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2d57a1b062652a1c50c56e9bdcd4f7ebba84c9df31cd3c7879142f35bc7a3ff50b025ff21fa3b1fe7567651d859912366bfb81b527a8df81f4499cb793650f4b00d9262f8fea411aa33688af3fdabf8c9a3c52b85b2ae18e209d95944e0ae216f54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbc6b7146d538d21dedfe2ef2c028ef44e51e3b3036680fc787b7254e98dc8aaedaef2c99e9505c03d844bfe3c22f995fc69ca44ba648acad6f06dec75bce752cabf3dc59347b003f8046fdf4dc7887c1d50108b57d2c861f380a07a3d1e65a96ffa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h710e0fee8020031d8fc8a23dbe34d84a088e45ebffa15a640db3ba78eb1a059593f115fe8ccfe5164b7e5e2091d622b3227a00817e277da00fdd5cac3439a60794618568d7c47c83b8ddb1a66dfe5f2241eff4bcc3f37a797cc8aacd396352430fad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefe7193fa6eccc5fccf0dc7c37f92b9d33b44752c48971012ffec126bfb0ab80811e9d420c3919bb8181092fdb29947a0a541351539164beaf540249dca02aaae4123471df628c540d9743568ed8ef5b089a5cf68be2547b386297553684dec0016b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd44a50b828a145e11f5759ae737020a37b13654dd33ef8cacff634fedb085cf5af7037d8519d4c621ad1b4c3d9ce99845d90d0ec6ad14ce671ca0ea27d01d4a5381bc2cb2d6199fe601ae35f12c7ceeb0a3cb561406ddc55f75de89ba62db58f8209;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57c3594ede881bdd48ac117fd052c9ce474c332037538bffe8a1a29ac4c278d4de6d3c3fac5b5a558f6f5fe9b75d517b430c526c77112287a02f789ddabea9ecc69062caa3cebf617891bcd02ba4b181a8409af9f57f3516ce3582e17a62e6950a6d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88139239d158d53a73a9ca325cc6a4171fce87ee365b74bc26f13404efb59bbecb33a7dedcf19ae74e51133b7db66941392f54a82b380af47826ece8c7e003788096f09127361ccd30012946330bf4fd91cfe0ba7257c66b72afb43e732325e1bba9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdbfdeeb8efde419ebf61d47b22493ecf6721fcf6dcf93a688ea5a49e1f475d2d50082596dbf6f82254b0f6ece2f3a64597f6458095a73b094c1b061ddda1dbf7bde239e291db9eaaee6558189f1bcd692ac0ba9a62965d76802863b63309e2b5e76;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60f971b53eb5c133ccbb813f3c27ed883c8a15ae7577d4131e2481f1e49f44dd89541eefd95e2f4fbe771a22553d164a1d8d9fff884a162c031471c4a4b2cae74f503e211a7bb90d2a43935aba8aeb120f20340b81407cdc6ac1405ec8f090a8876e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h88c451a2a44d5e23df13d048f7a714485f9438db3035d109bb5a8018f80455bde518cc2c0e64aa50a93ff27df954bac14e05fa7525dec65db0e6d53870b605546a29915adb1851e5e7345a2aa7a2755584f4b00aa8ea07ff3f6f878644ee45820c7e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1814532b494bfdd8826bed5188a4c77a5e9bf290e2a294697474616be4c8783b221fe0134d4843ea6b2b48f4b92d857a3e04d046ae24471c2d34c6945cc0867f0430cc30f4f4fb34196ce07005d6ce8109875e33bdc61130b273038c5f49bc1d26ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1882adb4421073000b0bfd8c558790a9368f37e546893fe82edc6995c2e70caaf0a205c331c2eb0b743cefd773f6de2b39af5c5bacef5c4e0daad60f8cf47aa077c22b040d0cd703a101e0a6c8283fe09cbc142d7b8539af3abffeda6a66ccee4061;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he4be55007b290a7217c5ac34c58f4b61613bde57d34fe21c91b9d199e438090bdc3010cd63e763ffef9b419c2e1cfc7007db2115a2327114f17568e9d8825440daa666964606d9594f0ac158e123f35d671d0c1196b7c1f215926714110ea86b8d3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he88c08a827d49f3adfe24ba8512ccf8c4c5d7a23bdc1f0b403f396bf54eff4f5423a68a22679027f25fa760dc33bacc6b8917413b56016f3e7378739c71f101f2106d82f8db06b4f4007514db0ddefdae510f8b9eb18af0f6fa606626b86a2b55c22;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76d2a01e01f813e5f16e1a67fa2bc2d7fd4e97bdc3fa7e13b8144e80d18678cedebd889176611af506690406bfda849aeefee7a5a9ef1be9afa2b31c5a85789587069d9823addf1d91c16735ac97917f36c330f258dd90c439d8f2e6867d8e54dcfb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha66e7373b12a8dd0e592fd4dbeedb5dc77cfc7116a4219a8f5f640d929bba7e76ee5744513c999f51077f762459dd6d57ba85fab6962aac3f72b6287ddd09a1b4ab795da372a4b6b9ece9eae830cf8d1109293f3e024fcf7646d7c7da9240497bb82;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d95dbf0c816a71f74fb9e4b62ec2ead6cdedba206b1cbbabfacb5576887f9b96e170c407135b9cbb42ae358294832eae2f1eb48bf97265a5e26d26d927de120a8505ca40f5e7a00b0cbaf523f358344b162da5656e9c22dfa0e0ef2fa972e5e579a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43d950e3b2af61c5e69d4997f9aafa256ddcd25a66773fe992d1a09eee8ffa1791f52651211ef92a619cbc0c0e974f4072f3feeb888ae1c105d0ac911324045be9afef660dc9a0521f3bc512bada4210906b12553eb601edd2aad8d6472dc0f4857b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb927102aacf8260ee52c27b8ca9987fbb3c01dc30bd382d45202cd63ca093d44c4e6d9e2cafa8cae604672c6787ffa7cf8c34804e97fd604a048215ea8e03199f4d7d983598b574baac93636c799d7938e7578be70bc8abf2759a9d7bd8c910db60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he301a1ce8ba187e926c28a33dd76dd5371560e1da81168254ce7d8653b2145791e7e1efa5cce6a6ea746697c5a1b3afc8c0298b6fa767520c96cee898828b521c4b4db2db1430bef6a5554ef339e2b0eb92c5947e128c2c724937da0e6528a624bc6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4dbbe05038e7ae021011c155a2cbb9a6589c28dd173b8670c10a1c356e201088ad8e1002eb869e4e44ad97bc3b8271ac048f61b72d298296f95f8a404e2cd317e615f0a7f12fc617bf501bb870d495b6d0d5c6de572068783befad381ec3d93a77c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb09384253eae9b0f12f98fb88f3402af7c6154235887bf754949a43dbc50488f78695f30bef514bd378902f00918ef9a808e49d2caa9366ad295afa77a6d3526fcefb41e855f428d7c3f59d071ebccda28afdef564b69c32f64bdaee35206735d15b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c481b634e63bb4f73a9776c16d8c6619434386a9c772d75f04d7932924ef338d486f6c84c7e88246824b31884d7af2b373e9849fd913b62ca7ef993a189780b5e03062206db0c3812e9660821de8a19b949f240dac3e7036437794d05cc5ab9ee9f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c50b00f6b9d147462021cce93c0ffe0631791662dba526edb4af4bfc1cb7a3d46f5563c37114834cc2f3e27f8d9aa0c1be3915b200f20ff737e2841c7cca1281d5cd764929b8acdc68b02c8c5a5d11fcf638d82c69c523d023ef6636cab46b5f94e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29e585ab29ab28fc6314500f2d257c3eb34f03902f3f76ec07f35a89dd996d8639334f8a3a1cd1d4f78d0a51073e8c3c9079a9e1b348b0ca213111f2dbe4852db17ceeca70d7e4606cb908a4593b8034742ea325440bd647e9a68e5b81a39ad53435;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf72ffe44448fc07979b00b3b592893dea6a154e9ee82cfa9eb2f033e629a20c19c6ca7b434abcdb4f1e983d445c9e887984cc2acc93c3ec2634d9c3f57a4545f7536423b70c5d45b6dc4372bbbf75710daf8d82c7a94ab2a01688f98d48736b78978;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99adc24122000ed14d22cc6b2ab9c5445ade5b7104c81a8beb90b057217af6c91fa89e3e0e1eb759e263a7eb3b4b2571a80927443bbf51ea3636cf093d7e6b0bfc357bf7d946c25bc4161e703e0fdfbce691720a82c1722991b3c03321fc1f4d7d68;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2757d90ed6e7455d6b7ef0d53250bc8b10493cf350beb894cd46be6b5646a95a1349e28d5ebc443ace39f8389bb8757c259e84e502dea11749e7854196a07d94d0f8bd2996cb1853cb7d780f47a0d83572e6206321501db7b5069455aaa966e2a78e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h700bff73adab845719574a4b8caac8cbf9ecd0f2e55b1fc255740a42859e0313c044c6d90114ca98d9c7cd43a5396bc28e250c7bd7e6c871737e19c450b419f8553ec1582d2d4fb344dfdc824a2cf1f62e8b17ad3ccdefbe496fef7d11860c88e200;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0e12e1fb8baec94400af6f322174df95b07213975a605a8004e05b1880a82940726d9bf9c7df229d1a1d1eeb28ec7e797ca16e03462d292c08fbd0c39e8d26b479bae23db6452edd52957b0d9ec18748bd9fb25011ee463b75c0b4538e4d676a75f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1bb1c8a9f781b1ff3d4019c1a5fc72d6d80c7ea57fe2931ae659c86454170fb064ac7b6e4fde8b7ff31b635a2a4ac0e1338272ddacef574bc012eae72304100de72a80599008a746cfc9d47251902a4e5b0c67482f699cf2438942d178aa88756755;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h338bdec88cd1b16955c0808f1ac8fd4ea5af86eba5eebe26446531c516fd6c2cf6162f6f760ea3941087d6a4f540c1f759e1cdc0a84fc6dd908fcc3631bffe511001fed7f6128403dc808694d1e7e21935e6ca4eba4b29b2f97a09bef807f8ac7509;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac8ee4583b332ef94992e36b6374ee9c7a19f4f6ff1ec9481cc9a99d938b720a49133b2cc53146ea338f45450f9f750ddfe0fa2554ad82ce28d153a608c3ad5cf6f11173770a86d1507bcce243fe7266ca1caf3d8635e46c2b1c182045c9763667c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ea77b96411617161fa384c18ad37aaebee86171ea795a9a02c3915a035e7b94716b5c64bffbe08733fa167e9a18c1f300da399bb8a26fed9302c7a8a65c806685bc42531b5d8ac515de8102c2708396d588160c081ea396a0a6c566850064268372;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heebb4681de53dd616c3ea9df44c5c4e3a6811233ef070621a8eeadcab32e76be66ce1712e9178eedf564d5463c57b922bff961d8b6467993bd98d25dbd55d7ac2f771d55d7ded5b17cb29e138d3648020f0aa247b1e212bddfe1b53f0774751c431a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83bfa3ae59805aafabb12b4589b1c2e29387a9db9b0a162cbcbda136c1498f6103985c480819d749cd689d569b60ecf7c5a75570ceb46943e74db36e7d8c1f9dc706a464dc5a2d1a11878d6a3c9a0daaeb7edc5e8cd6bab31c7a0f34def588f6b772;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h45ca6941d1ef9c87217fe4460d1eb8b0559a58e72fcfbd6b4bdf07ecfe3a32cc2b07a73d42f3b1695c9464d04b09f8bd8c421913ef705e492661a35f4860235c8fbd756a03c571ed5316a5d920344ac942411d56b1e08cf813f9083dbe78813e7e54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h293a6e300c75ca22481d02ecc5c76c8293cf3a32cb7311c2a7c2418d722551e1a8a9196fe858fe3b1760229c96b72ac4a5d772c162117af4ac01789408c871a0214c92f6a05f203466e759f26bf4d1b3f161610ff38151e26b060ef8672eb4c907fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd69d544e34c5293933369c0c6029682aec36f30a7411805b32de65299a07acb9c599d0017befca436d9c2ab9bf410cc46e6f102b74363f16fd63108c877b9c906f28f8757768cba352076899b5ecc6946c3724b6933f4317bdff507b483e66643f15;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h268f5d0c7e04538a445e7d79fb56f81383d94a4779aa46de3809c9f765ff2d461c6eb9c26061ff9b65571af87fdcd350559a4eb7f7444307bfcdbae3b603ecf0a18756c261c02a9972e1962b3c4bba4d524a94f8ca5273930c6f098d5754798c157d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1c3b576cd2d34036b83e503918bdee3cf2c79c0fae7cd00f13c5d4a9b89c3e1498a8218ed11cabd1aa70cb2d9e9386929b1dfd4d506158dfac3af5c705a524f8cdad3733e62195fd3b2c3f5056c5b1a79252ebbf87c6879ad968b9f7a9aaed0f044;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e874cb8d66c8d93d6b5032b5e5d4efb0a3cd088e74c47715f297c14aafd85f5bba8e9007c95ca88df015dc4defd5cf10e68718c1834ae960e2c957010523a1cffaf993dde439bbd08a88d7a6b2af18cdb412ce21938e834e431096b1e1802b38694;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ac4234018dd5d7908a826474d809102fa3eb96f020f7f56f4d9b4130416f7a5b6010731919843e45201b4da79ac12d33c37391de31900eaf530ef6763aa7b1b2113caa00ab9c79545746b6aafe9ff46054d3399f613b5ce36aa8935cf3176b3d06c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h81872e97f4d7b53c6390ba509db8e4d909710b19181e52effd51c16d0f8f949e8cd833c599e003153ca04513c56e6d9bdf0ad825368d10fdbbe9f86e90ab185bb63b770762802b2bf15bb3d51ac706230d7fe15ba47cb9bfa3786740dbc6aa6f5a22;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h587a6e63a4efe6e0b8bd834ba2961ee8425d0b368aad73229dd29a785f90e076a52bc9d94fc68a11c47e897ead32df56058ba45938d1d272866b6d41778e5ecd76c92735a5c4e398c8a1ef08474adf68d9b4e7e8e792fcdd87b96868b93c6212c5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49be306f526124e68557203ab4c6c75b80b1242dbf884a6695c965f581c14764a49ed76aea3c60effebf69c89e710d94042aca8d349cd32b76b39a28d0d7f7a073a58634d61f2e72823f082015ad823c0bfd8299e2a3d2e28b5d1a3c1647bcc97ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e616b38fe5b609bd5c3c53b2013a94286992c316fbb6a59beaa0e3f3dc7361d878f18f1e460e0b704a676c1fa633e1899399767658dc89a6f12de7968737cc6480fffae30328947fc3ccdf1aa417eb80ced335c380924ab0079302b2c9133413cc8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9987332b39e3725c07053d908b2ffbd043575ce905ef0492da97f32a98ac7d773bee87365af7e0807e79af03eb49c9374ea05a0a4aaf7feb151001095480b24a49735fa7ca082c1fffe78bcbd2885aa406cfa09b117b753cb17f40f26ef3343a14a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h651acfccea480e1b4b90513f623bbb42ca52874687df46f5cbde5f0dfb4166bf04908d16e2e9db21a652336e75827e3cf48a829ae54b2d57eb87ad7d9ba3f784e04f8184126ba193d0d17644a2be0184f6ac15a4c8071f854cb3928e28c7a0b9b563;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca9d2e608ea09a8a6196f2032bec74681a8ed9adb146c0ea746590b214568c31363666435a6079981ea529623866b6ea9448861286eb024b68627a8d8b11e835403f86a995ac8806e24054b33638b2e53050c0c3ccdef017cedbb09f5d99d0212f62;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2285331134d7f40e744eb7c9f7a439d7c35289273c33250ebf436ff90773b9c49219a78397721d124e059c20e41aa922f62aea6c228593d400dd7a9a375f079f11386e44ff3c816104a72f3e4654cd2e9326004df3c0e4abec2e2c27bc4a9e7dbdf9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e687e303c976db64d907fbb8b19d7b5a1d0f26f9f793c8f6aedc2c172d5057b2727998419074505b5555b62528f39eaaa0afc6b38739631027232addea36ef7f27d12bca8305a7f24363e0a2fa0add1e8faacdfd983e621bc288d3d4cdb0171a6f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1706a782be73ec0ee07aca3b35d7d5e6e1f18bb24911fc429f7e1a30ad7e62524c6a1239f8e34c025ccc3fe26a9ef6053fa073904bfd001ece4f69d0a3db946eab895351b34720490b8a113dc1cbcaadf5511c5ff4370eced32671226785dc2bcb1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89365e3dd454921b25450391542bb6b2e44c7f35e8ad4410a5a87a91100ed2e245783fe0260d287fbe4b2be7a14055906af285ecf47416323a53d6817fd2a6b2dab72d2d5102eb363be4d8cc02e1f070a1d49b2b5ba6f9abdb592d73a63cc218b0d6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55a4c2fb0dc75fe6570ce6e0cd37c4adeb7d094a8d74dca1b6f328a80a94bc8a39dd9371c10028d81b27e2fae472323444420561c1ecad8b9e37f2fdfddf36374b216fe61daf7ee5422387dbd238226e0dbf60543c765d25bd73a406b9f78e38226b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91f1334324a71f4e0c66eea79f70a60eb20e87b938a1def1648053d10a2c163f2478cd9be164c6a2028e7f7fd9d1f0003b708a2f7a931ffa5ae8b2838b54eb8d56010f80b683ac87be00b3160073434fcbe63e632bf644f4e8d355cb0d232a2bcfd2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4da16de21f46f4fa9c226951c62187edce2ea131a26495e684e7bea184599efb136cb1f024d98cda4a021f237d0950c5ad11dca645e5d16a0cfccac3387d97d85daa4f52b18b0564f1efe4d8626e64f916abfc17bc96d09baf506f828ad63349e671;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5f97df118438b41fca5bb5a2e1de88f56da5198d464cb19ed4b8abef9ee366829f882d9e7dbc91ff5974f462a5d463c177cda9b8186c8ea5c652b267348573c83dd19ace798e950ed586b92719a0294ec0e0e5a12cb5f2bd7c3418477b23c034aa2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc201cdde600ba162c2ad4c2447009a098594718621e0f28deab9718b2d14ad7d7bce37325ecc866379d5587fe6ba57f3b136d9d1a182abaf86d959c777240b486d3e93b8b18c540d16c6b96d7238581288c9ccbbfebf064c31375095a762d6f288c4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h687c0d38d99d48a320b18a969684c17baa37ee6682952505e3eba1878406c037c780a4e551d5084485d9711dd51bf31f2ba5e41f01aca4eeea0e6c14741e140c832cb24e325ecc0b95cc674b2dad93a8ce947aee37634a9acbea32dbc3df358df8ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52917ff6f4d4f5fbdd151865ff35815504ea1a7bb5f670b83421d8ccf08b21d13c4c5de4660520216baf24428c983382a4a5aa14c16567e2dae65af6cc7142e7b3f5b2774832846d34b437be9a2c4fbcd44ab237907c505aa824531dbdcb90425a6d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf71d380c06c5f64d3fbf7db24e91ea3ef58bee2942cdc0f26224478066da2162768390b65a51f5914259d3239bfcf3ce14f43f28c4d157e498959535782ce97097db125d2cdfb02a474f332254d8b3af32b42f564e696719655106cdfe58b11a1d97;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h419ae69c22e32e0e9bcdc546499a8a9da8ccde25146376ff63c7771b9c5f9230b85cbc9199ae8bfc6238148c49ca7fe12547534a485aa4c01cda3fdde78b442d095a9aeed0309fb656e95dfea87de461a3e7097ad2c9e0bac1b3ab3dec8eeb0e957f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h33a45fda0fe5c49308880bd39279d6bfbcec29f4b7bd34ff149bc02fe9d0e75927b1e7c56b1a63e91917609b6538d41376f4f686b2ae0c2256ef1ebd943ccf9aec6ae2df6f06ec6a0665468ba04979ab8f76116cfbd922451432eea36a432412075;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5828cdc12eef93eedf67b9f9d5a98a22a3aefcfd9bb6b4d79866cfae376a91375bf6caec37530a547285cd32afcfcc32a53c797edefbe2bcbce20468884b1074f65a406c30e0dbd69736dea0214a7ea0d90bb35524e987f4f8e556aabfcc1d66c54e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h930aae6fedfcb54bed30bdaa599198b2c2e545f74a591c0ebc344513de8c2e8001ee0dcd82826eec347800db1fe52e0ba84a8d910af9c15273685de966e2e18f269919fd08ee8b9c719641186d74beff78776390c795eab7a7ec1cb3428472d359d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e4eb5c78eb5f77b7c738f5b183939a5cc7309df567d375c5cb1141ba09f68db43a90aeaf6f6ed841c96684c38f03b727e1ab57b4d893c7e4c5cb5185dec6ba19b28b2fc13d9dfc06f18440d97918c286d199a86b5639aeb37ecd5e282dd2a589c19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b2d82f8444ca6479170e00d47c20b4b49113fb07d10ef8fe8c6f2e53073595278600ba078dd7df571515cf28c03cd5ab2595e21a927af03f88038a6a8e1aade7752a3ac9f5d623f8b76f17a5ab763fd4235ed84071468af945932d63ca0fa43f4c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfab569955745407cd2d4519b28a294fa51c77e69771c5339195675e20700873a98d7e7670867af04067ea927c2bbcfe043641e716a0d6d67ee29c73b46defbf0cfcbe813e426ed3f11ece58ab8d30b2af53fc6add4cb630b14ba12d6412cd38ef7a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc94e82c482d442bc67ee7fbf0e4b873a44bc011fbf61e1e45b32c04e964bcfdae5f9a6081ad4d7ebeb2a07a988f4dfb1a9c2381d1eca53d3bcf822fb23025eb7290896215f9aea823407bcc1ba682a686e1fb9b0aae331db25cc800c52bbbd5bd5c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e1ea50f50b79aaaf84e8a23adbe6ded2a7e10b75e17436bd579a4dd02554db71ba759e3a7cfccbe0be00dc4fbf9a5d076264d19db4bf53d69c16a6fe2a840276e1611723781af1240eb76ce084cc791f8a7581c25e77efd49d7f2f74f2d83402488;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he98a4d2537be8960425b147c8bc38a1bb327d10397ea9f3adcfba2c7c4a089a230d03c857133b6f3f3936aa0776d11843eb843ac18283be11ba86091fa6d4211a8f6e9cf28c781d347492ed2fc99071445488990ec6d7d0b4b4717099334ea78a236;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc8df59ec3dd792d3c05bf1c020d5c95d4a8b37fa7fea549f1eaab4c1a10158e056379365eb929d061d4e374c9cae5eff11d9f3dec1f2445b47b4ac807ca687af304b0958240daf43dcd74944345e8a594f9db26504badb3928a1d7976304336dba12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h516f9aea476ba8cfdb9a085d3817461926893d0542ce2c26e2730937067ea161b8f5533ed34ac45834177f5be3dc00727462d6dea24ffc821ac214bb1b1caaabc3935efd9a906ecbf8cfd4ecf0e8f8771d8a76eb4df579852fb1e58fd18dff4e6573;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f5c3ed496bac011aa2af64bcbc181197e209c845ec49e1885c05380919881d1346156ef364d3c13f8eb37dd97c6a3a6f21ce909ef947b896b48149328f0643160600de732baf260d5c4b39d0104ae5119c0a802e99ebecaa927cbdd3f2549bdb7b9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa821a6cb29939f4680f537e82964a82b4cab7a3b4473491ec573adabdc7ed811d0a3234165515c3140466f7e6097b2ed945da389b141fba5f16463d0276510a6cc9984a07cf5ae7453757bc5fc256950542e19953d1fc701d5b4c017f78a7633eee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf24318e7ebebfc210acd628ce758f7171f64598b1f2d0dc89cdf498ce5123e791ca3d451aa00ef17fb28859f19fa04b9a5ad56389a3f630bcb30ac0ffe6585b83645195db54a259fdf5dd55b1ba2b736d31c58a78828b1244b2dc3aa948ad78e36e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c543d1522af687feb8166b536469aff56120ad32c5c9572459ea2184cbdd86c6bf937d215a638117dff22aadcbfcb4015f25110db13077a8297847f96ae54fbbdaf57effbbf33c61569a9abd8ae538f199bb840bb50e0fa5419b3796484795b4cc0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75f549064dc79f9ba8e9e0b956892f74b7cfc23125b2629148c180622ba17845c67c3aaa8db7a54e234e44796334d208fa39f5f91cb048c3f5720d170a5b79862957608d5c0250273f734c7175b487641e04262fbf274b5d36a641a2ac47c2e5656;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc7c0812bc83f43e43a316a3c4665193a04896cc387e9b11b27fbdd2fe9cb57cf318727b2e25d380d492a704a5f281ee770f9c5b24dc78d32db577c4eeba0f188afa150d3d144a65b0b2067d53a1e4e9f0c2ecf80e5458d53eecb6770ae32bb15fb92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2dbad5e433829dbca8994770b126f33b400c362e07dc9c5d00cf0ec2f4827291c1f8c732be30cc38f2c8194e7213fb1fa5408583b09083c6a3c6a260ec9f69e409b156107b7d0bf06021a950f012022c7ac0502a3c50e2197c0b68d9cace12db226d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h457f6bfa0cc4449b18f8f8d53d1c96cccf5336d429d83cc263434a79337e01677054b72c72d06cf2ff17f02b96a30d1b33aa69ce9987fd129c9ae51b9fd86f5e1e209fcdeb2ea7fb7b3ee6e24a7dc44cdb8d13f28851436ab538277b9ad23cc43965;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h527e758203ae2e29e050cb4e9a7db77025eaf641ec61a416918ac2a4427ef0f6b7a73ccfaf2093bba1c6d1e3599d67e577437eed932da6f26d98d859c6e970bba36f147e8ecd77e12328d1bfe1eba629205eb215ee2f66ba9d45f4977f1e1a6566ca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a5581ba42517f10f243954ac603e5d7ebebf65a4f8d06e76f7fc5abdbadfe0548a9d79c8c7fb2a6e933714d1b8422a2c2902e84e54cc34e8f6a9cb63930b6679e7e51a4f3c7a8c177e128076e166f35d21e162d63563f8d8d27b378cb037982e6d7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d546785f4164dd33ca91ee35a9bf7c5603e034e8101d820ebbe46a88ecf53ff2c8e566e9b90e5c6fad43d1133bd041121f1df314a720a36ea67a074282b223374b4e09b1e5db743a8965c0b5840201999ceca6d070321bf49597627746057e2b42e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h778ea0599681c060fe9841d9959a90a51330b7747dc8411c4d8baefcc85f3e0ade9e381c7d4696ed4e29f900c17062cb881bcc9445c9ca97fd08173baadf90934d1872afd2c01ed5680e2178845e4b75888e5611d7aad5683087f30205b891b89210;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd1924f89df82be93fee920c721cebeea86eb7f65a2e755b6fd0d2c291be2dedef23cd10f471a3718cc36b2674c74192ae059a916eeab15601f6ab428ecfa9fd21e382c413d7edab50f86ad91f4a639bdab2a63ac41a8a3d711c57b5f355d261ebd7a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe9833e457495289a4303345cb4a72bf891069e62862c42affe0f388fcd94bdd701c557fd7e47c3e6969a08be81ed432f3e5719a718efd274cb31bb5258514e40718805403625900b0e5025cf3ec163a3b78dc018d02b5b914182f3474bab14502b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h60eca0d74affe023c48648231934e71a5e036352e1ebf75eed051401c020d1fc6d3636e38c9a6e62eecf537f1ee085a4baf093e27c480fcf74c4a3b147ad9e00cb0522dc9925d10153248b4d690f2b6e65f82db8349b0fb9b6c330949a505b62721e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had9fd4a68663a3777248b7da3576bc3a990612ac5e9d35cd0bc32819b7923ee01a2537cf7514a37a368c84f56366706956b0b3f23710190764cb334527a829078507cfb8317d13e9bd434cf3b6d3d4301edc24e5975fa8500c19d094454897c2ba0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8aa485006f317aabfe84ae1d7b532b5f7922825138c8ec37faed98be11bc7f4af2d422c24d9f5fe9765c4e806c191b8fa994033cbfae14fea8a55bd6db1bf5ce181ee7483fe0e2c5acaf5f884d93a9e16ac9188e1dcfd2375d5db525532a772ccbf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb02e27c608c8954f9c4e2dc001ac671f7f432d0f486df7f6bcc585ac14d09785e3fe8337302761d8f27fcd99a3f76a5cef1dbbb55476ac2ce67744233f7aea4e1d82261589ee907c58cec76c1bc8967182b5b5566cd7aabca55cf4a05d1eb505bd6d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h180c7199ea3684da384598688ac578eb7fd50e396880b5bb647a168dc7a0267ab248f5113e3df04d0b40a1c7c5c50d463835f1889fe8a0e35eb56dcf501bee1c5bcc225e3c4be9c8281a8f834c02d10c5fc0cbe81e199b37412e84afb28841909ef4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf835d44010aecc5058b0b4bcae60f0ba1f518980e08e1c99fd24531863b1c0516c67a71815e6df1cfaca0b49371396f20e8526ed2066ae7480b5fffadd03aab9e957863dc80136fdcb640459656a687fbc81d3a6c4602747677b9d77a9f05d70960;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2fb3b146fea490044f29cffedb7f68d0d2cd6ccebf45ab96391efb155b5fad180a28b8cb5aa15bd335e6beceed72967fd1641ded5c45a6d47c9b83214c4150e607b0e477a664b34d80e8a77ca5f9d62d7e88e72e01472d24f0a5dbd81e815c39c4b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6a2724605074116bdc87e58c59bcf06fb0241cc412caffc9c235290c78fdba39f2762e92fbd0899258e4068ec38c222c9c838f3019f83c702bb25524c18ee8950119276b2ada15b7d221c1e6a49cf2fa426062261e8691212950155dbf7cdf65d35;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15e6c267ddc6cd34dc0efd17fefd898d6789ef38a9513a23d3804e9891a9c0feb7457b25947f7e7dc2b8c2becefe2fe78a4ff0ab8567c1db1c1c16ad7c4c9f46ec208b818ee9e6eabea9e13e9c59ab2aa6888c863549628475d41e8f2fe612b0e903;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha164a2585395de54ecf6e6c445738919fd74f5a46949bc09ec5b983e4bf6cbc79a55eabad4e75035b5f960b3fb435f3be380f4614675e106a3fc8123480f01939ba85bb9e8871bca2fc38d0f876ca1e775848589670c2de3109a477816a1f0b43162;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3440f6b3b3c72d9085b2b0b2482542047ea68cd83d5d4329b4a537e34b4a3e59919659fccd35b3f59339440e19fe0bc7a6f2afdf79aa901a9ae9038100bb4e7daf64c60564933d5e669920e10c77a18080e8e7fa07cdd775404c1e344ddadf37a796;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d8d2b592099474c87f638b8358bf275acbea504192d343e8aedcbb484aa7a75b96e9a57ff26b2d01ba3db713930fa834295a9bfaac498f810ec4543ca3981ee598b315b466e9ddf55f3f361c2cc376cd3425a07f534f9e9fa0ced823d60826b816;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d9c4b3dd83b38e6fd79eecf96faa1eb86e3321ece21db13d3f1387b1ef78735babe707a75a11f88e43f78a693f7f2a77498c02446da79f005b8e0966a76cd009b64127b21366531cb2396bd10e7910635223b09f783a81b263ddfd8f1861bbdb2b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h578611121bcea352d9b496db1d4a7386b33fba7ea6410d76ecf2c8ec3465a5f5515c9a0193f27c03f8c8579d0b36615f03e7f1e398370cf582b4718a8ecf8874e5db5447efce6d5c3162e664524bf7e30c324207f37ec4b487b62cb3f8e06d9e9cd3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36e686ac2dee9e06ba58216b30eda7c846eb8dad8b5faf88e6642c2bb25ff7c3435f73c1d644da5059a7f1292c85d7d706933a54c9f874c4579b6ecc4e75803e64ce7105cdd438b6324706fbef34612c4b4e5a383fe573fe6252342468a74c33833e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfed24ec561940aca3a6e57554f6011ef2123cde05b32e4fc5fbfccee0dd93494e44519fcffcbb07101ee5dd136d395f58187e2f4d1734b385ff79727465f8d2449353ab9340707ce00cc9d3e91b4ca7d969b897aa3306fb1463b2ecdc1fbc632e972;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbaf6aec2f5cd356b5c280d21b887b2f5624e40ba8ce1132a0102c836b3dea7a5d575cc67a9f423123f6ac34a35d8f21199ae75b17a70467fa729c579157d15d916bceff0af45e347f8ea6cb041c679c139749375b30c60a39de86cf9ceb418f2029;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37127f173596bb8bd3fa7e263e0f40aad2d1b1f983d649b6a5ff2b6c094f6f091fd6f6745652fea44289072239bd3aee6e3c486bcfa6582c31694130f6191fc9ebe56e723e4dc7b7a9f30c47f86eabfe5f51636fa06f2a4b9ef4cfac891fafb07907;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d768b836903a7608d4b74d9f3244eb6f26d3fd4060b5ead50742804adb92af90740d4f0bcd8fde0f2282df18df4206e40c82abd619ee6e0a1851182b5cbc47957bae8bf9e0888ded41383c47078f42a60c7f76028afc01ad2a0f3da990ad771a472;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf571e0cf4c79eb8f8e832ef93e954af0336ee11833f6da83fe05aaac9b910d4119f29327c9c96ac1abfbb7565efe7b56ec48caee3fc2cc1d30c7d39cf53418447ce61ab10de4cf48fc914bd58104d34a162b926146815de76e96755574235831f4f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf1c462662132eced8ed16d9c14505d30f4124e1a69087c497a949efa3029ab543a0f6d9691e2f2052014d85e63817780cfc63ba7e3b3a8f15cc92f3acc41209e6e56338f2c3bc91155c451c54110d39ce3e3a404f5fa792aafbf4692b5d5c4ebf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77f162c721b10aa07c1fe30508dd50dcec9d949e6ec6a4025a9a2849f0a8b2b87eb20543d592744ae1b3fbc5fcd3accc5e293192578a99d338f9e48cdb12eec9503ed4d11a589c99aefa5a15d5647b6fba87eda6ff2ff1e90560b1ca58942c8222de;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfef2da66c0abfae7b44605c81dfdbcdbadfaf51a70293b4ee09d6713687a0ed45e763837d9286667ee4f8bc706ea9ab1ccae39ffa6a5ab9cc6bb8d4d680a93ce303032dd00023c36a608c83a72dec2e5f091fca20149c81575390a474764eb06d613;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd149946f7b33d88656d293a6beeb97c9bd830282cccbb0b6459e2a995bd8dbf2a6777c73d3c54d82faed9969f98ce7e03f0f863aaff92a9314c988555132afe9aec8c4a44ccfebb5e662ed9774efcfa085fd90f2252e99ddee51cf2b2d3f0382b2a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca1443bb1cc83d023fd849baebe0db4e86204bfc48fe7d301464d2ad13ebef903d099980ab9bdeea9d4921ae3d0c3bee7b83f6c9908fedef7a37369c8590b3903a4f9ffdecfadcc37b266e955555adc2985f32d6e1ca8f50f2d72f14e19aafa155f5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb9e83a74ea40ceade249654ab96ca7a360d657421f6d7b52cb1d72048ee5bb54ce7d90c0dc081f905b55ccc6cc20349472bf9fc7958de495e6451c74e0b9624db6d026aec330bcf0acc7cb679b18cdc7e0070084ce0281fea9031af5ec02d574583;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h92e45bb300bc5c6e6686a7e9aa42e3543048713b76dc022c6c7978edd12bf77ecc312668c5442eb9d12869115059ef8d40906abb8643662088d87e15057276db07225a8f00b1e910a45bed9f9e0ad503e13e01bc4787f7752c98f47ea0496097d6b3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h108eb72b33746786dc389c400dfc86e060c7108ee97e5be6865f1c05f0ccdbedb6b9963098114b41763c904c3d55773ba57c656b91fd7f38a14ce3567e86cc96c1d13085de4eb8c003f493a8f8914afb155a007a74a80be9199ca80168fa58d3208b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ffa3ef516053754d42396a9d60df51ccbdbbb78d8dfa690e900388417b19a7af221ac434032fc92803bb60b72d3609776426bff1b31c53c70f42b3e67ba17cf37b6d59e239a453afe26cb622aa7489e57828dd52f78dfa8b243d629f31ad184ea41;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d1d63b79361ca78694744b9a3b432d99013985590a6b19d6f771a96333c7815d76d44d2baf6d4bf102d787b8be1aae2bd4f0a7285b24bddf4f5efb7ab365c672de2b8310f78a49d2bb2eafcead71fced0e14366e6cbe3dca0612f4462e5cade2076;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74e764d6005a7c8629ab38c14af2773360e20206f49d02870df890c8a200124cf2594f590f656ae057e7fd5df85d4a6b3a308475b7b3f213febbc2cc131ffaaecbf9fd7b78eb9668a762cc2e95a3852ea5adc4ea7871cacf994f5c2064c704061ab8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h455a10c0788d949c56b9b9575e315100cfd51fc31d91779c6d2a60cc6acf88812dad2a44efeb3fdd0a561282f641e64b50144236d72b7703179fa8d975fb0f16ce0621d6ac18b9519fbb8f85524e83b9f517d97ae28370338828d5699112917ce0cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95911affe65be4a6829c6ecc91ccbfc75be7d8d1347a6892eea6ce7f366a5324b44f8fe87adec8810ce15796890e9f405e5002a672a1d67d47ad97e7b0daf4605a694cf353412bb2ca8214ace26bb5f9b245bad6e44d09a56d0b8b84af7a931b141a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h812b4c01d1129c8a8082d3f854853cceeadce8c58636948999635d4810df37a6f5d845500e021c8ddfa904e08ae84760955ecd9ddb736b8e74468f3a4b02587ca94b68361c9aa482265221ef3d5a68f88b565720f94692db36e7f65e5dc70cd583c0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9692a6c923c9ab61d4d0bf05a360b29dc156be7b293de2c53a27bd6d5462f2f70a1aafdf2f825b662535443c1897b4ebaba01eb225d2f2f550a0a6ddccb770f8744f0b1e9fab858043b12c9acc18b9b6cca896d3ea5401d4d8cc34895b09cd5b24f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6a566f1becd46a857ab8a0025afd4b11f1e6a4c1513c3f44e752f8e46c8e5882099321e3620a4ec77ecca31abf43fd6ef97395c137cf1c6d9a6c6b6b1aa99099d0abe873961f666735beafe663a9ddf1e3e4378431fd4e88f7f028095a4ebbb0694e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha816164cf44a51f14669e5c0f5f1922bc92ccada0351982493b0e7f5b4bd58468a3d29da56ff8a0b141482503b5375412ee07d4fa2d66b1ceca1004a869e21fac037c363386b95bf3317603accc0e2305ef1d968b6d39518c6b2023dc86f73992377;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6cf6df677d5f230185db257fbcbe01baa4e8d82ce1329221e7e6f7eb313b4f31fc455f06459f4f2f9737a33b2f9a7e6c0502ab3a58ac9e9b7a5b8948524c829e03a6716238f12a8dc0d5ef4f69e1583daa7579f116aa3b048fe2c9da2642c7c108a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1264c547e5f2ec2edc8f778aee3f4a821acc22940aa8f285541194041c0bb7b52796d7d5e9ba63c290abff5f77772b64d84e4c73ecc9c9b72e772490f5ca59ef14fd60e6ce55709756f0eccacba44098dde6c10a63166d5a8b5258f3a7a31782e3a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3cccbd74b55cfb7b958403a1e62a4e507dffa8316ba8843994781e7d8e57810ed08a80a4315697aad56a684d434e4f672a17963b8a1df19c9dc588551af5101895f6538cd6b4130d2a2cbc2392c42c3fa9f98f9ca1a33d47beb82dbbca4a20841682;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b19da5426c01326c59485b8b256457b924b957151237673dccfd43a6a6962294fcfae4b9af37948280a74c76e739d9d5a77f427e6a643b1287cb415e825b3794567da55f5b27969e914e7d4bcc256d444ea178f9ffe3a55cbf6a9fb746751a43748;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f6ef4385809c1fa42285306ff7ba318d1006d9f6282c44786351234d1fed0019817272b34dcb534ce9793429a17760db03f44615f9edb311e2925f80308465793234f650c1a9129242a2632cec7bce210bc44c230452536681418949d1eea0bfe20;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c6398ee5084e4c97a099f0a3e97e9071c409c898f64db4f3bf51472cf7c205e889072be71722fe328b07e7016ccfb445a82cd0e3bc42d963e54951e850d5fd5b2fdb45ae82c4bf6a045f444bd0746cad96e3c5167828058d4a8da09fe5a332a6af6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he038fbb17a563d90f5f4cb0bd989dda0e3a8e310d5b4cba8c5a4c9c8d0a8f8ac1cbe06c43042d249eed35fcdeb99f42b268042236a7d4f780464ddc2fcc5b6860c14e888eed96d8feab25b7886d49a59be2c5c083803305630ccfcbd2fea7a00dbc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3eab3d2bd07c7cd83d8baecd019922e2d04fb1a2557546bc9fbfc17d77cab67f4a38a8d70c9eac25e24c0a23342a883a3a8b001076257a685e4e109226cb3000f817adb7f95afe1216513d1403f3c010ae7d5f5463857e37565bc7a1dd0f4cbea675;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he074dfbecb75ea10c5d4cae0baaa672a540069574d6468cee4dfff90ac4ad31e791575d5e75c779f22809c434087cef96a088bb3e6a8928d2486fcbf5ee310abcdaa9b25af64385665d57bc90f3466163500378248809263010937a4bbd83f4e04bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h915cefc02855ee7cb8a1fe6e4d219a8d1ad3f9d8c3c5f206318b2c407a56ac5df2b1cc066e22c5931b6559f2429b75c5a30a858c78b362498968ebc127bde653a794d07c777539f94fe00dc6ea433a31eb1b020830b14844ba0e0485e87679ff09ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b54b4359ec38f5989dae61958742b1181ebc5ca48ab8d9c68a6f0fd3c6166a2223ee92bd32683195233fbeff3b2662229c9affde8a090592a27da4834fb7716d755c35124fbc054faa8e26d98157bd9e8a5201de1c8fb95b40b896c0ee2f2dfa90f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbd22f6eb740bc22fd9b1619ccf360c7f7480ba58eb7ca0d9fd689d62df712a7018254fbd67fc59362024862235d6c4473d6d6692d30c4a082d10a622ee8dd443c5d831531666d669c96f3ea7c4ef1e2329a5f291e7be1e9d31b3f6453fd2431ebd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7161ce88a09f32569752acf566f2130de77cbac2e82d307f72e6e6387ed9a095e50d896abcc5ba311a8796e177142292f15046e75552fc34f9c6b43ccc768c1d7ae47172992c1cd3c542dbaf58f601487a9cb16e1653c6e19279846c400ca7c1f19f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7939b99053125700fa163aa3ad90482b42af9758e4d6dc9556260942200fd7e3ef7633d39f14ecb8dcdeaa7b08eb2f7cfed36ef2638acb9d32d185582c895ed25ab82bc5e8c0f670ac8cdc6fd48e30686f1fb0127678f924197cc063a692586f25ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc61a0bc714fb995c35b13a221c2a112f9f579a957ca7a6424ba457cc236ffa16ceff91766ad3142b6cc02c31c7e2431ebdb4799d44eefdbc9c9bc30101be19e407d070c1f6de33c539bed9083900acc3e7be13218f4990875416ec0ba95806c8e5c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha10310bda29f7a82830389331156ff4751996022b26019c7e209137c2dd3544218873e9c9c3432ab71384a5270fe4c16ed3b8b7714ca7426554f54ec3a60ef323b786fc8435d4a9b9146eea450b191b69302ec1b0c3961e18824f6154380fd94bdfb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcacc4bec5b94d9db57aeae723d5b9d8ca374949bfc83b04994f97134c2d8b6863e5788bb787c8b451c82e268e4fc450638a698f170f1122cb438bc765cb0c14f60fd9792f28fad45c07287bd22b20c461650d51e19605e3fe4579c1d938b66543fd7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0b5c4102da0d34ece98fba9814f67bd4e82bd0cc452ba5f4756bc689756d66303719d8ec5de2e8492e043b19c62895ec6d675470b289ba30b91ed7d1fcf20843082ab18e333c184d33deda47670f95f97b6496a3e5df23664b086176c4a749c7663;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h66cf500c98d9da58015ec176dd6f47b00abcde49cdda6582616d5fbf5a729ef2f55ae1e569c404b6af30202bef5bd936106d49160393f3630fdd1bd9c0328bd569c527782046adfbfd9140a6fbe0a9ce4c9165ae2c086b11966388bc688a14f7aea8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h109358ee220b69b21f4c4a375b3348ef3b1ef3666c3f97ce4e6d4d2490306fc7a970cfd92caca16f42af6d009bb0ecc86799d0d24bc7d1dc322aa53ba12bc953122562cb330f38e3fe9a6b5dd6bc4e8ef6a3a1c5c6b6b8e12881f5e448aee497dcd7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9472667e92410dc08d3f518933b058f957ef0736d61a197f5abffbfea0a9829c206b3da6338b232b113143696d124a2f4eccde9722ab0f226fbd09cfd78a517fb188082200bc9dbde3f41d795cc3de3f457546758dd9cdd9cfa57075e081529b81f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef55cc577866062f46ea85668faebb975f59bf106cc438206c45eced38a716aaadb80d74ecf8d95f30ea78ed062abc1d0a56db0823f76a66927cb5053c33c854cc5cd81d3dedf6b4a26e2ebf361a28066d3a96e0baef8c62762661f5471af340a2d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d2c032cc02c970826d68914949e62252beb7c91ae42e1301f09a5cc1ac25bcf8eb8752df1c3df632ee44dc8f72a939a0bd023bbb2784dded20aaae819e258b6f555d68b17b7a72613577a511a6cb353005cc00c30b2e61eb0f8459e99bbca33d193;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfe6b571698be5510760019db588da2fc51bfa0b794a858598e1f738a294e5576f4e67eb5f2f1e8c7944b47e56978868aedd721a56d2dfc7d9120b67244afa3ca7cde8791a925276f054be70be5c500c0c84757988a057a59e41d0d6b9e504603dfb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2466062f59472aa2ba1013d0eea206edb8b71d5592ac481c77d1a9caf7174fbc5095543727d0eead27a3c831ca57a08e49c9d826467be967cd30a86da35239e631edd14de2fb2085638b2eaefd4207074cc36d939d6f883a04248bb497d8d629904;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h14a703bdadab82ba4d814f80b29164266eb426257dd7081c0c997bb2b2f1aceee2f31cc604e3b12f0b3d52a821d6790b7793fb6a36e97f953e6e61df5c36caa1b1afbdf03aa2d865f2615b4f33e504ea2e71c5b4d6f48ec71fedf652b37869ebc249;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5375de8994c0ca1a83be92364528d1b06ae7cb03310ae43098d26aadd3808abe3e5c54154c224d8a56ababee8e0525edbfbfce674a1a106f4f03b0841f0ebb3e67cf33ba045c95cd300fdebb76b2f8521b06dd40aa0fe0a6fdb4f040200bb7f6b25e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e73b74b71d3f29026d7424c4855cd0ee056635fde38674b87770fd0ae605bf5820d57fe8cefb8413a3a5f0b9e88d093a806a0c3805c82c1e964ecca678a77157d48662d56cde02f7d5b3532589a8fd27eca29b9dc3aef5dbec8700553a211d4272f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb5a0972d1ffb26529c6be1baeebec131984dc9d8efce281519f70af31e4a967ce542b7d2c690f616ff055f7dd821e65187c8db27deb012862996d56d6ce0c42cc1673bc11c0d2b8dbffb8bebafbe23bd1d9a36b8a1e2adb1e0de475ee0e73a4adcff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b26038929d027a635e35a1eb140405b8937603a269bf27b5fb7747609c36fdfd2c437e4235c2e5bbdf27a4c58c11c7ed589eeefeae14e9f81e7e636b028120c87d25907f953dfa6a2c7d21855246920fec515276b66587f0c538862a83332a77eb0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb940c546770b2a990381aabc0b709b448b9780a57580da05a1f526b715eb4ca72842c63230ae291916d168402b7a8d80207e353014f1444e21a8347b4fa3d585ea46ff94927df87cf9935fd1eb6cbf2a4a6788da4c531056a2c55599f51fd740547c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he1ec4dd04de069cc547bf7426e5a5ae01929e2c6e98c5a86ef06358a2dc56a65a9dfb430fba6504eb04910a026da7e2e41209210217a33dd314039fe95244f0e0063a98993633a7a137d9e1635a3baf807e76bee4711743700d7b74e7897da1b4b6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2b83147597b78fdc99ffe56381565546b4b85a510922bf9905960fea21797d294b9d496255381ef197de1fa93081fc7da0f1d04e92830d20903cde744e6b8c021c70b603a73ccea966f4c5a444b1639e174abaef3cb4d157f750d161f523497a809;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9fc3a7de85ec11e9541d41095b55862d45936b53de5ef5b4c66b051a8eee4d71d8395ef1e5d0b23ed8f1472093c9082fc54418cbd9fb4b4a2e137c15884495839cd471368c34f1b19dfde8e7d660f856e22bf302dcf1a3aebde9816cf5b4764b404;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47ac9afe389049e3ab98fd537a8c2965c684d5c3db77017ffff6387e47cd6602b3006edafbc570ebc89334629d1a07806d88e79102544b9789288871ca1533ff4715c31ac02c218916351083df707746ce2fea03cdfc6cbca60f4cd5af63cdcf6b6e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h830a758d4d24e16370685b228ee3c373866b067218e6e18b97d1191ee7e1de961e2571491872ded0c207a590107e4229d49805b869ad2eb03e260d61631f96d2e5df28bfe10ba616d86ad5c94a7bbeecefe0bf5343c1f0f8c3f5eb5b010b0e7a473c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h764b487b46854c5af2b5bfa4ac3f2710af3408e1db2ef2c3f968777f64da013f86da23ce594f2d4c945537877d76888fd1aff5a7e18c2ca22d6979755accb9d0e392e171b81a45464d02586b349f6aa62c061bb359fa502bdbca669e912d4821133c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8d672822ed75729c9162653da6773595aa0c74d62bbd4698e8dcea01c10057d75b90cc7525c425b16a808894028246cc7854fc94665dedca6a03065a5f7476d05dd3c650e5b1de7ca5b160bc1bd230bf7877b53f960c3c89bc5cc4cd53e45ccd07b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4ca37f9a472e74a8aae765bfbbdc30be9ed1d7c40b42e51b57537f126079226e189e5152ebfa7226f76f6e6f32da7956f7897137ee1177e00257c2ceb84ed148cf81a796596d950fe324eb3ab999995a7620252d1aafe4f4cc11217b7cbfda67ee7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c0597910ab6dc882d59e9c437528457b433f7b33505bc3d907c8a9d00def4a4658c1e1482d827012596416c13e9a8e5af99d8c1ba40e1bb90f30b04641df7b4cb715e22a9781e968f56405528ccae39e5fd292a7eca8392cf73c67f2cdfaee4c90;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8c85ae298175d1721a203e229eddaf7d2f080451ffe34ff4721cee83321aca7cc3f4e9b956599aca3bcaba0bf1c9a9b6ae94478a94c2957b63e11c916b0322c1359af75d1c7580fc980eeee078a83da926eeaa5dbc2c908323901255127c22bd08ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc01c04e4caea729f7e2c5985567f27a7a61ff159762a65e766554256785be377cafeb257508f91e4a39dfb0d8af9ce72bc257d2da83a0afa5d44e45209629265dd7d2055cec1d731d353cf05e1aaf066819718bad7363c70250ab3f84b2ca576e9fa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49cb5f2b58988f0047799641eb7aa169a81768b62c54d7358d7474ebf55a2c5cc8cd358b19b7d2391e0d4f1c15b5543ce7e19c4c015938b1063ea5c2b257ed44b7429e8a0e809fcca9957b348114c7d7148ea74d187ee69733b9ea7515c679cfd6ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfbc4db2760b0f322982106f559d896a7ffd2b95dff747a5f5f601e9ba55982a5f7c8de4cb2526898372fbf7fd2cec0c3c4db44f2a2d64e7eff8d9da1bd81395b4f0cda667d8cd004ab5715a8a6afdf7f4719b3689dfe6924ed17574e42326a86dbf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h406b66daa64b5116220169f077b54841c3565b41d5fcd16587542eb65ab0a19603f59b4c4d62523b0ad6a5a0097bce53e681f4183f3028fd0a183c3119328190afa9edd726942dad61f3b2d43c8d103955e6023df21b7ffb42e85bd5a395481858ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfed3399be5495ad696bc336ac8a93a60487c59f6c06c350380eddc524d0d30f3de881201085ecead77f055d7babcbd1c1063a8655f2f97cb25f8ab9ed1ba7c5dc6dd6fd47227e994719789c8340705d4b86a2d20f6cec14dcf941d14e69a3c4ec1f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41a0e2e84f362385f71ed8073611185badac46e7a5c1ccc5a18bacd9b7c71d30fa179a60de17abaa67dfac78d9470ccb8d43f879ab29002d286bcd5b318afc8587a1745ea03dcb1546b37f0ff32d818c8b33b116e275a4e8d2ef4151bde306d03d86;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a7f8f902e65064658abaaae2e31d11f0dc9504f40dc7ddfc0d342396e9e61720013399963250191f511dc6f1ab012a10ab6c7adce9a5909ec23edf4ae467952c1bbd6a21b2a5545aef0bebdcc6ffdb002366488e2572fbece273e8ff70fc5776b02;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb71353c70395a4cf4383624141f434853a7db5cba14d52aacbc9d7f4d9d22b8b5f06876b7491cacd7db57b0fc9029ef518a479ff2802ef69cb6bfdaac35e6085e3f401a34e276061ab58762df3d7604c35b4aae1eb84732ef2c463f010f292a5106d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94d4fe1f76ba765f13324f7ab9c8c266aaa450a52d539fe3ef44c1f94def18606e4c38f7f297f39e955b0eb9e9d75d34c8a3d31dbc4ecea6431012fe3c62b82d7bd05b23a0204935a9e52e6a98f6a16afe71fcd02f7221035e8381fae24be3b1d566;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacdad911230bc3488a6bca2c7c198b01c14b7670b6e177d6bed797b95e268e694ef4cef34f41ae8c9433b3294bf47aa9120544eeaa1ad1adf29344b2ed0be510cb968688a2c7e71607dd51bdb85f076a98d4cad096534264311f3576f34853de3890;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41b57e33ec6fd6f9846fb3bde06d3f94d2483664b602e6f7a911163fca32f4fe27518333639988579e635117c390d3539d0fc4cc9dd72d7cd7cca06be3c56ba34b711cb47c73d3c8c3b2fca7a89f1ff9fcef68c49ec40de36a757fd6e7b404a89397;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb96cff39dab22f5446da036285fcb97f95eb06fe684a37a5c5b565d68037cbfb8494d048ab1e514814cef7a2d1371d517c5e58475371568a15531350170979f2a0c766d00f96353cea4b8eefcfbb36edae65fe2b41f1145234dc622942f926ddfd84;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h30680931b236754d6b50cdef8e6d611d76a1696353f80c87fcbe31d0e10111adbdfb71501b3ba2a6c661ad02a7b08c82e963cc4019b9a33ad887209634db63652dadec5e05b9a3e255e4a1ce3f2597e33d78228d0411bfdaf13c3d7a2846a4190914;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e3c30a8771bf9d8bafa42c9723d5f884e814b419f6ee92683b07ebba6e4f2fbdb8ec977c1206e2ff97d347525fc53867c4a17d7e62a22605913b5f56623364c1b6c22f3f840e5b7860a9f36cc888eff134c2aeed2152a1e815b9c99c0781d9c4544;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b043115a04e5df5c561072f1eb94816813f0a1d87713f72da5ccc82f5f96bbd63812b6c57e8bb095964de6992ff34b6d9c9a0e5d893346f06720b64c2eb33b7c1c0d56149726309678cc1aa0e9b305f4c249626a25992f6c1a78eb60e120807735;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf985dec787836bb2639565622bf4e05d0e700e8250b49706540e7a40a5cf811db4bef1190ff3455c5e097992d28502891560fd378776f0a6acb0778a0e905ac6abfb7dd8929fe91ef86f1c30db75ec06f4f2d87c30e16dcc5d6a36f4e1ea6438432;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6021cf4f75f70d303f52e9fc02227dc5528220e768850d32a4f52819b43f075ff3123143ed764753d6d535580eee2c8236220af553c6ee7baf23af66dd23e658d61741eb2c60b4067632435d1a612022c478233ffd1de4a5c17fb3b3ce3b8112562d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd7311de450302ef8cb84d8f0b9334ca9db93b45eecfc9810c1b24856ad99ff2f73fce58de854439de31f1c0dcb63f1de93092167bd5f651f6b83088ad0e4f928c6ed56d8ef9332a4968f84ce1c35ef852699103b6a4aaa38f7f57af3c5f5dcd4900;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7945d1c99bfd0871eb85a631b5109c3fa5e4aff82e2e8f670563d9d42081781824a7ed335bb9e5ad730f9f3778d226c5e15eff3b9d0bfc8d7bf9b69ccf0e647c7f56f7562a4c432a1615458fcc176167dedb12c82408bf5c70bd26d0f377735a4937;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h670fca5daa3ac82746902aa1200c949ba65af882187bc16b55dd64ab753b7767f304ba4160226bb90eab27a401e0800366cca055f97d686038bb25a2f5be0e78b552759cba6666034b244205f6a776c85dac1541cc80654d5cb928f9255e397ca1e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6905dcf8e291fa90d0515675ff7d77a2059519417815fe0dcb6748668ac4e336752cd89ca986d6f8a1a2bf95243c68f2b2c511f25e8232f65ea944c14e8afc2542b4610edaf884de1193ca714829878782670a580acbb2e35c648ec139772c4578c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h896f541d9bb262eabd04177ce27264a23bbb7a42841254dc4a3e732f4a6f8075741424f6eafa522c86bafb376cab4a0891dca3c3f73a2d77fe937d2b2fcdf4d0012e8f2ecee18812fdc0eadf8a0ae10c51cb81e970bd485c51d733953cd08268419e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8ea50cb5e735631b0eb86770d5d2f0eb949267865f9e740392b61cb872af804c766004f5a4aaade2e2bd401db15e7add63b323e6232c27a579d7f7453b056ac52872cf5fe78d97051d6e505e0290a6dcc30974db220a640f0f372407398c0fa7f93c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17e3bdf041c6211e99fe05c4090468c92ea941db7fae9bbf79370fd9b0f39525fd54885ae7fb6764b022d193463201301927c763331119d8ea6417c642697e464700b9bf9f9afa9be618c0ab144121df83d874963d148e2281379c09ef5df45020c6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9c4f6936e1a95c38c4ffa44ca0966a8ea9c7a67fb1357a2c9af18e2bfd4541b185928c161981d0afb940f3111a8a79f04a289b33e296011989c7bc42dc98458dcf9297bd086705b87e59420dfde328797015355f61e078fd5c13f07f34a75ab08e8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha59448772e2414283921c25f0cbfbcebd1e250b71b57e3f47fe6340739d4ba7f0e872edbfc1478a33eab89989988634f012d470e75e90a5f72f70ac926785195c4afff231c9407dd93655551bd537ce9826925252653b75ebcbec708d959d60a74e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd055eb3fe3b69e8f72a9c774d3e38b8b09dfe00b436f9bed1fda0b7642dd89493cc705f8340d3af9c3bb91208a7c7f30686aee86581a4434b154f5ebc3cbe2690e60d06308c60373a58f921915ea5b8e4c75b696e51ad73fec049b51102a7161a113;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd20e0a560219d4dd9064df4e024ee9d47c94192ddc66ec7e6a92c540a3a9c882e13e03e0be0619819a086c48ebe43a4aa0fa320696d3dcb3e35c90164d3bc1de889ddf5fc11d494567eb227cecbc1332bdffb1f9ff1f5823babbd3ed4a9ab85ec1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5d6f14d91acd94a4d863bf0e32c879a7b7c22a53df0c95e5279723aa7bb905e262b99640095b6ce62f61c95bcb1dfe522d10271f2e37b7f51e0c5ac7d9f0a0157b3b9623768872eea8eaf25ec1721124a6a7896ca10c9470e3c94e685de6458bbf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h356abefe6a7827b4e5233deedce5f2f73614b107dc39ac7ba847a8b83f9bd86758e15dd1a1f5d48eef6d5e53b32f504f3e15594aa9007eb2c7ed9b61b4e71a600f5d67743127ca9d47740cedab9c94dd63e4a7eed1a41cf71814f84d64242febb0e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbaaf1193cd68e66b841fd37b77efbd307b534220bae5c6f8c5b4685c8a750e21b3dcbe7e84afbff5fd9d8bb9a23c8aabf78ffd602d715d4a4cb244df0b75342f8a9230b9fb842d9398588370535e117a0b7aece1128950609c811d64c111c0267037;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h352d84a8d303964422b7c70c18d8217845e3604dfb3197b5f44b380e8dd15eadfca5328b694bdf45201116d3285177ff4a9a2b381d48c41cda9c75258836e5139163d23c9867328a1f9c8363690cf72a81e78eaf5983876a3e4389d84355c0ccbfc6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94cb6a991344eff3b2d056c054ceb0bf0510579190dbed0034b1f8b38baeda0dbe577ecab9f70d1dcd8ca0e4ea65e734909739150679482194d32b0f121620393db268d7e0e2eaf08e605b1d1e3f0eebb852a023825ea5572272f2a08872e158c3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6daf19acd281b1f9ba9eb75f404a54810df8e956c7831b95f16717defd099134262d823ffe6e740b4fd3f4197903ec17b11b78ad3c4c83b8b4f4e7cc242495332e1d1e66b375e2ce987b588e1951529d33fcbae3d04ba650b10d2b216e03d2b3a329;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5e3c003deef2b09727a93791e2cff6db81b0e580c30a70da6747d9bd3866e175789edafac51ed67d95ddc47f7b27280f62537b2b3c465209096876c87f642eeff50f2e993a8276fb41e0e71c2ac4b37d2d14ff3865ae3447e2c7e75290cf856e0a23;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h809188d65d3bd71ee30c09bb8f9312e51f4cafd36f36deb96b18cec6f950ac15c76736de3a11a7a278e9df560e299b11d26f6b20eb85fdc2351a84442e811988e26dbb1d3ff713bcf7a8f51e1d4c841df596bd637d046d7d3885dc57dd200d74c080;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h807073b5261079f46fab7dd6c516ec62e22afe2787cd527fa9b10902d520c7a801a80e3fdace650bdadc60570c1b800561956152117a55489610605a901e7d10aff3332f7e025224e890024e283d150a25f747fa0f888634463c14515d17ba682e87;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb7d134f8cd85515bd4c6f9d68bba71146ab7acd604cbcb1d2b7e31c42096c8b8b4f8c998ec6a57044e9cae0fc6d95e9a41db3396ee3f7f8397e5ac4fac2b5ac7ededcc061da8e27bd5b5da68d286405738081598894210a48d88f52654c931f39cad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h376513b978ccf225e573516108f9b8d03773eba600333f4eefecd99eb19f07ab9fbb3b5f591cfb61027b2b297a0b9127a651ce794cb4a8794b26f0e0bd38e7be6b6be018f14da0a989e51ae6c2d895c63f98808958968cf4ec0e9ace726bc250bfe2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb1772c86e1fd36d57e89ea0ccb49ea64408cd4d8df5b32b6e38925603bcddd17de72afa5ae30ace6c4c28975109d987d0ef2e035ba41f3567c161d5830a0f901797d90633d74e53ba9c1a46977b3824887fbf4d412b22b9fcacf01e8250343a3e178;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he35e37a157331be9afceb6e1f6f36a4872965d241b727528634b20ac8f605f77f43d63ff42c386bb858cf649a389fbe3f19c64cbda93faeb5fab705dc0e375e03dfc0ad18f02ec56cef115fc13b1e1d497f5bf57eff29f44f3d9bc354845640f2981;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3b3c2508339bf3a5813c5b8ece2d55e37db743ed8ea0e54037da6484172662ebbbf51545b7aebc358c15ce855fb440c4a4d12e79654fb1ed1fbbcb34d1b711a2e01f5eca567d770cc62c2af599431a389bc9b2bbb2a5a93e17b790fed24e133c1793;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc170600661bd00c6608d5cf3724307f873ea18607b86c8efaf1c8397faa95d608d04efaa65f2d78d1c4ac67a175969f91ad267d4de4af0b913c9f6727bb40a4eb7bf50a6e493239a6a41f274a433a2c307ee66369183948a94aca9e6a5b2703496bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9500c64dbcbca4bb3374fb76f8f3d48ec0a83c0eee680f16fd1bd8f6035631ef27ff5065350ac5942fd1b874613e3a5004e090855f99b4b210d09254aa49e149715bdf11a1a6bfb4aaefa8113745a125e77ea94439f57361bc46430c2d4aff3e4775;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee8bf880ffd1601b9a21d85ddbb50dd76fd778ddbf38c3d95f53c539137d1525de52a63d967858071479a58ac4911dfdc1c72e6ce240e45f02acad6e69f2a2c2772e27ba9a0694e9f616c937150e9d0f078e9633b30b10b5c6b8f84a761454abcc5c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e61b5db1dbf46491bf35156f30fbc3920fd8d29f52f3d05e712ce63ae1da280a72f700676f669a268ecb1ad7244df399eb6a041b7496d142a44f39cc422d68738cbf81a6fb0419e3d1dab945fd96aa686be9a5d574e513b0f00903e72903ad369fd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha1722c45655b1c525486b33e82a49747ebda1e71562ed5af092318ac8b378a529b5d4cfc77a154c3d873f51f6c595b1aabbe02b0ace15bd1cee07ed0f0c4d530d58ccf1933d75078d2613c050030bd3c27591a332f6ece4f2e5827dc454d8ff45553;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e9cb35fcfb71d60481593bebb83ac49ae6998335d9052b2ef92db64852b6faf8684858d137040bf21a3e41330ef6f7cbbaaa0df125ca59192f8273f43021f979f52f69296640c174abc11ced34ff54140e409c4da743e24993b8d03415b76c48160;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce053cdf9cf4788da0d0ba3b84b4e1ca46a884104813edba5b401b8ba9b18d9c51b7f9959601389f623c01fa8ac8ddbd77cfa7be4f19971b25731ca689364688f52f1fd82a69ba363fa0e71fecdbcea1d6e68ffea2a22cc96a6874ba5c47ac63d9af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h77127c491f6f1f4452910b51657672e95c7d6c4e6ba6c51ae0596dc9f8f76aac7aa966a9a020024172efc813e8d6df90b3fde11f467e95f6028557260debecd8a10bfce66f0d004f04ef54fc31a8136b56cb60d6797746bd7e5b1ec3fc5ae8088282;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2f312c4cdea23abd6fd33ee56ef5824af76fe3275ace9ccdbe1ffc9ea4a1314a82778728120ffb4ce2866db090d825c2f0f2c7187559567200f5ffc334abae5736b23aa2e8283e37ee53892603e04625c4a52a2d65c6d34c01444d970bd515c8748;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha166f025ffcb25594e62f5022a3860697abe94e1dee61190ac092a41125ea7290706a4aac6ed7347355414b79f582a246b84b4f2597509dd24728ef0f4a55de68a088b70f3d347885d145364b2cefd86aa21cf8c6b1f50a36a700097a459adce10a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10192d708ae76db447b17a2dabf99ef81973bb87dc55b39efb903d8289a070d282a333eba08f1f31e70bd1ce4373a32dbdf2e5e3242de3f2be0159da98c187f0d93136f9f59fa80255fca1f50d4e868ba1864f95e6f30c04ced58ae98eadd27eb503;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a373d50efcde71da49faf923baabe8cdf2fc8e09f9aadc01defb10e45095f3afb2d70a45feabc68a6c660b1a9fa73f24e4da380c06c035ed7f848eade061c3963a3710a71141acaa27e583b588904a92c552aa3d880b1220cd7e9a310a13d21f91e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfedc5c1e24d03364b02f6d3ee8cebe77cfdd12d1f597b66dab6df43fcfb351dadcb9cf35cb97267829bd208e0f4208b2a4ecc60148fbbda813a2ac50e2c7f5b64f6df597e541e2aa96abdbc3c88fba402706feed9fdbe3f51eb4bd7110219696d98c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d359fa31527f4581b44dcedc2da3b0701e0b00697c2bc6729ab11918f3adbbb25565f590e3abb023f036310a5dbb54356ef58f617d5df29bce12a7239cefeb2f599fdebe88a25f146476752a2c5a0c7950e015cd5885e998ffbb02d9c666b43decf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haff2dff3474875071e36ed2ce5588ba7e1f49b4848e9808226bc91b082dd97e0376ae4d889a7f4171da7bb5bd3b324702f72d3ce3697756149890578128be211622cee5f957e220f316360707a318074e5646369263f3e83b0a44a1776f3274615c0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75c3e819855c7ee2fcee80bde7499bfbb30940ba43f805b7643926b5572dab98fdf1c2e8c25f55d8fd36e93c1974a95a916f057c2936811472682d18fa649849bbf92ff451b7669f13e1195eba1607790a59fb43ac84b1e0968bf992fafa3bd9c59d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d2f8d4c5f2b808e277a677e05b902aa4b51c9fcd6d4af6d2aefa20df5366ac0501eb4fe46e7d6e842a162ed0e9c2635c18e6620c7d5cd0e2e833c88bfb4092ea47a790c8eea30c824241c5ba3c879c0d8d20e3158390f05131ceca27cc877fb3851;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8fc19df22c9e702a77e816784b804d6d4444b39bd2bc84b1ce133360a066b85a02f5851c71046741fb784aefada2fe0fb13bbb8da1fca30950ec8ab5b52f40b40508d1383839c99eca9302ab18217d87dd1a349b57ed8e452b94ada52b7ad6dc615c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h989b1b57f914f9e4a80d59c804b018a6831a4d53761a3ab8a241c06e5844dd26f2bd35bdd5737c548e0c20cb62d693105c9a330c166ac29207769375fa8888d8a31842c313f2e3e7e9526db2006923a98a3b18d291959c5e3d95d37b15c7b7d34130;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58a7e5afb20fecf0040ec91e834215b25999f6df75e0f9194367744ddd9ec59a6e5a61de905707e63656f9f9528cf21b287a346ac48dfd9712997cdfb2ec269147788ae0079edcd9398d406aee7933bbb1f4551160f17f66115cacbb4dce165c4447;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h486437e9d17a74136cacd3cc6547ef1a2c94fd1f6c218977deff10d4f2eba8d1f1599a2ed6f8f5009140e49b8d0098bae737cce9505adeb00921a054efcb710392b9e3b1f40e5fc5238db6c7689521a8a53032aad884a718d467234fe537511bb3e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha146e180ae1b2b388c142c4245334fe7be812f1ab597007880322b1aef6f6f08f5479151cc586cafb825c81c1a331d6a9ca15a3e72afdcfd08cb54106794f84c47e1e55976cc69822f9b4d3dc9e1e651d5b1470e57c41f16cada162a3e3ce2da1e05;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h87d5e58359edf17c1972767658ae2fdc9dcfef52238e03bc4517c0f5a9f2ba7620d751c377bf9d04425747b196ddd266fe7251c72791b367b89e46e4f531b06835c3c1c6747ff81914f12f7f405b5b4eea5a7f9fcc433ba33239e05eb6cc169a2048;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e3e421bb65978d2b4f0cfd2a10c86b2233c099f67573a727bd3c0c26e2a9efcd974710cf9272daad4d726730f5301d9997cf3f38d5dd179ff3a4b50ce638cdd5abb0bb0ed3df9f6bba50477d7dd00cb482f9d1ce44fe8b282146c44faec3a56579;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3b09b20a20e6ef4da3d75189fe38a2c717ce844694629c9621bd9c75f708bed56ba6c27e6cad15f1520fecfd6163e34acf0d017eec8c06548ebe98257b262828bd627824fbb49934ec6e09990dc96cec99afbe90b99a43c36dc1bc1eb7eb39dfbd1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5a68253f902a83d4278d6ae37aca8a4a9fb12e73fef698ace9d5ecc5b4bbcb4e75824a537689be1cafe9a5685f134cb8a3a97b8475714484b1af02e553c6dca4c8aac5c79e4326b40f6b020345c315c5eb1daffa89abf3e1403590bc85d6869c018;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd796fc811725bbdb5c80f9965fe25220b84c08323d052d08b55f35208620a7f1106e2d6d6dd80eac3af91a6b9dce368a6c23bb6f8fe9ae9cacdba6d5c441a76799a616ffab489693b2e8bd1c4530e5ab0ee4cf8346bb3b75bf59ab57876a3d8e486e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff9091f4b11dd6835e06d0346c723ef84f7884a4f1308caf948b9b85032fa0278065817bb75b19901b8c865974691106a214c887f98721fd72af0bf95209df1aad9d3fd36a97733bd067ddf2a1a0f9a3243b011c691b739fb903b690cb422371dea3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he5061b9280d6bb843167e550056478accac9e3f289585d3176bf4c876f13ce12d9d508fa900ba3505ca811da32dba9f70b41f9a685beecf3e10065b286d8f752886c609e2d0f153a096c6c67f1c7fd21f142f21bedeaad5867c181f2c10148291363;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h34dab9f78cb2607f4e8228e2305e95f8c223e981b41c6b42b8ee17f2c9ef47286c0f483fe3ed4bfa018b0089a767f757f6dfe0c37e6b7718c0de2ef915dea62c7d9c15f1e67aeef26d24151996f6fa8813f82ba663ddf83250338e1b53c2fe2734dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a708431e2e36bd129a605462a7280dbc7768d53bff9cf3a3744eee200bd01e81399024212225aa8c660af439739349190e8aa74f10771b8c6a4f6a5fdb17c40eba99ab422ba4da3841d2299258b0249d3f25ca46b360b5be2ace87192dd31bf6ee4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a3718abd0418c46931c19bb78f927cd69f2f73a39fc717db0c63736977b86d6bdf1e4701f39b51e71f9ed65de8f4fc1449f70ce61c814d5d8f94ca63b5bb9732c1766a385b2419e58c202e2367b21c06b992c497a6cf304a6403ed6b87676a73040;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h71829e2132e0d423244388d1d249a70f8125d3c5f416fdfaa17e34dfa226f8db33a41fd9c11e5b2e615b850c0e0a5687aebe74d0e3e6df69141bc250049ee36d55cf9f7d9557c8dcec6008a080a26586bfb8465a263c8043495daeb26fd80f69dbf3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd1b18a97141f960b0b9b07cf33068ec6e578346a24f1c39ba194cfbe90cf8c790ac1f8f6f74e6cbaa7bbc908a68c3b06929f37edbb13fc08c5a5c080e0c2945a5ff2812a35526b80a9519434871e2f3055b955d93b8d205b298808550611d695e6c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbd9b94f1c7ce9c71cf1a6cdefb3c659b5b6a6ed2099c8b9b304f19930d6a8e86f0ae461cd470d5d6a66a050a3849718a58a8187d2d71fd90d3bb211c83e86be2611ed5246e78b107a92e10e9d98aeee831f5c4c615571aeb6256d5e1946ab240a6e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36a0df4fbe6fcdaaccd885b9a624be55112af49288f9aae36ef123a7fb95cdaad916f29c6ef0ab0155b0c161886b61c3f1fbac69ee6deb01963863cff6578cc15589cbb64a1a8a8378974eee182df0bd54c658a7fd57c216e9f4b64d915c750897f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf6bbd3e9b76a1535c7947d1ba2d92765ee72526e2e1d065ccafb6ecfc9529f45d09130e95d620f4c4688a5855c8d085bc5ecd0afb68446f9c0a310213225662ff3e7dc2b110a61b5bba24341a9ec6c1307fbfaa449190e8458ed5abf2c250a4c5a98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f5b977bbb0e5c7c977362ee58a91bfae29c728ac16564b20154796d01ae293a8fc6f5d11939e15b871d06f39f1da1b27face91c47410c5a1e596ded969c6760130731ed46528a387e720a8134459199524baee1df3a25971220218b5037ee603248;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h526e84e34a8ea5ead71e29b52f8d859daa42a6aee7b22fa4d8319a5968f12819228a4c46f55fcbadd06f9add6cd073291b63d38619eda4a07dc4680295d7ecbf729a75017c176712817956cc7293645717ff8f8974d3f8303a4138b493d05fd5bd13;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5864ae4dd0539bc56e115637b5bef2f603b32615fe4aa273c40e70e44119fddac9d0b7e902491dfb541e9129b4053661d59abf25b6c6d290e718f41bd21c79a6bb9b06909d028e7991f500b98e1a24cbdf0f7642d1ced695287a893a36cc736e1297;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h11ebad0ea67c80ff92894d140826f557c29bbe0f84f32bf059f3ddae97733fc05b317a2b4503a6310caf0ada8d46b53ea41c7a96d9225662b1de8c7a23df3924184769f35eac1ac999dc7d15c2cb9b9a81cb8f8ff49e548fdab47e59ad059e4d9cf4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6b549850ad50f3f32b190d9919fac7f2c1ef32a0d9027e09afcf2e4fd91638f3b191d7a5e2416b65fd32b21f62622441ceb78d9fbdefa50a62eec7d4a62a6690cd48afc5100ad9c311066e5e9a5917f5ae8c804f0ceb164959c4b9a714322f881f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce779e31af544d368171dfac8b25e4969d78f756030055aefa7e6a1516006d136fa2ed349a07cdb59a8dd4caff964edd25c1094512d1e87b7266a40068524dc3fc3b4a7755726e25aff218c07f5bc7a4ec3e2e90f7b1b67e3d3ac88305fc06f9cc44;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84460cc3e3104c089398a8925d9928478e890a9d95057e4c168708bf34467bb4fb9f13643fac85fbb045863f649e06efbab03067f280736e00f4be7e240e05dce93fe1599dfcce596fbda0b25671613b586b43e686f665ea8744ea95d8ef8cb3fed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdc3b4fe1a0264c7a967cbb4b2eccdfd6273143d374ed569030219684a4ada19c7bbdaa8196f9bcee7621b55d34f260c3151089240622dd8623ba114015c58ba6f2fb407cf572853dddbc1c5fcad51a6eb2c2041ae1c5fdf9fe02816471e986aed786;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8815797a67d6fd5191854b8cda46733eb651a7e4085cb4ff95f3f517d5923a1d3e0f53993e5a2ae15233fbaf29b53bc859c12dfd03c3621683477c901c4eace4f92b4ac6a861a5369642c6a1795d26d3f5a245ba527b869a37bdf8dd9dc699b540ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31ee91edd08fe6f58caf5e3746ce9a8a971c98370db53ae1f743e1761bc5e37859e15222e96ee3f33b8d68a8994240680025e16de3a938546924a9025ab08779b2080e0efaaf68b84da03a22f15f0e29cdd95b49c16f0e45a2f96c06224586ed2215;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7bcf6ed901b18031295b360624551f7075ba00f461ac0eb6662ffd1aad281d6bfdc6595adacec338e5274e76669300f8ccc3423361f9d6602e48e2eae8ed5f5020586cae41b82330d39c19b8574439808edcae12abccda31bf3ce9b9995377139f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d06ece6401fea85fb95717c04d15d8b21be7f380de735d1cc316145aba6201fc3791233b997ee3e8bd851b0f9a50587234bd0190003039d64f0782d641da4a33fa7cfa4f53039add8671da113596f7f5a78fc7bdbac055d8e07a3192c0e3b693820;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f1f976cdde70595995052d97f161624f6390896564334726e1c88aec7a44d9c5db846cfcb001f3cc0e4115f7e808377d81f1029fd18fbbd53b0b1864d5537df3f985d1a366f8258fb9100ba5891e077c5c54e60a4c4ecf687a3a8e3682bffb4ef8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3804d68432b01c2ea902ed18c410a65ee7b81849f31a2f53b6caf40dfdffc7c640b2732e9799219bda3f35295218d54cd360f4fd765f145c21782edab14c511d5c0595f0a98fd91dab5209e43dce20c465a865d4a60b90ea18a8976b33cb82abc169;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h480c61c022e9f0e87d19f7e83fa8ce29956f6c1dd0b8f402ce097d92d5b6573bf389729574ae4c7cb9226bdf4932108b5a96402f320586fd93beb1f98ce74993abab60ae96d772485f2e267be7f242fb38f256e45c304e5e63cdbbd2393de54bdd06;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h936e5f8034c64ce1003d414028d65f542e96233d98cb7874a2b16e8e41ec585958b8a3ff2b5ccbd804a32003996752d456203d04fd7991692c7e6548f88722a4b957a9ec3d088c5229abaf38b7d19453db0fdf1548822444cec667268f311a710c1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf9578925c79c0cd71efcc49e4bfd20dd93f56deff7f387e9ae97fc220849c77cf1a4f96e4bf8371929dd1352f7533bac8bf9311a61e765338832da034cbaaccfd7e8f46c6c9eb05fc586cc47b40fa5e678e917b509ba27b0028fe6894414797b55d1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hddfdd57c11cb899250a5fe6bcaa6d72093f7915d86056c3bb6111c9691bb807a3afe74829a2a3adbce40f64ab4bdd1a6bcc06455bfd68226d112d47e9ec287b14f7f9289b9e3be9dc4118dfc3575766f91fe2d3b611a6ffc790361af7bd88fce3f78;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5841b1698adfc35e8f420c96a71245db9b8c49258b2f114d0a401ee8ce6d53a47ae3dab42b592d860911dee5edc04c13471600a34ab595ba442f3768801d4c00df6b6dc94555e2f4cbc63a10b797a2951fd10d84f09a531917f864a209faa1db4611;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6b0377dbd480d03098b33820b281f4ad115c26ffb0bd3cd8e7dcc8a946c0cc40b1545215f24a2a23b232b23e2b9b750ec564cc16145b59977a1243866841009d1813b038a54346aecb9849f8d7ea166ce45b1de8daa5046d83847812f1fcbb0dd0d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcfb114f84f997a8710eb176f60de7a4f52d6236087c22334b8793f2af6b2d66229acd591f2010405e91e02e1d547a63914758d118751d1678fdbdf3a1a5cff8eeb13d947e87a4c77fa4d88d79243ded0029036791c5b27e5b9fd690659a01a488b31;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcf4d7e1cef9d66b7659216491f7ec498a1dbb668ed9c1c8bda695706b5951930c872f99c8ff55c855da6d5646b6284ba5c8db1b9858e848b9d0beee7a4e4e5b8516d9d6a1812cacc4a7ea5d9672cae9fef884570931d907b70695f48f8e97b593987;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h827203f1a9b5245b46fa7086cace307cb7c2a403c2dcde309e55fa1372b0a567d83567e874c1e3f25475412c177b20da0bde7d4df2941dad8ba93b0a57176a30c27c2d34e345c2c7ae233381aa277f8d7ba3b6157643b277420273a98fdb8df50042;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4c7ac4a800c01174bd7757da19f86c20869eb333ebb22e8a3a8b4ee61bcc2e2abf979bc33a3ba6ef297fb9fc58b29a56b247f0d062dda70b5f65310ea0c4f4f278468946b288fbd770266d4d158900b6ceaebbe479f40448437f85f6c2ea6d7d291e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb431d749461246c138119f1ef2a1994ae0d601bc4acafeea8074054b0e6713561bb43f0c5bffd2da97b33bff7e118691bdab2ee34ea47e4637668a9fd09d66b03d3ba0b845440cf4040ba35bd41d0734e19fb119ef675d96e19d9fce27927767ef94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c107fd482287dd569953f3a6fa5e620ceeacf8e24a1e187a9d9309bd0ac0823f1c190e92a494a3fda2bb0827a08ccc0bcd296b34483a624f9fbe3340d876c87fa7cfdf9036874157d421fad7c296cf93a798a98ceb30dd44535138b0a56d80bf4e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h562f2974d75effb855ee0bbf9c18fd285505bda11400edbc72394ff614a94976e8c7896cdc3f68c08fefba34924f013b7554c1e198d1cf83a3afd1078df01582abe73f5ab87fee9d29d14fb3ba6c040740156373a3df88d0ec2e11affa8bea90d765;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha486b1833fb7a6322d8660729e4ee881597c5a2e1ccfc4b521ab4c64870dbfbbb8ed5ea444640cf95ff456f42aab12fc39520861e3bdd29f0b66b8429bf7d3a5b51b9803d48bf167fe58366ddb6b1062b06fb010ec9298e6d07660a0e4456ab2422;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94996c1299e5af735a4efaba55b450de618bc1f1dcda5895a2d2ac706fddfd9fbac83482c1192d9b106fb2d579050e2657cc305c67d25e23d6b917a3867bab818a0dd55170e71a13466927e5735c7feca6bd2a7e2b7458973fa55d2fd9dda94c6f03;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h800a75f4f039325341adabd068939a16d9a75fa5be71fab58e26d42235b548f898b5fa5b4c5f12f895a3e8ff145c1cf766cfcea809e88950068200d5e92561dc76ab5b2dbd45eb6870894492e00645ec0adb9c3fc50217f654f716cfd99d6c688331;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9cdf42da84479b85284e805abc7318ac3568a797e1533e4cd12fbabe645e04377624ae523286dbec0e340b5c42acc3843ba4cfb015ec7641dcc57582f03dcccc1b07321757e1ce6dc55bb40becb22eff8bb3f5118373b1e4dc61d778c8f091170126;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20289d002c2117f5c535a57b5ce1135cbf60ca8dda8c97dc91febde57beef23a2b48e6093fe94c414eaabf0a469a167757b4991aa034f8d2cf960ccd8503f8aad4d4f9a91ca472b1fad5f894c319a55ca169c0bc54e46dedeea268558284f722ba37;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79115e43427e6b6771340c006e2bdc11427a3f0c0fb3a221ef1ab7165bb1443167065dc852cb717508dc0af5dde0e79e7ba4c645c05c9e633e54b4cde00fbd47f0283a86d6e217411b20c6645863a60becd140b2cd6600a400795992997997d0cb09;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h785bef28777f5611a21836e35ae7626be7bd1c05ed90a30ffec5eaff9e1f9d74e6df755f93151d8cd5fbf980e30c2e6bad625bc3b86a2df02354842f52c61dd18b97c7c157c9b1b8d92774ecc102ac89d922f293185c64416e1a565243fa0b29dcaf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha2481177ba65c3e980abb4b9f9ecd25cb4b0415036ea57bba01c6b2354fa739ff546a0b26b26c97be7d56bad51906f9361f500a97163b81a7d4e8172103172a4d42110de8dc8c57531caa7936c0e04f464ca84c504acf74bf05d01d6a8e57c70871d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74e4cf6e3717fb5f857fa8c2932b6a5dcf940a243acffb0e41449edcbe4bbc65c233d95d087f0b197d7c6c9db233db0ac193f2109e4135195c867ae2e2ff5ee11799f8a6537ad0e9e44e002e1f71aec6e5291ef13831fdc9b8317564e93077304207;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44dc1c70d9a80c352cfbd56c818a1471f53d411779ad6c3ab2e00c428a7e6590d592dd425c5b28fd091c9a32e4d22109b56d5b170188c3ceacf9c694b28cbb1d294e7841527117630082a6ea02551adaef23bb1e9b99087c2e70c4615bb9fc64291f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h191e2331af6221e0cac5eb1ffba2de1af7cfd3547bf886bfe56c4ec1675c7379ef95f18209cbe8d9f9e43de6edcc89632b780ea7599d9b6d9d314a9011c8fc914da8a2682aa20e0b6a561a44338dad66943afa1e29b9f2ffd007be44007b7e70b5dc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h185a1a8bed7124541e7530fa7fd2eabfdcb498a7ad95ce1dc96e42afc297a2665f09afc6c0dce452f525baf85e3f75af8d1e99eb55bce5ab0bade5c346b21dd4804d2f85c05938940db818c1c626dc5af403dc45667ed48765de2fb1e5d7e8f33fd9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee8cda65e14bbf7a1fad4db528e2b3986b41d80a0ab830db99925ee74971c44ce21d75be605e3bba7b5dfbbbfd04bf338886d78d7de9d62656e2fa640dc3f284bb02913c888c421f5b43c82cd42f4529403c3aac8b7ee41377e81617c057fb367e60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc7bd87f1c2133bfb0d6ffd180abb368d0678daa2800be840cba777b33824783347ecb92bf5fa2f8c15b1a68ce24652c30ef96491e2c42cb239033a31273eab92a94c02bf791dc5d21617a535cf4549dea81923befad7c71edcf1dff9dc26ed8f042;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca9ca3e9cd1d2f3c86fc4b2262efabbc03401b3d1bcd7f8481ed8ed725060c48ba8225abb0e8242fe35654aeae2efa21f4135ffaa8b648aefd9a6ab7c44eb6dadfeda16f78eaafece0a213f4c8bf93db020adfe808462200555af0ea89f6a79b17c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf46bc918bd138596898786bccaede134c037cbd32e21ad8ca965bc9709b9ddab3fc514cc5fb7558749a854cb7e7f8f8a7e006a7e63f4c4e2aba927975ee2e0bed582f17e0ab749356418244ad2563834bf7938555a4f9dcd889f0a955e5dec24133e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h408306a7723962e3367dd45f32cbf800d0f1b317fb32716b4b0941c855b93cd2658d0e162c4a2367c4d4bb6bf177a261e68986297f2bd1a5de665e52824051f42aadbfa11eb3a6a3974e08dd38fd069729f82ac1dfb3e48ef4ce47960ed642d14806;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fbba599cdd862cf88b1c8c704c22c0c41e006cc0164cf2afadb6d4dbae3b86e1b4d060da1d65b388556b350d63755931d686b04395c05c9f191f6e7300cf10d1e204fcb6ac1bca942cf83de765dfcecf3932083f5f471b511072e690477f9268a4f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17d1194b872ec0bf3f30ee495ab73a7e5cfded403f9ab84a36a668e99d6946513719e5db28f934f9fff6aabd3d78aa33a709b61bcf64ab0d463af3175594c99454610b9fc3f246a6e8222d672aad0f2eb612b37f96f029ed6bd3a07afe32b44bf8a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h770c21e906348f33574a44168cfbd21c61d1ba74ddb12e90c7a27922c49bc70a5a6f1d924a9e82bce2f5a257e08f6aee79f0915c9721ce6eb809e41b7a2011de74dc42a51eb454bf7ba9a433847b220e93de41cebe4fa90bf19d2d83a05ee0212bdc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb9e26503fd917e7268de95e96ab373e58b6ec273de5b02517a5d6b778c081b321aa9ab20b16af61d6bba8dec8d3bdcf853b5c5ac671173305eea793e8e6399aeb97fea645247458e862031814bfa36c2ac29489774b226e25ca722a0a917e5a9dfa4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6e88fc42d04f391e218e90eaf10c5bf759d1e75eae90a6b2ea5f71fadb55844da86d8bf629b7f95f7b1e9ee5f9becb5e024dd138a2869a458d6f8050271ccd6fa98776fc0d15a97654b0a78db1470fee9c25808c9fa0485c0769532b4162aa8119a6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0542ec36d6fc8f0786d107f9eb813ecf8cb40abc6094c1e0de692e417c5ec965d653c06455f3467365a877bbe3bfe20e2bf06e57cdc105bbb319678852363ba070e8a157f37369376e8be5bc0dd888d33b2122295f5af29c9cefded8bec0157bba4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2681f99636bb09f650ef6a834e0accad3dbf29704d99ef3477dc138c2e2c62d1f73e69f97882bb2057fdcbc84c5d546f2675c09247b18836bd74d44c8d25e7d08b50054629c07c314b652823939b2b790438797df36fe210afdb8a218a89da15dcf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7cb7158238649fa167f2184138321c5b1cad753e568c82d83da5334fbd74fdc222275059acc04c251a41bffc38ad632683f222b058dde363a698c52bc993d4907bf2f119d4e4214f38a265debf1f7473515cb9c7c6c465dd19c15722f05fbb550e64;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a0c44f665716acb68f71700f66e71e669178be8aa0765302380921bb0a9ba89834818db2d2d61a6589125c3cb6ddbd732c3272e4d4ea51c01905174e27e972232a2bd329b5f456aa80cd8c893c5c2b358a74a451a3995e52bd10044a975dd0132e0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a37888eb7746759440bd11b6a085e0910178cdd59ffc8cad4d64154f48f017bed7af18fc569c6622eb67e3407835c435766e34647b275c81a351cba57014a702b2a8cecf8c4c2d8cf4be6f85e9e1043fb412328f4c8d18e73820d06e63e44d1b71d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18e2f3848467423bb5914b1af6aff2a010eacf3340d57100b56d7d424d1ab998423456050c584abf69d8a933a313ec889ece5d4a17532f6adb4db1fc070bf312f0faeb266d1c0266da91d4337fe8df53e614e508fe8e385f4548ddeeab7087b5b74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdac9c02c300351ae79185573f0fd2df40f10fc7a4a16cdac9f7974feb17590ae4702e136579ae76867405011fb8783e437507a11746809d7628ba6e4bfafc1c72519a1c6b63ee3bb659ac0881e47551853fb3aa2ef563b925a0434b065c1cbeeaef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40ad68dcf03b1ae26a2f8c8a2d2abbc7263b1923f1a6353aeb285653ef05178a654bc9d3c4a1c497016478c4bd1205c5c47c866251641e3ce02726ef0d9ad11fc2a9cc6010744ac31b9bfea075e642eb0c24835e5768ea34444c2b0e041324a3791;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h178260d3483192e8b424404fd4d6b3320e499c9ab080ee27c81dd053a8ddea7d2753dce80e342ffd6717ecf7d91b85496a6909f230cbbbfb7557c8b370ed12e7d1b681e8900b626de98fc4b9b0efad69b2fbceae81ae4617c4c07d7eb1e5adf13bbc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeb02bd900c9dc3a650f41cc5e1b027a4473b1ebc9bcee93957d3c8dea3e1aa1f1da794b5a028066386fb18d1ec85b10398e7dfd0b2ff24911dfa372bcb35647d6884be10b204bdf2c88053a6a1d4675dd6ba87304d031e1cc313daaebf1fb7398fb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb4ab34138385704b7936fefa57bbe2d1884ff9e0e8666ae3e2522fa4629baf1c879613c228d44b5c13f9c03f60494d29967644210f9b9ab7a8131dd603c6db2ea85af0ae05a9e58252690072b04251bf1569ded62776101eeae5b71d002b1121b242;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f96ee26029c7bb7aaf8adbc5867d0fac64eecbead282ec23decf83a3e87d4aca277a30a04c2dd3e3c633cd6ab9babb08bfefee7fcbfc3bddfcb2532155480cb42ce979d42ea20eebc7282ee1d86ea4de3f8e5987c409de50e348b3cc6c8cbe74a89;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13a185f4dc4799697c670b99627eb2ba5ee98f91f8de14b0c53e30b709d89e7b92e3c664fa5c478f66937325ee205395f2b71e507d642566dd6c852815c74ded50f30144a0a2ee49e5ab2b593ff499e6787ac1e0b2b94528e6c11aed8956d5a7216b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdeede7eccc57748a75e78da28aff0fc5665500d9bf30292cd5a7e78163d8806af56d604f5f8b6a3b7112b9ea562a9bc4ea7cf8b91eb193e708714dc2c9ce900e57c631fbe0a8d28b19863545743866197153cea2043d7c8b0dcd7f872efcb117e456;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h717503aa93bb638b82aaa7950194db074649b7fa81928da1394758316316eff716b570547acd603f33464a0d28149c5f609c0c92c3d91d97c326a08832a29dfc9894a5a0cae7b3e67eca7624a6ca054ce69a07abf67428b228e3a629fc8353d53fdf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76acf9ff7315cdfbda8291a28c08c016be24ffe3cbf7c7b4f5fe205f881675ab143572eeaa327bf67de05764c8f9e1a4c231fc0b0940ad8eeee35ab24f0a701b14bcff5385740912379903a417c8ab478398e7fca044ce70ef2ce72c5c8392c5490a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hae92b7c58e78f47f579f4cdaf6e5169c6ee93b7dd845149984b212a96313ee6f6bca0a217319d20f4b920b3f42de418f0699743a495e2f73b4a99a8f7b1bb0406643320f7d4ab21b4ef3f5a08367dc3d3dc1ec6b1452ca5fba6f16873d992900afe3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3cd259c6082a770fc238b347e335108b7c244bb8ef5de1137a100e5bcfeef8984c30f65f6f93d872be00a1a07f4a2b5b4755cab068fa0381cfc2474953c9888d8ae0452301198ab8bfb9789e1923f06b691fbf7cd7065773becdae051ef0ad3f0fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f8579fd9e067bb20d49a143f63c2c6ca4d60754ef6279d64dd77a8c2a9a30558b35a1b611d1282e3819a1b397e6e92ef0bc3c3ea6f366aa01358d96b7741d7e0ae2ce9bc215fd827ecba68681cddcf75390217eb1a58f902972b489577178f02913;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcdf0ef777f1d450d1b4d575a093156260d3429e7254438723cfc683108126012f6d785cb29ca802cc449c4247adbd4c3c52339323ab148641eacb4f6e666410e229e0830a217f8e35ec9324259d9b0595071985de1c74726ca190c43d27ad3461888;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8478fe3b85f4f6d84fe7dc299806680b55558a3a00de045e6af1937ce2285c05e4ee2e5709cbe2c889cc25f5be15627fd5617ac766cbc6bf9dbf5b73c23753e6f3882cbd92687112b2db4a957b03442bfb9c28389cbb7ce02a35a36cf225988838f4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc19ce1b75c17dc463f30ab211a97660a18e906810fbdc4862d38735d3b165935a032ea37144230af4fbd45fa8676d533f33557bff6de40dceb413022fe446c88f458d2c3831d77fd25a17c3ee24a32463befcfd3a7d021a0b620b6b5e4019ec2cdec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b9a08cc8548be6b0a599cac28e2dd7c18c0f0ba3d8577e9cca470eed9606122b36af43dd3b816f21524b8bb062d9380b1a9c92472e47953c5729388bbba6b7704c3ca40b620aa7a498234e357a7b6402f1dfc8a9d9d22979baa03936fa0bcf072f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc2153e5d7ebdfad467684315c416050fb8fecea5be1dbd769276e948aec85ee68c506446a0fff4477a6369c939e94d2bac2fb29ff9dcbe25dc9f256b158a621737c136e899ee3b892f5739962f71384b97761229e91b4a3ab1b03497ebe3d6aa8622;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habf35e5268b05b625fbb095f673439026391b24a4fbe4db9237583c62710516c6bcd4049bb2ddd61b811290d30013d360d2fe74860ea0f70efb7380f115b9664693e1db1120fb450837d6a7518277cb2e322c3575b48dde4629c9df198584a028139;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd804e04c15dd66bdfe630c7be3319fe687aef43eed9c92e8dc173271758ea9b24c142cb35fb98121f9ddae0efff44f30a9459d2bc50b4875e031d7622fe9a60bdf18181387af9a467d62dbdfede0aa944f09273f031dbd02f8e3d548e2de92abbd5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h293759cea3bc01070fb58743ece194763e948a60ef70297d0c08c1a62ba5a20299fde82bd14f40282e31aba52d8ae33748eaee1100312e1c25062ccf5bcbdf6286722a0b84b6ea1bbc61c5be7b2bbc34bc343826b3012116161ce43708b36781531e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2ccd111f00c4e7e25d29dcce57d71aca343727ecfb0958c02c1d2642f2cc945857451da8bc6b7f899a5e3915a5ff90dc94743abe05eb0bf8f8296d4b94c4447f2daf4009a81a10269af3da809034adf9c729e63bcc3262c1c3a2d01d97ef9a1e305;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6bd2bb13c6fbbb42b95dc3d8f98fe77cc4fd056666a3dc6c1d9c2fb47dcef0890bd34ba9ceed71983f6b5bbb3f1d29a422b78bef6f2aa4bb64de5661bfe4e5186f40d57fd697d5ba68aa2f9e0ed27f25e5c4043c990e23c70f9e825d58b81636afb9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h94a90c6df3a62af0eb784f8fe37804814e46d93d61e0ba0da449a51de11a972c7f3525e062de3cf48198314224806697fa82b0b97098d9b9f864f4cc623b05cd9d659bd72c549be515853b2fe4e2d8c0bbcdbaddea10d7c7ca7ba9f4b45d5cb0f429;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h56362f5786285af4aaac52624bb90a2884b6d5df15ed8914f3c0c729cd3b45deca62afcc92d7ccee81f86148d9622bd675798d8ee10b19cae31bd1960c51652c6dacaf51604833c3638a3d0bea70fa49867eb535c43d0721e84b2d3684371eb3f5bb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha09283e91aeec9274354b7ef89073d25c95ca08ec134476af1f31986c3aed7b27c92d71a749bb5cd8569f2871132b5f34cc294e6a87c2dcaf97a4503138f07a93421993701b25feef2a028a0d2fc4aa5745b8df6c60c258c5475a8e4dc40de26a634;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h631fe7d38faa61a082f86161d11f9a4af50cc1e63efc50cb8eff8ef65df416450cd0fba201f2f9dc251f15801b5f67964517fbab4a5b68ba461d7f9bb4bf15a378976436741e4188141bfe43e04e4f7e9d1f48e165f5874f18912007c4cf62bda438;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a0c481e8a93bea895caf72116abfe2db3fceda65cdf4936b310a28195548bdeff2367ce317f6dffad4c591078f7d0edaebcd6ca558252c0a6c4b441b5a565af1f30229ad41c3ad4863ee9351509c98fddfc56716e919b4bcae614614631f236a9bc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3541b454eb578b6488f33ce2efd6bdce92146968cb4dd3907c2ccfbfe4be07dfc58c74b256cbabdcdca52eddb0fcd2608d41474aaa2cbd8149e753e89beffea4b57471c0a3adee3ce2dea557c718d132e785a554c567debd315b8f7f3aa5af9900;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hff1074bfd7edd4d0aa2b614bf715aebce2ada86b43369eab7ebbedb76aa13a607148e5102c251dc2356869adbecac435d9fa167ad929433d0516fa8c76708df89a2910213a80b8935673163f9a1538a1d408d08e1117f8407ad514eb7b6ddaf16aea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50cad3c63e270baef3d7765ddb729bd6c45e4c073d3e3e7ef478b4692c2b9cebae81129befa0245cc889f0e5ef461a69e4c21b0da410dda3a918af62e3f8c38ebc9a7c93edafc875f47ee2a465571258e9fae19833b82d3114468921e000d87e3a12;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8fb69ff920cf2faaf6ae01306a558f14b38ec6f395954ecb102131fc2667c74e96f3f909b7b88363e88d565b3b589ec68e78570c8f01ebe1e94e5c64eaf4bffba5287d58fec31496526573d3d3b10635f04b3f858b164e8d4ea276b84124ba0f8ef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36199b8f535c0f64a7c885312ee2c127f9b299cc932150ee929e213d7e483e13b4bd886cb804c3b51219cef896c9c6c908c0e8638d4e9be039c9d00adc68432a6d6da8fe6fd0c118acb297eed9fe451a69d96a310098f3f616c1268ddd99000fe4f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf991dd862aeccf169315783ef09ee4bc704c9b9597d9f33d2210b3cf8ebb70b2955aa8ba505cae7b07ea043783d918f0398d08cd52ac59fb20b811d884dedd4f4ec936f1ada0c2123fa6a8600cd1fa7166feefa3ce59ae36091193b0b6d53075ea7e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a4a65b061ddaa4b14c49ad291f66697ba4eb12f2216d3f906aa24bdd7f3142181fb32cdd4f4cc1e2b4711c45c24eb7f1cdb3a91684f9b35db00e29903fd4f28a9d498f42ddb3ec0e5c538b3344bd18caa15d638aab25840bad38f34068b5ca168c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a2aaf37f30629415870fdbfe3740dd0d2f5c6698565b1886704cd45d8002d7564dbbff0bc1903f25076ece96f78d523c5d517de704a823916752b54f84deca365dda6c826703a3c978f639000ba124162ade4721569b792f7cbf6d80ca0528d98f9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba2ea1ccffa6d38e88d06dd85b36e0a6578c8b936d123919d01d5f19d6ee52950fc80535b6505a6f89c7c1fb96de6d88e0fe3c6520db73d1481009c5feb47e5a4f11659b283f6d08f376dcc2549ab9dc8b4d87ed718b7104e9ba8c1d3ecd38d29dee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1de81515e2562fa26348c8c3d6663dfc061e3f55ba48328b7c1867c0bd1ac804b13cc78b9869b52d79628b438e39dde46e7e885705e36c80adcf6311ba91e678b270dd2fa190218cea1ab18d43043e5f5c341cc217c9927f033732c5b77d1fc3ec55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hea5c14df98efae06c867abd4bca23170368f7ddf2ed5e309af321e6dce97a60b6996b1de470582e6aacb1206e2cd98bd0b6f9fa31bf3683c7d4e94a3cc651f0a41fa47dbbb36a3307c9f2e4e5a9093538e7a166b79b6860004dac2a56f2d529dec3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd514054336450694d519158954af2480ca7f2f3e31f9b418b5ff7dbd5e40fd0ed7b97d136f9c95eb77b292832b072136e744136578d122e92280ea9a37acb49beb2760475dd0c4e23a76be1986dc7f37c91e4fecff0b80837f53e4ab324742dffa2d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6054b425034bacc3c3f2c8477e5549f8e4e218143f3b8472664eb1ac813dfb1bcb8d53eb88c86d6407551c3d73eebaf0d3a33c2218120475a1e4cdf74878d14819e94a0ddb5623657f773466aeb038ed9b693d23ec4da8ba099cda5dbf3a0b4a904;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd21678928138497f8086ccf393680211e4e4dd7fa21799081c7adaad53466e4f397f66b2bb14bf0db4d45f266c97876b2826192893d241ce448659989445065c5152e97d004362315b24a49d15c775f1cef51095999b0cb7f6b13e45198921cbb38f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcad1476064243d3be570bd0b09fe5ff059dec7db1dafe3f4d86b209c3428e2de574c23ac0db1e87f0f207ea6d06418d2a50956a407bc966fb99fbef5f7b5e8da437105eda3cb7940d9ce166e1736a9249b37221306a54f55e74929772e82f700fc40;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6c15c9f8242789f99c4f8fc8438e9603aa3c0a19f54697b75798fb2d6ad689febe9e69aeba2d0b65c57fac50ab5b01727ef6cec74bf4faa289b4c3c5c5b13e3e335aba2aa40d7143b3d1cee89c079bf188bfce042300ec3ee0f350708544586653a4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55de931afc0da33342faa42d3edc2619d6e7097aaf45800aacfd18175facc7cb9e06c1b099313a2277ba1b87f77bc4c6ed633a005473d2684f1cfdd8e60c3deb722ed4ddd877df35bd953af4af1814d3d71b32cec11a24cc5a40c2472e5a1b50fb8b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haefb9b1dbd94ac6790086d49074070e1b7228d59a803e96095cea2be073536acf9859a112bd8db64a969552666dd4013ad0ef4082e3930449f2e45ff7320c9b90660a848357e7b276971f420672139bbc28ebb0cd83d7e330f9f08c940eb238ce8a4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b5ce9dd700ec9e14f0245fb8d299d35a609fdb3578df4fe5f0c8b9ee25bee87aff7cff3f0d60096aef75e88cc19edde01cb8ad337fe16f324663080653f968cb80d12ed5d9f284049c4cab2c372c3ab30e252d2138e0883302d7b708c32f5d5aa1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a1857a97e4f5c5ff6cc89c29455bc29394ea266298fb6d114dfe1f20ca05c0bb7058425f8a897f37392039bdab8e28d4d27ef18ec822381212a59d387c9fca2260f9aca7cb5e4820cf0c4b7df3e3b0490be3224b9e68c7aae3d1b4f0fb1c5a4bd83;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h648e517f73c7b6bb7fd2896830cb915ddc89fa3bb4fbc87527c9fca62d01ce03ad45b5097763d32e94d8615568baaab854dbbdb7160eae9f5039e01a1934255ddc395dfa51ae089d21a296929c1f08e644f609f237d7c658f3d9dca771a155748449;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5c5ada3598aac549d088a7be0ef12070a8da72f868ed767e180ccb6b54a2985897709c41dafaa06f3210592f69c4617810a0c8f046c59ee6eb95e8e36d74db9abaa8336c9017b9a07f5220f2801c3843a3c0b830391d170398cf48d7c6f15994e455;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83d9e6905033eeedcd6a53d435a48f2367a879dc0460f96ecc13678c399743d97ac808377ad09822650fb92077ce7bbfe0b47cb1d415363475f3646e7ddcab15274076ad04d4ad1b97c641b347ef5ff7e975c79318792085bd0cefb036d980315b2b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b6b7fd2a528a2a4921d512e11d201303982cdae9aac51c322d0f6d9d0c92a699db9f72716bfd67f98938cc53ef75c9d4485deca273eb0e19967d8a04f8a99ffb4d920d45734a49cd38ea6baf9857e24d012fc3248c5d8f3840edcf400b87c3b558f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f9df98aa948847a5cb16a80d22f6f2e9f335572b32b795006e0a8cc04b5d0b857005514f5dee1152992e37602a81c65bfc61d43d3c6417cfee58bd21b80ff0b1e0674f7f07e71b1fb7febf69304be7a93f8dc89f5f72654e4b74da6d752ac15ed2f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d89eacabec86fb9885b8b1a4f68767cddb53aab4ca736901cca805340fdec1d612a8366a3cf393835f0f8d1d1838db23a529d2d7386a27432bcb1f26e91d8901ae59d57db98d11da8f4f653c85085cf16552ece3960f09d9100f920970a6af0ae5d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h547b5eb464555ed492fc9da7d0344f4874f34ee9584508a255f101350bf5bc6a5b234209471fc6d461c01589dfd3ddbdb584436b44a150d2c0872a77485430c237423ea250269b882d4fd86210c85a1bf95fd14dcc52f0a8613b30420afc881bbeb5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f7a96b8798b7af21456aeb224374b816786c1bfc0c2bc96dbfbd3c8336d8548be73f45836bee280ffccdfa4c291dd247ca31442756091967f0858161fb69b7148c5f96ca79f4310470814dd61427877f75a854a29b2a7952f1862314fcb0a544e58;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6457925bbe7d21ac2c58fbdc30cff036cf5e87ce6fb80ba6c966c09aca4988830447850c56e3b71ceb5227bb217ff4e944f2847797a45d57de839961d5f9fd9047ba5054b09e39da1e0741abc72b1a90ff69872b50ae08a536ccca47064ffe11449e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5772642f90a32e739c052cfcdf6889f1fa58fe5ff2d53b178f0162de2497419f80597b9b9ec92815ba93ed0260f0ae7468c91ef9294f16336e83f1d0e89a772666ab40bab6108f1b0bded003dc0d6f99e6547abf3ddb8d24040badbbda7782746eb3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5b23a6be77b29fe228fa11bf1da3748dec4978e75b5b342210782c2e2979998441701da74b2bd1aec0d4d82a9e72043747c11217cb99c82662715c2dc6b21ac5f037ddd9d63217a0c90b1dfd75b0cf2c8f80eeb77b0d2dfc49ca6dc92a3fd7e4bd19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4679cf0a504e486ec4f104a538eaad3104866d1bec97e19470f0f2ed97544791503eebe0853b9ca2194d9d596d826d8ea635e2c9f4829abc005283f5ddce1b27849e4e1769af262c23411e1911291b570bd6a658e5e7819c10dc7f14ee2b99fa847e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe9bf3bc90ac96688fad9a88bc0054d1984e292b198efc48c468845fd63099d445eec3da82a7b35dd9fd43ebfd1523cbdfc3fe2e617700e7856fef2f0e306644081c3cf1f8ee2356cbf6959f03681e1798f3bf0524e27a736cc1579b96df016f4b03;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e9f132c914681c072f8683ba4d2a493191f3e9c055fefca98ce59d20c6e3effdba727a75d1c938c50ac389b6e13d9c3aba150c807a246568a9b34efbbbcb090c70c36438f954e88a81fbd7cc110eb54488ea7837cc00035fdaa243f06138b1fed8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc0413c23aae917bf400229dd68d75d7cab77346fa1458314b92d01719fb1269c66abc8610a78077c47127a92f48ba1aa86a7654ba927af4bf87fcfb4d261446f86fe5184ed6dc880fd3cd50ad1454333a41ab411ebaf9f8a7756526be02bbc2dd92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h796f2439fb85eb1c20546b0e886d444d1a5d86d02d718007f9755cf9febc332b12af2d71c32622f844c88cf0299d6f025ae077d733eb7058e33ea4b142d0b57e4ee78c36f594b52ddd548d8bfa5f4954af02f655e40ac4ecad6b11d2a67454bfe95b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd859f879f1c0965f74029c792c178866ac39b12eb4882d7dce359e677b63982c7a54ce6a2c0dd935b6c7895501938efdb8d36be009ca67cfbc09d7330fd28a91e99cbbf94956d26c4246c315b2552a34bcddc315d01fad59fcd5008204191713c76;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc55be3d41150816832ed6eaa3f188ba40f589874baef75a0948762563f889edc140772a9e0ee1708848bbb402fb4caadb9da49f49857ff533966b882c8af939efdd9a3b2c8a4fdf75eb01933ad4bbab4332365d9a16233e6cbca0643be83bba27e6e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8dd7cdc1fa8abce805b337350689af6bc8730965e11f9141857a7ef6d31123eac04264cd0474b0bbcf4f1f9ab89069ee1fa089323da615da3157df695917893f8f0dbf4547640feb9bf0e58fc93dd661e7735fd7e24b08ba26cec316c0e2b12f0a18;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6abd1e99ed6eec716cf1b976b9ed4c01947cc9598006c97c7169f0cdcb93d702ebf200eb3ca3bb847dee062c19f64243c736b01a64701a178e840cb93f5877b4bebd8759432a8813434240b76a56f858fbd34dd3a6a1a901365ed8191b8fd89042b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h231ad2c1916450e361b3d0fa0bae53a2ce6ae70397068aec66471153ff7bd4ac1e141e76511589785e54ffff6b20715431d1d7e3a17f9810a20184ef5f5fb4ed954aa14c7bd860fc6e42b32685516757c2cbe56478ff67ac6d94a4b5f7552291e0ea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5fc6339d788375ffd3785a3edbf3c22417320613f8f1b410a429fc1ee1618596fcdc95259b242d98e9c23d38febe859ad160707c0e24ba3420e7f5571f807834574016ba9843100acf37d60c23d93c8b7ad37ae91df32028289e63336a4806167c54;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4552ebb91e36a226880d78c7558475431c766b6534323c4eafbcd27cc3a92d71135e8ee830cc2099a6616157dd02340ea44bf73317923c1183251db82b25cfce8143d79ca05fb7948862ddc68597d879c25cc068c6e101d09b0f14698160b304ea4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f09e20106095b5cb45e4ad40c31815639a6e9de923c52c12f90d13ebef7e5010ee4adc1251d26691ba3b6b1594429d7aaf6d9964bcbb1042ef2cf0bda063fc9baf3251e20cb498667dce66bd2d018955f7ea8b3d2e38212c64bd831109e6e13915f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21d84bffffd33ba6ab99f3983270157cd01e84b5b3bedff2150c0117d3ce81fa45170d9b40d55a52b40c25d37774a14928572172d80ca220f5feb3782cbab578f66a3dabce61d1e04a28778f49a0a5defeb70564f47c6b45444479da12352bbf43f0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbbd8eade93c1c8e4c42998afee0c6438f060cf4dad2d42a2a1aa88cd5910d72a68fd5239d202bd5da297a0bad1c11559e60fd1c1e52341ac2fc2d7f4740861f52c62345562b08ccb64e34f58dd1955ef68559a349f7bbdea80462c9a2f0cdb939aed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3154afabb00be3f614cefb8ccc10a3d8a89f5e9423ade6948588555d92461b472da2851fd93aa6c6e2f26812bf059d2cf78f4d087984795bcdb35ceae71f84cae600fb252759e46ea437b179cf55c5f4d43ec479d034b7f85dc2f6dcff044017d78b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h15380b4300b7e5e18f7770f50dbcdddc8d0637f1521ab140bf08844d941190db25bcc9eb33d1b6a57efeb3ca8822fcb29ea8b713c28206b3c6eaed27c83f71fda76b49e40360671a7addfbf20d2ea05817e074994b5cd3c80772edfe587021362a92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h933e12269e98658b9e8ba20795b16d6126e687fb7f7d80ed0ad0350342328666ec05dea78f6ac08ce0c371bfd7cbb122aaf0ee728b5909939c28f8ad8c8c848c6aea4af2e24ad8fc84563c93e98c98d7360ae1121f686f9d37732cfbdb309e7a13b1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29dca5d55e4bb8ee052273f080dce5de5f3610f1c36cd9c5b031901e00379713e4d94dc982d7b8721f8a5aa1fd681dc08f145cec5e22f5f400f4d2783289835c7e535fcfcbc8d119dd8bcb0a3ed31808df0f60b59a5c7517d82cd9971c28d5d05208;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba48887b7002d501d990455d78cdd8da5bc9066b6d1b982482abfdec60b698ca250f67acca243f7eaac31ff8575367782f96c1dc4ca94ba26c228cb577281b3b343b24e198b4c35321c18418a008472d551897b6531daa368244f42f864d16c9a39d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd262db6253bdfcbc7ddb927a7e479793cadfa299f7a7dac4ec658f8116dde795bee2343971e4f970d9834fece84ef414c87e62b4a0fff8c22e4839fe45e428ac8d434890c5266c5a354635f716da23004b399867356b945562a897f83685fa787564;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21dd24dfa2fae6e0fc7f34ba64892a89632a6f0a981388f9aad14c00ad9c23f6f5616598e5e9e9cee6adfa5fbe87c036303b9cfcdac08a3e4f9d5e9670bc969e35fe88134b39decb1d22e4b585400d6fb05963a8b35138981fffca162aff029d1c75;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha4f159ab9bb413bdf465ad260970ecf9ca9c1e41b3eb1e6b793c7c84062e5b47fd22b4e72ae98fbf82ddf83f981b0a3f9cd634f5b95879a9e97dbd4a0f7413fbcd256550c9859d19f3f30fa399b3a968accb654c7bd96594fe3326827c1ddba4b195;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b3592ad74a7d4df58d2415211cc1cb4776f60d2db1d5836371376e10a47d12951d74aba405e3092f07396bc470ced6d8c899c98045101517955f70de63c1d8340c4501717f4e37c7e375b96827dbb9c594124426a4fffe1ba4c9682a81a936bb3e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf5fcd99977e1c43852bf718c870e745706509f4de33f74d8c9a82107ab8c9d6e8c12d5800c71e4f3e246271a5010cd6dfa48048562c33a1f2cc4ed16cbd4e08fc3be4d127b03df238f0fe40507830991f966b5b8e0273eb839dc05fd3f3238fc7575;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91027e5a73ce15bcb7753cbe0f1c49c5aeb4524d6c2e90cbf529a3e42cdbed45944e649037515a4190be8c60fe0f036244781e901b7c31125de07dd63a6bff2a81c5e5cad376bba1214c5ac2e3785347013c9e31eb16a7a5b04c10b87de56e073e01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb2babea35e4b72390ac3febff633d1c838d051c651e6cdbb9ecb381243273da40627015ee91b30182bab2e909d644c1edb49ba791ebab12239d94d3b2d24932d03c224b330a32ebb026c0a9cdcdab6ee4bfcdfd18aab7399d859c12409bd9fba202c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18610c5dd76a072d122a56051e6ca614599b90371fc9b8d9df25e3f1f2a5a4faa5745e6c188a2b42de7dd4cc6c4f5f1c959ce439a628d14e5cca03ca794289e110bff0816a0052ebb2b136ee3a3d8c7aef603e1a3593f0cba0ae920d834ed71da88b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h90e5a5d11ec022ab54c9aac2a93aead11c29332fb65e5fd9c160d412b86cd778dde451c456346740598719677da763798778447123934c3fc9254f622592c9bc5c8e12a492672dcb77aadb83d2f383c2cd6271b37eb9ca0e8d332d358baab9f1b93c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcee5625b2fbc581cda873da106966a6edf2be4433301dbf9eb58aa8f0329ec57b8ad766d1779f8e901def9b7b75ef002e900e3ffa692f8028dea942f374912dffa3b804fff025056d83f8b80498dda76eced35aa853356d297e114ddfc7cd0a23a58;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'habf48648854b6d6a25176311484aa228266310da666ef3d164969bb4ff25802d5638842587763fca1a2316d428a6f03de974cd7118e70d46f9cd6488d622d59df42291336d0af52c4adda0ea5e818fa4e078158e1d2ab4b6b4bca35c882e4b962aa4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ed34bd5609e878deb9158633ac7c6f607ac792814b8dbfc19a793516219710cb65bf3588466c23d2e467977379120f39894156fb7e324b794312f94ae011a4e043ee983348e610ddee96c65e3bd0dd7a6be6a7a2d77810c825e6b4f6031eed3d6c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72776678751b9cc702fbf3a271a086da9a1a5f17fc64dfb1524f1d6924d7fa66fe99495a7d0c6e695349b2a759cd3b0d72bffc492beec5a0b3a7e306b9cb5d41e936a5fb035224b46592db5ffb53714b926222b177e128fd8a3d6d0a9818e116df5a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd55b8492c6b77f22fafcdc181ed9f2783bef7618793dd35ca400cdb6c14a615920cb43dd1732feb59946dc293f0138a71a85fe9451b011f22be7b91179b84543ab703c2f7119f6e377fcb7994b7ac8f759b1d8d2b3486c09ed654e4b1e0488d44d4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h74fb9c6e0e5f9aaf0237613efeb186679f91168d74313f43ad27cb24811ef3fdf4996cc34c6d22d613490971832918f97204b694f3e4f44bf1ccaa1240fdb67afd48cbbac6d070e8368e6d08dad568f2e7acd03573824a5e669e167f2a3b45337aca;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb7a8e8603cc82176dee0258423101658a489e7460dce764d178de93512a2cb716f19c2d51197aa4955b2b27de044c06da256520a1d3cca36227f775aec3f58958543319a43427bc9844b71e8f32016b9b2c2ec233efe92e5a4e8f0a44da8bec3ac1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h311f0b498ab0ca52c6c92d249aea35d1c0ac15fc3766e4f40ac34942f74f471740e226b2c68815f7f1299188df859566b3115dd5d32531197c7e3618bde35cd57309f3c8af99b1e3f76542185f4726f189d48e165e5f5d8d7e06ad465c03dc086b8a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1e19b565da2d788a6c39f9ca47d4c186db9801b257de672379149ec68fd80f8ea63b61e1590d441b46a63b91cb8b2a40450e21b1944e804e0d1f3b7669f989ed07913c8d143ab39b340bcc3013133271806fe9d2f2813c512d3636af52a7566e0752;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d4e3ca47a38e5a4dbf6e72315d4ba33f36c45715ef3cf34fc3e637926c170211de8f24fc700419dc1fdac4f86c3353ba239859779a8dad51e1d2f6b868f43ca80d5520fb84bc20a799a89c664c119186376a02341ea16c5aba3b81883aebf0fc81e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ab74f8d20838c51825520792dc6c70548f4077dbc2b9f787fa29e9625a7ed12392b07e2fd588e9568822246c68f3346502d3c8455e40aad2865222ef41f5c3f40573b0f169d99b02343d295c944176d9cec34e6a98d1ad67b35e125fb8aabb1ffa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6345193225ae367c3c38b19e9d9be7846fe5abf66b0a1999612c4834d4063cc6173447836811c1f34338d44b1be20ea15fbe97ed6dcc5a2319b2688f3e59872bfe15bb14c8b8938fa52fc9f730edaf6dc97186122293c114ee3f5bedb02eff3973ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2ff80b5a41045117c6a7e90f73489157c5985d505addec62453700d777a83d3c17ba6e616c83376de39f5f6fb34eb51602bb5508894619813e00b30a47ecfa51af1f591ad2a6fcec67c8fdfcfba2d9ccac6a3f104069271b0135692ebff3c3d22169;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38c68ffca2f399648998e9b55add49b890d7e51a32c25cef537c9a6f0f3701b3addd209bc886ac5cd1c065c2e67f6a04872413b4807bffe36c654b94be824c025b4ad95b164c59aa7c2ae3ac6c089de3eb8c931c29407d65c6883e039b127f3a4ba2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h130f9b19972d3dcb56a3b37b8ee49dd2b233d4718e6d96dfd7711296c6a3fd84ae1a64c37aabe9c80df8d66be51ea48d9ab3960938a3822b4182c7dedced93dd69f7a88254ac1d8f6c9d4131add822145e22a744f9e566348f6c575d770fc44a135c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6f6d1178bccaf35ae6fd43476672d2d2b0da78937f43ce20351ca72312ae9950cd2009939994a5a3386a227e4f446211bfd61bc64c3109d6a12578eb97c64bb0ab8268beb08eddb14ee78ca88f9859ab64e02e96a8edbd52995ca5ebc249eab79689;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8814c2601fca8e5c534d93422085b2e429f400f15d81a057ef14193e76bee00052b6c09412fe7b2cbf6e0c0195d95a68bc17d002ad80bc94932eba7c9782cbf2b596887029f02a9db5e6be325b0488c8115b8934a193085181f7cd634f57ffea6602;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc20513657a8da0898847de9e7c1caed5db293d51eefba443d033ee3a51566db26dfdd7d4878f35589a049df6571f1c235d9bfa33f77e54808034b313688890dd3d477d4185f4ddfca5a116674af31bb74f964b4d59abcf97ff83fbb33f78f221d19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc997d12076a87cac030da57c12ea62eb3b935add91da9a8b3da06a192e845fc97b8bdf597fcc5e8573186fe1aa07aef745f14965264e62d891a091aaf98b6a55be752ec191ed97a05b119c6e30f98fbfffaf201e4280660c5cf6ed5d255dad3b16d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79246fb1bda73ed090b881474dca6e6f0ad1d0ee8aa0cfa7b8bf24c4031aad598d7d8c201eb77aa5156fb1241d86e996db54bcdd5ad25e633e17a1aeefe7d8386cf77668232dbfc593b7e696ff407b5b1e2820d25d20a1eebeb389b45fd652d91c7d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h882accc7453b5a1f17915b9ff8ce544fcc622d3f8ba7dc27346b7a4071ffb1346f22267383804970e19197c4401d26564e3acd508a5c4057d10c67315c77382d1114450e72660cbec9404c4170120f6ef71bed47d66c048c62921d788cfa2284ba02;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h895e6fef03698ad15c1fea2e5af2f9a68a6a581024aa7ec9fb8e342b03f6b743828719a0334ff872a215cf35aef3996c2b18c0cf6e0577811c2df4264c8bbe48356bf4ff5e9fea1f6f8a624ee9e199ad5846c4a87d433b29399d87f52cd5b5374072;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h31fe174fb65bc52c7f1d45d4e5e9efbc9742bf8a163f149be138894cd31057f63d61ec375189af76a693d2f077f4c691cf3c27ef2aa8c8d253c804aecc26596fcf498a155ee3c47e99fddd5a22de744ad0b8a5b64568de302d730d4ab151d938b5da;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb34ed9c92371e462edc29c3fa603c4d3b95b3ee47f59fe79128d947e3a88af2bee108745a04736bdb3380e7761c68945a439eb7472ba2576005a93390c432b05019c5998d6d550204d360ba8b041ca98ecc279cac094c92d66ce6808cbbf137891c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfd3383f5a06aa1e78e03683035cebff09c62cd4a460077ec9ef68f172749763d622db6a5f789d40fe50caba5e4db1c0f3b1363cb0f9a86ca1690aa3a9d6ba84840d74b6e06b7fc18393864996b26d41d035daf766fe6294ad973d4f83a76fdbdc193;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfc2d46fb4fab6ccfd54514c54cd8e35ae3c0c37a1a695919d5da01dfed40fdfeda2daf91e5dffc06c50d2356c5b01f72201453077ebbd0dd52a618f1104ef27bb23599dbf95bd53da7ad5dec3200810830fb2861d687df54d3bd92839e433911621b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h18f687c6a420487a5122763051bae720524f1de4a785c5da35dc30d75dce3b6e0e273d06dd69a767655cdf3ac4ff8f15cd2bce52000dd890dd8e2c1956feba7ecd78b0f00057abb51e5b563cf3c79d37340d175b619c5e089bf170d2eda26bd8bd62;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha8fad28f5259ce0a848066edb683e4fcc6202a94b08fae271fe48211dacea87392a2787066033e7d1f6dfa83ae186a6da946980b11acacc0a398c567dbf56a9d3b0b9621b7d21dca15c0ad890af5f19b98330bab87f03ca84fb1dfc731ed9b0f79c8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21fca6ec30702de35b92a1ef5bb0a5ecbb2e88cc1d529a0d2d5e41385bc9b495480cc759e8ea61c5ecac27212feb194ba71358cd7e5eb54f0e647718f8d99c96242fbd900314971318849d1b28d43809cc9532a80088b6310a6f810f25658926ed33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a99b80fc15d801fa19b4832ec74b5a1e95482b6848b8a2e8ac5eeaf91521db86e817945fbab98ba4e373d55783650a41a133a64d3e589e57e09fdc352dfe5ee925eba55641dc544c004679f84bc9a8432a0e82db25954f077503feb6f2cc551096b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d0e46909bd66e9ad439672dd708662cb6656e26e2337b59a2cc984bc21c89e986d1d546b2901063fb6bcf55812c059ea153d6cb8688024d057cd77cda0d9b0cf1ee94450f64abeba6e70aeff50298cb5b1acbd20d3d2345c0f32b9a30b59d4c4e2b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha85452e7ba5fd8e11f7a6df05fa1d92a599ede19b84da42d3d6e73efffe094a4f80d44f1424857ac51d81d1a2d86f7c28e0ddd9049836618c87d2e80770ed3b7f49f13a97b55b7e8c0bba23bb3fc3121e6982d4997f603b104513b0bce0a495a305c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h858fca28de4f417eed1b80d9a539edc76ecfd500de088282309b1cdd96d2000785a002d7154f2fec9c1708d35e7084571b8377f9d0fb77e2bb88fc54c134df52ab78e6fbe2d630cbc42d9098d8e23a810f2e35bc6691dadd6ab0f52021795611a3d8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h352ecbf4fb7ef0db3b10f51908c87e0a1cb0d6e71eed573270078ea90cfa62bc0d4cfaa2d96d34de0a37cc6442a36fd7687bd843253881e3d6dc7b1138e0fee11a5bd5f2c6be247de2c000e796ac8525539dee6f0e21cea6ff77e0d54cefe7dcf713;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3e820e4572c8ff81a01a5e196966083bf3434e9aa658dae0006f774b8821edbfc40cd25ca79e2d81fb501063dd1cec57ef4a6b16f182d6f2760e03d2f8a67aa51700f296489cb031ae12279b0751c067de9f6e1e4045645bfd1e305d2a66919a4fb2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf744ef2fa499c8017520e219f790d6128718e3162ec67c81b6e7f2f7e0f167c8a3e330fa465bce4a6873542b2066076cf0573d87a994acfc358343850c6f2c315216422630bf467688c07d893230eecc3c32174045b16f14cf4203273a47a068bc20;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcb84f45fd2dbd2087518b5d8bfe69364a6f0f0464c0f32f69301ed574077e366c856ada252b371048bc8a2fbafd4afbbca6d41e692b091afdac4f3d12a5f31b1aa4df51bac150b64d804c5a17628d2dc41d1afc835ec13a411118c9fbc3045c03843;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h332b50dee93886e5d9f3b6ba889220682439f621cf1a9f12e4e868b232456446c9e7bdc6807afd2b3c445ee9cca452834b9cbce1e9bac0bb76c6866c535ff703398640071c040778cb7aebbfa752591afcd11e0198f139d8ea0f05785387de2efdef;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ec6d8ddf86bd017c9642bed95ae64f74831e60a59f7d09377c03ead8024c50dc2720f8eb1c73e23e40a321c01aa94237d9a5801a4d3846c72c63a43b6027b9a41ca2c2bfe9ba7816f9ebdb57f1cd7cf0929bc81fa5d266f1bf27ec29cf690894ca5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h21e878357fbc724f7987957adaf05585342320b188b7720320c8b601f1008c9b373004069e9c9c2c3661197850124bfacad0a6858a0bf5a69a1344c5ec9b0c621ed276fade7d0e7ca6afff5920eaeb55302d2a3a45498ef10df6494853bacf5dd67c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9674a2d3713994959f5e7e0f1cd87a21a3fa5f025026af7b3fd684735d8a09fcad684140c0a5ed9e508c5937022a331899e6613050d50b5a0cfcc510ded8eda33507cccd52045c765130207d0b79fba0668728c1396cd1e1f440e77d4770b69050d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h668d3622716c99a7e7e8a57203f6b913aaf9e507d9ff44e02eb1cf1dcac09811c7b28b169d434fc2d6e54b065c8e03e54aaf27932e5ad81dc9c1b8709851e1895ba2460e5fdc213451b42dbcc8dc9dbd174e263e439303271bd93b120c4cb9ef7e7a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h112881ce05fdca43db9961352dc25794db2623ce7b1043276f5eb13fdee3583f2d65815ad4499b3b39ce8d325430213553d949378fb6748c904d8efc3a10545a02a96796b08574835979f7e6404e454d6068785d775632028a8ac34bc9b2d92f12b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h93fab4daec9cb360b2868e0ce26b99565bca67f458002253d6f89eec2ddd0f747435d46919564481d6dd21993417a1c9aa6b8a1c9d11058778eeba06449e680929320ef4259af3f50c092dd2ac2a28769e6f7bf069248207ff298321904fd417a26c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h114cd04fb8b64471fd6535cac61181c4e169d4b961f55ad83bd3f88a40d4a62fcec8d9592bab89c27cdf3eddea8ea971085c01a2335d8b94e1ecf5942a5c3af9046f0e9aaff31f11695f32dac0d682bdd640c31f6c6b2d8d3a4e9b72ac3e032800ba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h710b6e17401cee21c6bef6b3d129799eaac5bdf6821a0748dc94135ba6af59e127774f5f3834a7007e8ee1bd4c55112c01a6617ab0b972f01e8a843594c8f05974165cda916792ffcffad8239e46ddba130039beeffcf67ea38c2867d8d93386f695;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc86d3bb8a251b9d0c995d1c61a2c76bdd98987aa587b330a401c2dbd5e9750b27a6c00846b30fb3580ab7a0d948427f80586ac1a5a6a946d8153a4b283a34e34e2a867e291ee4e045a7fd210be9ab9332bbba9d544946822a81a04309f74c20524a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha56192b06448ef2750ec6b819e87dc4e6feac61a0d222db33dc325653b599cb42c5efeddce960d5ed1e3c1382db4e504d8861b15820f6b5447c8b9919e4d95420905440b1937c97b43a00966834cc18fd1e63e208c6509ba785c4b7d06830d1570fb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc5aa667afea2c38c215f11198de4430321e0b63f056d1526d5bd9f2694b524567de85bd61c245c49b6ebb4dafdb66d628061c9baed1c568f4d751ccc36dd20443e30cd886184cda06b6f6037b266998940332215623b27590151766a9ef537cbeec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f5e53655768fd26f8700e94cc9948f7770fc1ca9f9c9698772484350927c3a6ede701d43c4defeb60d72b52ed3ba377a9c9d0460e4b5b3aee35964d64626782f0eba31b63e7f6f4e6dcf47392a524d2338783830b60ec9b5e1d99be8f8562a6b454;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6ebb1cffdab90048f1f675e9e8940a7158097a3752495a12a8026ee31e020a14dfaeb6734f43e6bfdc4656e81b30293ec7d4f68c20e782c8fdbfced46315c11445bfa7d4e17b3a3484e138a07fbfbdf377a3e8c2d71e2dcafbdc9d8f898036c14aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdaa45086fbd10aceac13de10d483d15002822db7de5615e29d700393d58f969c22839375afc10369a936ca1353582a677d1f4da1651b8fee723dd7947d8e3f21139a6a921d2d416b09709560d9509265562d097ac7fe9d5f4bea890e326d209cef01;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h973fcaa81bdda752b22f8dd48497d833cbe44e298fa7b4bec9421b80b2e0a51d46a73791f12c71c43ae20aceacad44bc07e8383abb2101b58a8fa3eb49341ddc884b19b5674172af68fb37fbc7f5711017e6573e044d49db608cb548bf0655826e67;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h347243a776ae30e15ae24e7546fd1142f3c57f348a582557d488e626d9e4696936a5c006b1e914b70dce69a1257830cebf87e842f942df4f069f569c583ec4b9d33f0327ae0199e5eb8d92339e8d13006d099719e01fa2abd3f938380690c076e2ce;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b86e90db235e9bda37557788dd782cf885dff6a437569da32044390e29660b5a5511ad40ffaa4bc52521a04cb91b9349b5ebf400607bcc598662a391a0fbf31de1272b94830a36421b245bd9ac66856582f15c3380a1400ff80dc878d4dbc684fb6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha6953b7182878c4c8030dedf3e2bf618fd18faa5dbed07f160db63f409e76a88fc2332c52f15a12e0e7c4a8fc9af07f9e1c2edc5083e445ca8570f816523adb6b79fc232fc39410bff79bed633c4b53e13e0f6f4b4cc2bf801210e69c1347bbb8951;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha3e814ab2a886206f64de9fb4bd5b98a2bf2f2c4a89505fc39efc86641eb496e6b856b87fa7d82a2d16d78180b5a6c17299bf83e397b62709530958cb10ae7c842373f7cd71acd1a8613de15fb5ca16150f4e6a0a686341163f4f59c81ce8519005d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd671b2511f49e7f204cf9122c29ad64ba9c2a8dd115df06eb20c588e23b3a7440e7085281b450184a3a9270a955f8dc708f4e39013c3700c36d8e6edd007745f1a9df626c29f6657e30a7cef031b3df9b7083d3474c8ca94342b502d5cf4bcfaac68;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3c54938fa66f729ad4b174045ba5b2a58eacfc5e3c8bd3535a94c43e0650e6b47c4001d206b6a9556f1fc05dbe7501cd977c2b396b0cf8e998b43c709dc34c6dd8830a60c221368e2e0671253d6054baa794eeab938177c6ec458184c7b0da85a7e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b196ae0e29e91a00ded4dd99c2f15cde52848cad06ba567c1b15261eebf719108bcbdf6e77c4a8f9fa63d20d9c4d918f570d63684fbb4105d68299f1ce1ace0612d490d00cee42577986a773575ddeb93ea32b0fff5c9627a7bf0bd3f59063c0af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4f295c0c83006af75560eb6a42ba99c6136ad53dda2b5bfc05abfc759d1b16e7067993447748d6c0bfe7f274ff1525307a9a55f61d6491f22a8eb97d8199fc234ce6fcbfbd7102bb55a9c2ac4cb233b40dac6ebc9c022b64e7dcddf792939f3fe2f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h29aed5222e5ebfc9db85c2747d18bff192fba5936a2803d1d21a8e9f92f66ec406953006738d29990dd33c998af566bc673f2bdd14f11c38201057f2b2bb6f064873c7d6fc9d1b6deead0bf222cf68b7e51a00f60843406e3df2e6bc43aad9b7e899;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d63e88f96b453df103560d14eefe476fe9dafc1147766852bf55c8567321594021f3e63f607a1d21a9e8ea1f972337473cc71ffa5e954067e1e1cc2d84288171778717afd124361d4e68fa43d1bde26bf9c6a00c20816e7d2d316e0013f96295538;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2e0a9b6758cfa62a628cf1612617eafa41635e23af96e2b414edbc023727b524a9657dbc79c2df8f80dde8558a43df32baa761b83185cd64a2959d109ffa4cb9b1f02d9db01131395511a8d257e55255f57ba5dc45a062c91f5d9807a32fa149fb98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h117eed998c34a399e01b864c01913c4135b53a0fce2d395e1bbaa007320522e01ad66f2011b26431519c64bcda286d1fdb3dbe833cb7a8758ff52852ffd3ecae9177cb3269c5967f73d89674e6a4841099f1ad625b45d0cb00395e56e67ed4ca8532;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc08e9fa2bd9ebe9b801ac696a00c8d753860da47edd0b8fa98dbcda21d7bffc981620742112e797a493b0edca54073b740e964207cccadebfca1c471af5f210657362c963d7f243767d67ac3da4b1d3cd448bc7cda55af79a74a9a2ab6f2bced1c3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbde7ed84472ed2e20f0b37705e649c8cfb88207eab263068e1592be3dae22968270426ff78595ba1eed76982d7bfc995a4e88821833693e6d7d2ce9842907fb33ea0b759f2aa5c802bbf9affd9cd58c8e6391586382745943bd354aa749117effa48;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6d04324ee31522e0f63767093c7ecf0a525cf582fccadb1f9f911fd34b96291daa49c40b1c291372e8fb6b1ff9a9e571f98a0f4f98dca5bb8dea6cdb825e4ace681f81ccacb58e23befc44dbff036dbab6bbdba85d7fe17eb337c2ecc2354dec29a4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89a96ffef2566439d8d1d2cde8cd8475c28215fdd9ecbc1a59838980f5054d82c681b5cb1151a702546275b74f77c1934b4688bccd5b4376f9ee87e3771ff753f1c4b67390949d5f680045fa9d029988bb402030aabde7be491958269ca2c461a015;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc43cd4f969c1554f999fb3cefcaabdb17dea878bb69b863bebf1f14ad13f74f572eb115bcf88f02d5d792caef46a6d79fe3df4d88c05a2cf8f68968769475c3f183698d99f0c498e6afc4c6d50065ae933344786a92c2a838bb72e1b53acf9dd4328;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeda77fbffe6888fd77fbc3e46fc92caf95f9a60d1602470e12bcee6fd9fa290d44660385ff3d96094c47a848480fdb7fce6ab86c19cc00975afa5cea4744a85dc9bf89bcd80b670243ccf7eb64e6c9c85f88496240ed402ed1c45e0d472d1cc0ea7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39040bc2d29ddf00f9dd29712b4fa5bd68b96ff15006bd7d7391e58a2128919874afebdb5dd2d554bef5865069ed5e710a975ac28454080f69c52fe58c06f56ea9d0830bc579b7daa66ab6420a76dc2ae1de608762981ca31889f1a7462c8b0e6948;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hef84b8142d5f9843abe51a50e19edcf539559fc68c9901ddf1914067fbc9b7025a3d43fb95c97851fddc854633cb6f26a25f01d43d019472bb6e41d138b2fc4523d20f02f4c22f01374320e4bafe4fcf14336a69c9b4377943423d7028bc89ec9c15;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96c9749913224dc700f2726507f4b9e4b21a12eb43653b797ea1036c1680469ad2fd9855d55708e84e38657e24220a707304f544d9de96f28a160065318c3fe521ec42b80e708324a29f82f4b433fca0354c91127262c7651fa4db285e6f6c4ef978;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5257ce2b8ef7942a9ccd764217ab5db21ae8604392ff6ee11e647a0325f8e88c8ba6f6cabb52ae1889774378ff2b842e484a308fd6ec61470c205d7420e46edf3527136565a7f41988988bdfa48e654271fc373e693c3369e3de1d60f7172a63ad85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he0a6f7a16c897beb609438482770c1b6fff9bcef09f4d9a9daff8a2c16c0da13794b87ce5e6e01c3029a3b9095bd75f8e3a23eb2602b290fb8d2da84740b2004385c1458251af3025cbae3aa0f72c5578bec4789b4a2e53140d6b55cf23e3a4e3002;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1f4715ea53c58b05d002838a834c326bd11c6c3b80f59a136a09858503b09de30a2fb7e594676bf75036a0146a9b5739be2564f428b864c9dd81323364211490776a465b78210017653dfcd2d9d681ca6491e31feb17f3525f3a399d1f4d5fef5d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf25e560a7fc1a9797677ce8573a1659f7a1075800bae7c81159a9310352e37c73bbbed0059ea1dfe5a474a8ab91cd4e0b75b9df4d6024794f4aa03b9bb8dcdf788ef341020d97535e2c7d2cd030c3dc974699c2dc227136077e0f0db265cde8b07a7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5a2cd75bb2d90b65eaf94c3f0f8e3da64ab4ce8eba06366c8208c673a01be94d2e2782d915c0d7b90a801a34d45f11b000ad21b1b9fdb334dbf14632eeae55df63b3976baeac2f188c807114bca7108bb8bd9c29bbb2b07d0a5c170fdaab13588393;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb3fdb93925b2b489f8a71fb04d5996827befae7e77253d29bd99d8e88cbf05483d9cea3ad8162b946ddc5890bf693e893973d65daf2abdbcf9a0eca6dcbc22da5cee530a9a186c476640ee1b6011e9144688f4c4cb30a8333c43626d7bf4b95af2a2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdee110c0b21faa9cfc74421e95fd62436a7156c9826cd02125564725190b661f4a06df05d80375bc5971d0b1a4f22fafd933bffbb0e7c1df6c982fce82e541fdc3c98d71557a8ab13662c52acd215bb82df4d5f51eff1faf5cfc6c302be134f774ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h99498824bc1699fb8333e925f60826e5f73da4f3cdc6f6ffba5ecf6e02d11d77fb5565c4a328da6bf0015fd7cea8b638cbf14c17c2404cee56cc7fadbae57e5653c377c8e25ff9ad3ecbeb746e1f8c6a9440f6504e57d5bf5054997ca1cb8d547561;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd72ad7f281f3190669c98302f9b98870f48422f4c42f0389ff4967bcab29c33c14634baf0c206bd51c0815515b3f09c6b0c2af9c0e6a99e477421e7c5193998208ef5171678595cf43b4db5de6d1a4e5b140fc1fd753105235525299bd31076ec6d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h241a10a3fa4dba13f31863b814560a6b24924952e27af68d71ad78355ce0963c12249c68377478b3e36f9e00e20e00746768ae786530d0d805a1013136782aef718512c3c51b220c5680cb452cd050ccf6fbcfc5642a363fad2d85a6d00af103488b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbe0dd4028b79be9f7ac1c7f1df8494a89680288ef6a85f6ef5de12f9a908ba2f4c24b6118d28c199209296b9ea5d9e235b53a4a31a16ca94dbab386e8fb91b772062922ed36fc389c91de198deb4a34881963bb1572ab94e89740ede950721f3aee2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdec654fa25a1d237d742843d761a48a949d6de3318775f422deeb7843ce72c9a44769f3542408f56a65d829318a6201c3855cb096934e296d31750bf5e8d8433764e8998de992bcb3d547fe04fd77262065cd7dd58e73b0609d9d5821ca5803d4561;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfa9871fa8b646a74b24cdc68a3b7e13c4dd90b9ec55b51261db52baa26424b4abb7870b4645d28ee627652b8b7043da13340dda203cc6ac11818c62b01536780a72d6671ba69c39af03532ef0c6fee3ad19a02dda2aff16f66efbcb3d2a8d9c52da;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d19f54e29f9353acf6bcadff60febed655dc0427f5ae685c5e5c48b40ba1be84c3869130761ff85c780977db74cf08be1fe91b7fed3d9e1340cf8d79077b5214be54e45df2bf034d7898ce76bd78d0e4530d85f764fefb99b89debdb4768d106782;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba0c14b547fbfa7f1982159515599cda2409d6c8faa48a17ff960a49162c3aff511b135e6f2ce858238f3f375c824c742a548ed232f13e61ef074f454dd40331d53bcdf4da75f3503951a2d72e698f88bf1111d4bb193bad23d608e961415b756258;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5fd910e75a0c530648c9b7899ec014571771f6f053839b98083e3bfdeb8a0ea55f0eaa84b501cb15a454450fd33ae44bc3e28e7be237eb5e781e40b318d5e0ac73661e19830dd96bfc019f1e2d58334e339db3195110a9dd3260631b5bf64c7c48c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfb287fdf1e1b3263cb207c6b4d38ce4875356ee6bb37d99f8781d76592d08c243b9a7e3fcf107939035c6aec19ecf45ba6bb7acdf8d2ef8839158e0ea61d137fd5afbf65c64d7a2cf6eda720caa5fc4ebde4343b58e47a041af42c62651440effd8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf9f5412b25118b321bff2ffbace75d08b989ce0116459f7f8610c597ec57a4aefe6fd21b71bf2326ccb5712363771319aab31ea36d8bbb6ba60e4462e8e7bbf3e0a0d8aa69a9c90be0a744e2c11ddd48ab8b54ebf5be8bd0a74e1ef7d0533e5c0f74;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h79188eb1c55f4e8da20f0b320ba8b3917a396da3258a5ad50f5c8499ee03beda44e1c914d93c7902741ce130edf771d2728a1f938fef620e838eb4341f9b8fc6ae36ec42abd677207124d5faf74e3ee12d44c5c6280365132ca50f3cbb65c5389fb0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcccdc6a0bca9951d95665a5a4540f38234605099529b7f83ff126caebabc5482bf63b97e091d4c217de86fef24e61eeb948c1974b8b240d6a12c13e3642c2ab39539e030821718ba5a3daaa5db079d9d4ea011d52ddb3ed0ae3b2fe12664425c5fbe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8eaf1972c0e06fe38cdafbe509d1f1f1730d2a1bfbdff2185dbcf27785f49ac32c07d87f86beba5bdcced2f3b79516b123ac01ea9da463e619924b3e4311779005504a1a5f4e475d11e157ee9d0ac32aa32aca698f8f00ae3c4e08f0a7b0489b652e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3712bd111d9f2d4ee7c84f2740a4c3f4382038f9b7980efb3549088f7cc519dc34fec9a154f68c9a1d0a9e7de4183f0b077c55830bb4bb6f26802df5c3a1a25060f415fb07b389a7615870e474c5295003a4511d6f185f0efb48288bb102ead0012b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8bce3732e039716a26391fbcb4610df365827b30baeb738eb6c53e80f6663194538a9a4a0ec4a06a96fcd7cca3a41abee4d3a9988b2de48debf2d54698850cc3524481f0802e169fd7e713305af0c2811156a562fec011995e96bd1f123d38d68b56;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd66f575596a2199945c0f8ced78eca549d9f8e433b7d824a9d828b2cb9c0358612cc942fe34c73384b25806c5ace7f8848cb99993e995958c8c0d63018333e495912c6ae9364026eba0f1b38d256b08e69a981fb2f194f1bca6c3e045d2910f4c22;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h91a6f7f9649d042163d7725520b64bacb8b07f1e419884fad7a726c614e8cbf60bf727d5c69659207a1556d2b3ccde50fd470038308e95c82f237fdafe1aa1d818acd578ad0792f65d70010878b7807fa2797165258c927be91e0e7fd284eb71ce8e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h868c573690dacae7bcb87dc4f5ffca214539e0c2b54c62609f13a2e5b749f7278ca9d3e08745689a9641432639f70e68eb07ab125a127e8556ff2b50b89db4b1f5eba37e49a81dee5173ae0bf705a69f468081937b3e163425143a96a1f7efb3068e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9048a01fccd171341b0e5ba46b13e7ec8beb8d0313f55bf8c719a06826bd4cbcbaf247de27189574f8d4f298867e06882eaf2a9ac6e84dfd64ea356429ae1056d891d6d8b79f414a59b0eb022b4f129b7b7751a59d7d48e3b86868c3980048a1be11;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h25307c6e491968cba791d0a5d4eccbc2e7590606b7d6154eb720b0e3523f33aa8944a258b5369b2f43b4ae7400f9639ad91c2becc52a835f4ebbf12b023682ad2443405c8d8f93682996a51c45c6d0648a4f1db7a836e48ef50e966d1b3d7461dc88;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd009285b2946a1066e1f85e3d3c81fca9fa5eb1070e316ba17e4452a27ef33d191af0d676ab47b0865ff19ff35a33b8acdb01337db82dc711f85880be57487041299cb3ea13b8bf86ca63a81b1f3f9c7f8b6570ab794f81c6799c203cbfff8db21b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb56e80b7463a0e32555064b7668444e3fbb2ebe1f8144f7ee74638c47dd28ef8899190f9c3494527f181d9cc9980da5cff2592c0ca9fcbb3db5ee175da5f96997ec3fab644c29a4fe5875adfada5c3f84517768c6ae1734e2f39c50d04fcd5b2be3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcebe7e8e482ff1f18fe6a7ce4b3681a0c37cb6683a9123d207baf4c3297cacda73e53449aafe0a557f2abebe5685ae0c97babc9cbb73a2282ffbac45aea3cd5a4998d7f300f9cdb74b69b96b0ce3ab8f050c2c401c13f5feac6394f62f5bf1d8a7a5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb208fd409179a8de193ce4d80ac273e89d2ea967a079ffaec1d74429ea13237ff76fd2910e9674b82dd4616a3646e46028f3436321dae758663eb5233bc5dc58ad5dc72dd012daa8bb867c79d11f30c4328c1bd8975f44b3429effed536639ff2911;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c4366550f48dd9b087180f02b2ca4dc1dc79be7d49b167112c62edea04474b239f2c10b1fd0b8d4d1c2d7f7be5ebf07291e26210e44aacb1dea3ec63d748464d1a089333ec634f49efa6d084e0b59bd7dcb6949ae6fed6091232e7f322f324fc3ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h89cf7f74a60d2e534d3edf952929d3f351a9e70f5f884a5c1eaf4165907c729bbaafd60a030c3d97188916ceac49e33c21c91fa82044747f7756c2ed079a7942ba03a4cebb33cd7cf01be700deca91f702567d2bf0011bacf3a5fda5527922b0a3d7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee2a183d0cfbc9376bb1cd33156ca4abaaf939acbe79b4e2746dfafd36bc622bf8bfe05e5b79803e3d4d0d3dfa888f5b7c4ee77bc6d097f0038d542bed824609d31b8f4a8a2a5d506da191ecdaf101adb561fa45840a9a797fbef0f6393a171a564;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47fd82f829f97fe949e9b78277907971b74ddce16edb03868cf2c531f29e52023291ef8a84a08523654840040fba5cbd2dd1b0dee3c3fe31053a6f169e45628f94e700486f8534c8bf36b8c7a3a1994099bcb921812b68c1e63c42140fa45041a557;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h995bdca9888b0a54a6c8ee1aefa30bb5a174584fda60d244a8efa6cbefe368ce98739da75dec48829d0eee697c4e0b28b2bf9846a3f7805b4a084a9b5177a43e7b9a05a2a9e98f4f69ef737e1f3f8102aca5de8f2695bcfa42fb255946a785442ad8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd200c34b3957aee015ed8ebeb2a6323c09f6a0c34fbcebdb4d32e7d271029dc54571a6623704cb47b5f8cc7c526a99c9e7eb000a500bc011d297c299480069be84801a72fa27988f014398970f853385ad1a7e174bec3fd5e54a5c8310fe40bf6eb0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5f495cfd905f7f2157731b760a4c0789e600a7ce6f0ea3ae82ca8c7da217b7675bf4abfcac3f3429a8abbec329d7c3b2b40eca5d7eb91b8e9a640418e8a049ae7c845fabb400cbd679a2c142158dff9f6cbc0f67cd3e9dedd0713e3951dbbca21079;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e82e6b4e08bd1ffce9d42520b5c6346166a1753f6855414f83c1c3e39b5f97dcf48e0256be5683352930631933f023f1ee8edb19282515844a7ed5c61494505170c90a9df8b69574ae28f89c95ef1a23b0b3b33313cef12805d062c7db201faa4cd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7db79b066fc9af40cf67b6c8756982eb08065adeb6fdf6aa7a568fca865f2255e6d05466a507028c665837c9883ec0ae09f32f441424d6f1c851a2f3aa2299ad704e36ab89cc8ad0b1b533340e8bd609a4287d30f41eb308907f9feca1f2a1a3834e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h57848f578025ba99c872fa2c25574b499de7bb74dd929af40d7ffeae0757cf856eb97df961d830fcc1279c8a801e8899f89349ca98bec498520c041e245385010b01362c025f202424ed2693300bb2bcd9f8c9a4440002de880680f5261a23b95d0b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h186d56e5ec8b79c885e840675c1879cd1c8a7bdca9c9f1c7efb154708a77f3563d7c0c65312cdaa0ccd91820a9243d6453e48ed00d5f72130ac5c0f1c1cc2c1338722f39033cbbd5c4c40a2e611df77c086cf35090e568cc2a2e166078f2c249833b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf1831ba6b08449dc5c329bf2993ac0d41caa980b47ecf96c62d8f9dd225065ee9047667af80207a46728f8b4e6ac2c6d93afe23e16dec6c688af7a57f3dc9f435684180e3625185eb323ab98064e8b0051e975165b05e2b979b7ecd844a416b6c08b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h10f7b534f4808c347e13ec27b95573f474e41b21c45d85978aad7c0b7a4df98235001660a94d012e8367388ee6eb6c922ad239879a2372d25c3b635274f5a544f48cad90a0ab129aa1220b6142f945d59f231a95b2f8bf336523852dc9525e213e64;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfea1792921d86dc00dcb7ed473940069c79ceeffc27828771117b5b37d17977537ef3c372ae89398d350a9c973671dea7b8d165af07e7e162e0ca24de6c386eef481671a486a98d64d44890dc1e0da7b0e16d7eef65a010838de8d9f238e4254243d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4bae82dbedd994f9851989568960b0736513bdf62179b1465b6b2246ed61644152cd3557e386c0ef84c1d6854382b10cf3c378c6afa94979e2519454b941510b79908d35455cf18ad6249e43520a4b07f341ab86999beec437d5980496fdaaee5947;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf70f44bda16f07ffe246a579700c76434f176cf7473b9a6c4e29ffe88c4ce80b504dc4b00fdcdf37abe95553db48152f97d5e82c0d5124c6a60cd3c2366cd7359b94efa388413e7d52640e26d14c753e4f21837c34f170fc5bc4dc1166bbe07cabdc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h727b541482c510e154fa78066b9e48b47a7844a50295136fb77852b64b017b5ecf555bb240eaa3ee856c418b7c3b304575c55f1d1af286a54eb974b6a2d14a297cc411f893da558e647becf1d6bd401a5ed50587323e62611561350eedd2460b494;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h44b964affd36790e127783d3a09fff2c2a288db26ed280110d22404329847b9640c89b8e4f9d5a524aa056f7b22208cff16e17350fd5e9e00e4802ee3c058e3cc817c7b39d7e577833a38f90e66faf0fb42278232466f8a683cbe7254eb43f77749d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9ba18c230de12bb41df2694079bfb2f1d773d4978aadc6923a107566578a191a2bc072c037c8dd09ca9fd8e9eb1df2356887a24c39ff9a9d21c9e98f8749f07bac9b156dabbcf1dedb18b680807ab9af421c8f642d7c754e18d94bd3165513b11b3d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h983b2409fcedc139ce2d5d8d77f34dd4a1ebafc8b717a9bc5b22d0332a5a12e5aa7237652593ad51dbd6f186b036c43ff97292ef433bdaae827e1e64d4251dd6a82fb4ef4b00b4317c896d3448c24d45bd7a8ea4b16b0c5e18a3717a214108a42479;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haa73c2503d2c1b92f5d77b71d08a45faa005fac5041fcc4b2925d683a1914bc0ed2efc5096f33da724a53f9d6abf6c09f33760fdd1f47f1b49436508850d4e671265fa5621bbed0e4cf5750bab4c9cd6f97f3bc84c16ac9a3c4626ef344d18acd827;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e2c5726d140b4ceaa1651ef3892dc7a615f9a508f8c8a1cf3556d2d834cbe90f74175f26b10165339acf04ae56a45e7ec385bfdb85d8d9ae708ea09b9964b3edf69789853f9d6d4f416b52c4953b21cb8744ebe05bc5ece0f10be72160f9396b0ac;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hacc3a0ee3667331d78d5f0926e3f6a3044e2ccae2cb6c1c957322432b537b32388ad79bcec6d4df810948ed53677bc78b2c6c1686afb10b057c675756f522f52ff65b9b7dceb05a5c2b43bf122b29d5c29760d8afb4647d46dd8e9b465ce44d1b88d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbde13c09a413f752b433a28b7d541bd8d458acc7b8244acf8ac2452ed57e275bdd09c79b7fa0e3b9475e9d7ed9d3d799f91b1ecb384821dc9f1a0a328b7301814d91da1619c2d9a0549bbf59027c1d9aa790ef4001b71abf1a6e688764710ec54487;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf97a20edfafa545e7d2dcdf536ba1b0edba2ea2fd3f265f8e016da9aba7faa873fe0ee11dadb4381904203ffd03d3efd55c7cb981f1f2f50b8924c0c5593c463ac4d7c194a63dc9ad5ea5a49ba496728f71de7420099ada478be3a5dc039496abf32;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd45b78366dd47d66854271c691af258903a178c0dc2bbfd8a248125486b860010d05c3cd347daa2cf5eb328afaa7921d7044734a9aa1533048fadac99083f94726d6752abfa8f1443b8636cc05b42c56541c5234653bfde99bc7e101565735783a96;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h884466523a34818027af49309fdd5c31ce10023e6f9460c5f4606b2baf1391632115efbf2c2d6d51faffea4de69639f97bdba1df0d7126d93c590bd73eb3738a725b1315e1668975c4f438065d76e38fed506b1119661eb35d3da4f763cea0710b23;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd4238f5108027144d40d14675a607ce6e67519b584ff6fb205e7e7f8df9a502b09cc719fe906c3b6eb6d7cad87aeda4f79171ccdb03f11541d12bb39d9280db155bb19083659da188351ea2d0d5938ddacb7dc2aeb3eb1b7c2466d99427a9a54e2f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf2b514802b7f44de9f50f4ce7078eda9622afcd5cd1c55e1771fa1061a5ae09e56db55f7921da19fb8e2cd29a274ba682113809608ef458ea1c4512e13640068b5866e9c6dc8040dd652731657715aee5f7c462d7aadbc9f646afe6c470cd9dcea0;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h681ccbf8bc9feabe2feb7bd6c7dedcca569087a5084fe53efd9e4deb5b3e6f59c63279d1ee001b863ab212b6d8fe057770cdc2afffccf9057c700ee91031307db72be95c4cd750f976a188495a748f168eeede4a978fb8512cab654ecea9098f030d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a243090be4c4084c732367c88571c20583d531886d22e400fec82095ebebdbb580e5838e606e457c234904841d94027ee491d061dc0a3913a9a4cdcd29c247c7257d358db7fcefe856bd3c22afe1ca54907cbc78a3b7d7306cbe872fc90335dfc7c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha670e3248ae1dfbbdf5af1e4262bf07308056ebd932f264a8d68a49e3c86244f7ef55b916f0b7a2ab1e22cbbf91607ce612f0c843d3d369d9bc7c08f583110aee00e638ab236edb6583bdd2a1be8b68284b3e98be6246384f390b59f1e6497a7c9cd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'had5cf3c37da2076653309dc51cd3aa67e2fe285d21467bfba70969eb770a238f60d2e4c6c26649c83f1c6a86dfb0707400037ced6b08202761f4603ebe3d5ffa01ed7fcc14cad2b81e90a6ca87b6e8c5ff0245f0dedc64c43679eb83bfda84bec7af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca6cacd07376458247a376fc677d48848550c523d2c57842394e988cf4948354f7875c815034f2d662d8491c3c8d880ebd7c54826b9dc8fd78c713e60bf15f2a0f8cf5e32136cd0b0392d86069c2de94dfdac49bd550a761177d08d79b171fad655;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd76381a135216270714f81bce16c59e1fc9af54dbdddb065ac1af3ecb4bf48a0f2362a590a1aceb75015cf1fac276369def9c47d606dab2164d4863d72955c2d813c2ebaa3e5df95603616b06f61bd6e23a2ef0fb3c331faad5c90b28a6ee2c36f6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcbece6688bc97a5cdc358975b4a3d040cd8a46954c75bbed57538a6b73d685d4f70f9b03aef365ac467ad7bc3732cd8e1c265105eb8d63e56a5bfa16f24d96e29d1b4053a632b8a550c660e194165a71a4161dbeec2e5ef0b8a85302059d172d6efb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3783444398ba41f6c04ccb5defca7e7d2cceb244719c3d6379b9deb382b16e1b9256993b3d097f3d406f525fe79d8304f5e2202ca5c500e41b56d90fd74a25564360511db9cb3eb8aeec530c5d84b34dec2622726dcd92ff8ea637a54aaab90b2d61;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hccd9aa8b02fc48837fa89b1bb402a860c272cd09a3fb6f63ebd3cb2e1f0ca6fd5a2597c665c90a4866e7b76d9d97f38b77b8e7c8f1d7d467c3596e23846f2cf4682037c5ad17e7b40d0ec39708f5be9e11dab6cda438932dd694906ab2582f652a85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h647536ec65b429dbce3711c343982a2d6ed9848903c8688d3b918911797803f6623a02886ce269a03479f1f805bd2fe0860b3aac6850c9a0b137dee730376642a4e33eae8df5600db0d1ca9b1ef06a4b272509d4ced5e1e1544a2bc15de647b32cff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb29b3124b03a582c206de30809861d7b96075a61881d5f3a753191a2a58cd6791d89fdb4dacf2f1da5acc18ef694062164fdeba7c3822db122534039cfa32e0983f99ea3494cb03119b42e2ddab515f1e4a8dc18329f9de496878296ad00699cfd5e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55d86dbf4f505e63a2c41f39be410afb18af17579916e42056b478191ad9f3a116cafd750fabfc3ace145f3a84f295a2c21fb958348fc35b78f88fbed2e8ec6695bbb9bc3f1718cae33297c59649971100c09133bb9c9d882340595829f9a070e266;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1d89cf3be21ce45fb69a4be4f97903329db06bbdbaed8223c4881985449e32c8679cc89ba10902aa6d0590ad6512e92a2aa514f8e428cfde9a02db2c7b04076506903796520077458a883e27adc743d2d0353dbd774497b828506f14b39b645c0bd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h52d10aeb140bad1182427670dbc48799f23ccf9a3c1dba292ef72c459f818789108fd6f17d9f4bb93ae73f0eedec548085679031bbfa444d6e03ebf758bbae6e7882c2f51f2dd84a4485d9ee460a2d6d2978fc08001ae010ad6af9865af3bb3c15a9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd6b216a7e2c4167767623ab8c8ae0316ea807d49f0512d26aee31d7ed719e3eee6bbc34453feabf35b260ddfafafc0a4cc493843ed727f5377ab044493b478dffa05cb8f0613f59718111106e8c831ea2fb653849012785325604b6f9c36116d15;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf0ae232da29c7cb5eca63898c97a596ccfa013336c1ba64f58861bf2727d72439d1c25dcf1af4aa6c78b1ab678443f4f017d7850358351c4fd590f306aea79914808dd93ad4c8e9f808b1c738da9e049f5a028530701a81e1e2daebe83cadd95ccba;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1541797a90df78cebd1a3cdfac2b7f7d51c7b98604c92f0e5899883f31b224b4fd8ee17992ca600901e470097a709541281f96fa852ece0ba4ee243c4b9644c2e97bab5a357fd88edb3c04467555f44fade915341aab4a69d7c51ee891c29305019a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf6c38fbd1483b83a825fbed0da1a2eccbe199f126808b39ebcda2b17d8ecf2392b89fdb9132861984f83f86d406f67a7e5c7910d9df931e0ea41ebb95643b16a6698f1d4cb370fc1c509b45e986ffe03c5f2bd01752c09ff2cc00e5d08e7fc6bfed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6dbedf9547db1743ab677f5ee070f26605c766e037a5b79d5a6e2946327b1d6a848fcb146778c499ef89f13ed4684fff3271f6e33c630f50cda8ec1471abe58d4f39b1d405847747baf330cc8dab784094236afc2c2e72ee84c62389b459632fff3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69e5b5ebcef5e91fcf6f6130d739e06cea061f0c48a783c3b7343f5a3b49be142e9c370eda3b3a156b287cf873a1fb8372b8b66903fdd4d87c16ddd73758ed70a8edd66ca7ad1725d0da2bba615984405497279b3b96a3f6c080b8e107b2812a5f92;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5762e0fd125a815c7539d25a385f2257a64b11f505c634e056f8b4fe2d39fa9515dd0998a28971b007aa8dd427d30de85dc5eae7616f3e0e75f8b9e6699d4cc95ce6881aa4f78a7a842d1c9e276f8c2b36bc6f98b0a5de86571eafe38c0bb8a0783c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he8d9ae325d9c8f48a620426cc4bff4457f8c13b1cd40164c42503e508c82e73fd7132e9a7316e6bf8bb4c48a27f96ff33afd534c8f6f0a4f0d867de7bbe9a9393e42d0e8f44eb5049dd3e6858855f79a4defa0fb1048a9397092a5b599ee69b59884;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfe7f573296248b3cd9e8bccce7691e93a9177c55c2c85abeba44a8c089bab712ebd72bde0c73bcfdc9e9594674750efec6e8f8271df7e52d0c3a9ed26c695bf4e5919782e033890ac915bc5f6e223d5bd41413dfc0267c6f5520dbe93da5aa7fb4d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3f8337a3b1ef7e13deeb47890c1063c8d5d1f61a415756686882b66724c02022377b1991fd54f38e38634fae98775139616313e7004aeddb73f580e6ab23f65345102f13ac794636ce925349721e7fb410595d1f8b1126a3a5f2c5e4582785b5e52a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3462acf2a87ca1a63a91852c5bf72ca6216fadbd3360c567d0589bf0b34cb12e95dccc2fcb75c666fca66a955ff340c665d25ee862539d62446a877d6d83ae611f301976fff32d55d2a97057f3858e2a4469f89d4c06203619b2ed51b8f8a602f8ab;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha338e999ff602c92460af1e200145bc336a74f86ed951c6d3852b90d61a89fb819b8ade37ef3c460e26fb717b31a82985026347d1133ea60f0ac4ff22062283dcdafedc179fa6a768e84cfae08d029e3b889191818487bf3831683ee7d1a5be2c688;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h518d35854fae10ebd8228ff91c253301345f4c31c43f1209ab00d2ef58f0a29d8a617b4fd7ef5b928d041e1d25ce58982334416380bf3978443a7a75be67d3c5455a838ee1082291d4f11201abf257eba414ccea7c8265332ac9cb95b50bf938292;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h5fe410d22e77369567c2183fac3b8c27002aaadda763feb3765f49ea577a3490445a0f9da4a003fbf9a555948aee7d0bf34f8ef28e9aabb44f2486aaff096408ed0f984de52f4c3a09bbb79b6034c419194ef00bf88c41045c30af8f2b79edee7ad2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h759bdbef78cd407b5c72bb54bede239503b429e8ec2fcb4cf37750c7eec23b726b79601224dc9d3da01688686102a6eb7988cb5a68845f33bf0b684d0dac74e003bce5552f929212634f230a87455c7edaecab1d9596806d797ef8ccfaec7abcb4ec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h19d040a3afe98e916a631132b193bc8fa524aa67b8c26b2d765208fc9e98e56a482b4c6fcbfddf88409cc637a5439f4e93850e704b24b664604ffa9ff6a470cdf6130914e30afa096e22d3b0608045328d6c1a57b9b76aade1f8867f80f4d2492289;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd16b526fcd45c4fa0c7a0d37ce04cb4c2681e344a12ad7eeaf6062724708ba0e027e900dede64bc45e4c222986bf5b7b822add592ae02f3f2d4526f593eceae90d45b6559a4c9dc85c0550ca69955bc758186d8a0df7f02f89d154c555f6c1ab8a43;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54cc5a1d4a8807658c711d80361645be11f69507118bd2d5afc80b77670d4f94fa29cfd060d5d66dff361bd4370839291b5e0c1d35ad28a2d32f43c51906a27a6e92459b8e2bb76a3780bac1889d2db20f07d53933181971b2f03041d8257ccf276b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7e0f76ed6ebb7d6149e6b4891adff252ba5b48893555ba75e670d698eb0af78743c8c1a95695467bd13ccef5f641828e9dbe6c39c55134e26b318bebd163fec64e683666fcbd5e12138e370ac3a3eb0452689d5f470175b5e5660571bb7b6eae47c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2642f48422d83e4fad7ca265f1c4a6b4d6700c5f4fbf69fa0e9c4fc9a2fc57f434cc5bb284b690f3b660d5b17f669c0fa74011ec0c697b81f0a4137be78e5d3d6707526d6d5409e3448df3cb2bd0392cfeae0204b4eda2664fd72e4889f48e6991b7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6b56d8d00b4b2dcae16054b306d1c24deacf4404b01034d87972ad12dcc7a322589093b0eaf2376b2d9348cd37623414d6730e809cca24555edf1fd2eb852a42cdde3f9f2bc3f82f1638f20873306fa91299b8582fa30cbf30c4bcf04dfcfcf15f58;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbcaf29cd9d3f18900ea24c33269588da58113cdd2718e600228693e6c1607b1545ac6583504253251e29c8d22b074e71344bef7afa815a78ef928263ee80dea8cbd954fad7b34da62a96f315cd8524ac989132d5b42ffedd944f5115fb87faf1a5a7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h229791493c079f821fbb7bd35e01c2e3cdc2d1890c52065f9c40b32da680679de8675412b56f7698fd69d2611d848e2e435e1e8a96b724ce9397fdb283ddc88b0bfbfd66df92e8ed57337dc99672b58b0bb8f9c37ec7ba4d4a20f74caaf7828ce4d3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h753f21b1f75ab95a6658967d856866f51fff36312c3c0b446064d50f4b60c7e01991e830ef2d71bfad7368f7bfefcabfeefd0b2ddcc00cc7da91e332c14de8fb8918c4466bbdc87376bd4365c33aecce4696c320755c1ca47c42a33b09dc5b4ab44e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4f88d7fc2c9aa8c437ede05951db4a77a0e2680d2f1de7ba0ef8744b447e974d53bd4fb4d09c34633f02131269cdcbc9978db8cdeb09f3033f0e55907433322761b7b16b75b34b15fffab291efdaf54065b3126c55d7dc66fc1b9fc976ba7bbdd9f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc45c030bfdea4dd9704d31e7a20ee8c6e78d7c063564938b54fc0de9a9254f0297b20feed5e70b8a26f761fe10a889d82881660c09525d9fea690de0654339238d7ff1f155849dbf2327125117d5ddbaa89135fc615743373ec6a8a9899060b9d0d7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcc807a6d8b59e0eec294e3eabddcea9a8e73a47adaab4e2265fd73d66d734dd6e7537990abf18869897d97faac08d4f2996cc45fc3eb4bb677a14cf2192c4258c40d60ce6ca39ff959ea9cffcc5c560793bb0347010cae08e62e5010971829c5085c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49b6adbf2966701cdfea68889f460c3caabb1803081d42e86b8c8cce1ec0e3538f56aaf39c14cf05d91aa95c476a3505b39926189388be184517fd45099c621387872420d971b16e29c96f19295f1b1bd6c43dc540b180cd24a0a555d97652e0f98f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2c93948834c7d13a2d250b220092da8d3e27b28f6ea04c3b2cc4f5dbec679529858bcc455911249104c9efd082a922355b23b2964654541b8887c452bc5c878f66a81369afdb42b63b5d6a158c4e9d25382bb03b1bfd99b26ae1d75a042d2e817565;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58e6b8762150e311ae7b8f0c454c5a90432b64feb25cd892c2a006b0cd0da3a69a4225fe5acdd4784f839129e1d29d89c1015d337cc8740b3a197a4eb06005b90a638a977c66736576659ce2709b1781b5bb5fea33eff84e9e20cf56509da2815eff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7158c728575a7dcd6802886783dc9dbc353e7413c29f6dc71c38c70f1abb7c0b01bc05e94fefdb7b57740aff0f22796857f95e9506f51938a4c00594a9164e82abdceacf1f14540788f6572d152e5ceaeae5ae1fae68f0d805ccd242ee9c6639453;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd91aa3bc64e785a70bc341344a6bac99ca52e9361f32b35a57efc02f9b0534e69fbfe21aa570ac2e7dbb11f1b76190498ef1cf40ef491ef2ec45527d89ff032fb29efd1b64a90e9f6fe3639c4b73ef9961cebd9ab807437723b0f3e96827695b670f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2a78ffef4a8bda5fb7f88883fd5c27f7f9571cbfb017c7a14220851eafe08a4074c17ab5d10d72bb27aaa7fe75bc7843b38dd78da00d28a0e57d08bdac50c8085f52180985a4a74f160c0f52e6d240c1df19d23fe8e329e2e108d7c30ccd62bb3943;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd7a2fc9525ae6c4b1c77ac511b80c3d2ec0c95d28c3118051d784895e7afb7715975db2b0a12d1064407f047f24bf402f92f0757fac169ebe96defd7e6d9edf493b0a96fd342c1a5eb42a5cc363f4c4e87d0ccdb169a220ef1fafc736fa4e947d0ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9d77c1cd06ce54691c31a922b545862b4dfdf2904618b2719610c2d479f10070f122983727d26fe0dd345d2e3a2363039a4850dfe898944139e455343c733c76d750f5a2a0371d8e7a2db7534e4443bf4164bbb061f044bd14ad42d049c2de91445c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefd5f4521ab890b13f35adaffb2a557152b3a4b748d8c22d59e73bc0013eebdf2655acb8383b11a7c7a2c65f823b4006b656437ae3c6ba34d2ed391eacc2d9d0f27c4daadf8c1a1038a87757f06e4823fc09ce628df69206346473c31d14b6f3daf5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4801f9e27bb13fd703f50078c768b4a372baa0b82a48eb5f9fd11ad4f91b9f22ed08e055cb76da397b2b5573d7d20f9fa4e485feaa9ffe88ebedc45d6c6abcddb61b437335c35f66d981d285b2be67be19e6946c9ed6eea242ae9880fb3af3c2b8bf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee7c71cd4a889709c284f7b8bb498040000a4b0e1fc1268703f1cb32304c740cb53b6b352ebc3784d7edb06adc46132ea41a3fd6dd5dfaf6aee89566a95e402c2f31103207748c9804ee42190c1cb99202bdd4fe69b5060bd29e3379de702b7694e7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5a960136416cf0d7c0d1b34421f7f11c6fc076955663c5a647e30092b34e2cc9462b4e1c746a3213c038f4f69ec7d52cfa8345acb1438f498d917a569c9a5264e22324a14a2d795600216907da899006963652e8df2e231c7f443bc49f69d7444c2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h35838a1dfa54fb26d76d9416aaf7aa919e800c86d36042d454dd025e066339e59594c238672bc6fc389bae3ccaf374450ab09c3383ccd933e21973cf7bdb6b409695426195273f5d07d8bfaf91d80463126672e2e54e03ede49a04d2b5d0c71d6ae7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h37386f5c63c0770efe4ae51f3b6fcb8d86d2495b222ad6acff9ed4200a6fc7b74fa9ee43bd9aeb63c236fca7777609fb1c1d050eb26d525bc825e588e9ac33b3588eb8e3dc5e8ed0b4a7782bbdd1d659b757c4f3c9389a7e16a0dd579bf06d849a19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h402b3af007d8164cf45df0d68432c4f3e0ada55f08a3bceaaad0746a0faa55328bda9771be115e12165d813bb424f15091219ee096f7c102eb4475d1fc154e2cbe75677a9ec9ef59801bffa79a6c2e49c89ec88ab700182d4dd9627b8f93475539af;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4fbed95ccb9bb0a4cce165de6078f6900f4293573de7c805a3e3a5a3bf573bafa4fcd6eb87dfcc572885e7371831a4b58d9c105006848fb8f7b8fdcaa5c4a035eb84800563f46f6198406355c56a7f48aa879fd96854360b7b39385f9d0c827f3696;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd71d02513bcef0ebf7c2fb44befed8d0f4c087c026f9e0513b33a74e28def9b8f518438d1e050f84002bfe2565f6d57ff74948b22ed2bc2befa383d25b53365efe36ded2adebd1384e0a41fa288a2921edf7ee059bb8c745a9a61bcfd5584738b57a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd6d3457b14304d73bf088a461a0db381bc822fc398bbb088c67cab51c3b550a598bf1e30d9c6075bc20e3f0688a56b0c60f55a4b127f02840b8522b023048dae9095f3a6d385e2dfd38805933ac533c1b237d7d43e9f6c5d322e96df0c4f45114495;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f74b062cabba5d86a4da2ca107ce38b023b885ab5ea71dbf77d41bb26129320f00f42156fb5e4428fb65e2c3088f1631f664c76daaa427c4b13c925d12b58b9c0e077e5c4abdeb2444f5778ccf5c3fe1c29b6a68fcd988ff93e4a10fd4a941d0f4d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h39cf25e3c2e6b8fb331ff108ff734b856501de7ef92223cedb0d80921c1864df654c09cc0b62505962b649d49220bb77207f504578117ad587668f55bbbff13f82e06f372ea6eeec80592e12d2fe713d5e1b3523386e72cded960b148543b8d57cbb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8798b6975c50cf50683daaed2b9f246ebb9aa4de1635d7dcc9cd2a4f0015c098b6c41fd49d9356d000d9c5275fa00466e106ff800e47d87d39ed1ead471eaf127dc98d8a7fecf9658c303902fcde64090f63fed6e41d11d25d8d2a86198d52672ff6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hefaf416de67f3c9bb3ca03dee120a5bd5cba2a510c7d7c1f7d48794cc81498ed21c09affe0a62e3c802a13d2a1c0da75557d5d4aa356972ac64266c965a254631d3477f5a1a7dcd5a3b03bd31db37dbe50149acf7adc93dd47e91eb226ceaaa47da3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3f66eadfc0dc20260186e4956efe64104b416eeaab7ba8e3356b0572dd8135d7442a3d4e4a274e8d48dfb81ab29fe4f6fe302a53ff66da4f214066d8aa467d72e5b465848518fcad4bb822c824fb8e7f157a12bd2786af1f51964952bf3814f6d0f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h17b4ee5e70ec23acabfcfe5bd60bdcce34a19ab1c2e4fbfb9d162dde3887edc1c057700a3848228e010d149db849a68f93a2af06b0bf90c7246d4730166511605c1e02956b06248600ab78ca4aab57c1ff9610aa97cf3ca28db9b859a5f21fff4d16;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2d85a72b96a59719a3c847b8d57de3b46536b076c6e852c9cf43416975cf3030e01826a54c670c89fc5985c3926ccb313b06e423b9dad2cd1cc245c7d284e2ad5020ecd684306fac5be90be4cb57d2658c1386e23504c2d96e082b0dd5640d25a19;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9955f845955643625f7613233ddfc8017f60dbf939dd8a98d268cb6990e46ab373b1cedc7833997b4baab2feb8bd52fd9c06896a5eadd4754006c7ebf4fff60460117d15b3119eccd41c072293ad658127b35fc9f0a779c2bca28a02a1a9dd655f6d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb300a4b5894fd8f76d9ad5d7f474299111e86827cf45721a815ccea0f7e4fc50d59879b0193d29dade499673f5cb76379a9359cafa0b9a1c5f1114a5e6ab6f65c17cc9bc4b6f1e17c8fbb5984f90a3aec8cfeae8be6d6f71595499f5acc62bdcedb9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee0e9db0381874a994361b9e2deeab0f555e0f91eeda018cd48afd837450bbd94a2e19409d1e6f8cecb5de6fe10d80578e0f47ea405431fe128a97e3ae8bd276aa3b103b39942fbae6bee4253f3061b70bfdc993e0df29c75c0d8f8a1bc5fc9a7c58;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6404cb7720d99f8baae1dcf2fb9aae4b8d59bd19c107fa4c7dfbbb55ad05fff560b1fdedcea2958cb3cf358b1648b22322a22a49eefb4d817c82efb700a9c75cc0e7dd8c741d2c86c65b2bd8ab04fb6be35358003a9044c4f938df0e2b30dbbf251;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h975c7afb83f405d1d9092a9fcca9f6f481c6a0bae3c79ade13d0f82416495f02926713c8f1362fc16e3b74dfdf339550f463a7be7c1563d974a48bbbad4505491ae9bf38c9b8bfa1f5e216c04f437ada450f55df626da4a8ff017cc52682d930bd08;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3a3778fe5af42b69c50e9e6681ab870710a94919dc2d559160fbc0bd3413d932d38cc894adcf62542a2874b51bdec3d0f7ae9af9e1531a078443743c113e8ad51e4bec3e8f14b0d53fc10f6d2ee142fca51c72203a0385b54780a3af51836a172864;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b2af737f410fcfdde154570febeaadcc1180b82ae4ce58a6e2f2776b8dec072e50987016a25461c56d1eccb18f542dcb919d52c3b95f9abafe1dde0594f47e4d1076c7d69b5127daa991c5c3ee22fffb5475e90331fec307e1920fc7f7baf509352;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3f6d16185dac3986ac2f8704ad079c83ec6dd5743b935f38f10f5e64ecdfbc8a28fa2b5a5c672892b72033f5d00970f5a7318e33f05b1fd511a1a955e5a199f5758d365d60e60867e937f04e4b555a83bfea4690007c882e0c5f524a8b273065d52;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h50914995bf6e96824a910dfbcd905fd1b6667741931894aaa4cd01d78757d23609bf45c72a98c58c1d0ac07ed0a5a7a6284386678a61adc92488d4bd81b1f0ee737db6251d684ec3d4d2f135b139e47ae4d0a4dc04abda429a7a4e9cb71c6e973453;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf509a30081e763fd1926f06b1e91799e097a592bd96fa3f30624d481c55524f8be193e0716c98a77492f093b5b6c02f92efa2da135a5ce08bb285cf0d4f2bef6d2223f1ce37796d8b95a68cc71bf08e6ac90731820bb2001ec374eda908a1534b803;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h97d0207e6de180ace3b24bc4536440f2caf1ea545ed0b27708479cce9d9d7872feb833caf321ed594b7c6ec721c97c1811e91e16385bceacb0fa98a53088c7869a8c8851d677dd5002869fa0a503a06f47030cecb7bc769396b2d26e1ac561ec179a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h49a6a7dd7f0f5513df38f9fb6de052189dfb8d6ea17548da2a8dbe7bd6ec835aa1d63b7e547469f53af32d1bffff911d7cbe9b4ffe75c49791dcc2c5735d362f0a4706372fa775fd35ca15473d5b9762d784e5455ed80ff42df61e64af605ffe3cea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hee3ef488fbf8f79248a76d57d9aaaada43e1201f7e6ddf879723067064a507e46ccb005471c4fb1f985f734aba90285a91a956e74ab680d543049e6f1a7017fa63c5bee03d1c660513966b4a0167886dba005d36edfd812a4ff6e559b8b33f13c3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d380c63b1c98765accede0993ee615b7bb9f3d95b9b20dabf0e7cef54ef48f52ca06797da303229bb022c6e9a34e67ede798173eafcdbd6a8eda3c77c0012152803e36a24a4d25e924cb673008a457dd80519007a70024746db5681960380c10a91;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d9775cc7fee6b2ebf74dfb0ec2a138149979e24c78694809d052e25b79d1086b7a7f2da9c7463062e03c023bf98044f4179488988aec1692765ccf82a4fd958905972b410938c43465661dcec19b329ff2edbc35c29fbfe228ce10f82c26bd30181;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h22ec6dfa3c2b64755f24c03d3ca4d9f1653acdcd10ce34bdc5200663310be58452c6eb6d13f38c2b46eea5f7da24c28bb51ef7cf0858941471f2570747ba9e6ffcd5996707a960142c921ed143f535f48dad64ffc9b017447d277f9bb0e0ebd503b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h16b9cfb0298a052f32f8ae1d276063c0e9d747ef76391601a8f98bd9ee6f0675118951c62369d395e5aed09fbd28bedeb9fe980f9c7bea4567886b4d44a4f27f03ac12a13fb9fbee64173f7c994112d59a12cf075550279e82debabca53e96b63862;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc6b480b309072b92441789e54afc61646b331ae78eb119cb08f7c326c8c01f32ba0c9d129ccd96ff06b79c8c80a52109c8422ff5229a53398166442328a735dac3dbeed5e2984f20a9ced3d122bc5ae7727fecf03ca4a965776214effe118f46d3cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32b21f7bcc029f87183d8e82c011a84f6d01e5888e38e3d341b0fc9364d69fa4561f18e494b412a22db74627201aade9b8aac10f971ce58a428bb1e935ed23e5d06bc3e644048fae7277d67870d933dfaf2774556415e817304fc4d18dd693b30d25;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h85cef193116573d7a6604e71d23fda946f7018b7251fcd399b7383f533538faa5fa67c8f91de3fe5474e5d1f841354b003eea9d693b160826322f1d5ebee7ff76cd54ab0a446b3931c968068bec5ffb05bfc49a070eed1611aa5769f44e1db32dd6e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bae32c95fe5597a0433fa5db8ccf97f1fb276af45dd99aaf970310e584b2dc91a3d371d1ee669f431d0b334c7f01c94dc5587eb4d29382e56fb78a53bdfeaacb8510c17546d39fbfdd01c84fb673b2494b9cb02ffb18d13c296ad7de7b29db79933;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4ad9bc58c9c090e2944911251b3d956a06a8c836064b5809923c31d32a237e7c2c0aa64f2e2cac933eed65b8159cefba1f815f32d87fcef598658b26eb7ebdef59418c92ed9a81de631e9eb66ae91db4c34c858646ceffd5768cd4db09af9de3b6b8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h475e90223713ff6fedc5b49e7707529ef7bb96db32e8862efcf7a9f91fc384a9de40b2ba9c42f3369ac2f1419d7779189bc5563a78ddef2b2a87a1be4c68108ba954763d330dd1f5144a6566cead5c6acf6bd61d431f80acd99b2d3871265f76cd8f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6550d95107fb37ba2e7ef95019d4d72c94351f2a700972792540856a960ff20d867255f6ea74a0a43c59cc826b5d9b5e076d7ba874acb7f43c9b3f5125a5a959149c3289323942195e25af272f3d2119ad5bde8e416410412d10aad8b729ba178a23;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab0cf50ba4cd696348bbd9aa9951a889256456be856b64675591c0096879c1f4dbb7ba681aaa80bc29f11d5914a37b110ba0912f1c8b611bcaa7ee42577433e31668e6b81f98e2ae2cb81d2f6df4bb6bb674a42746e09c73bef8a24ce93c3cdb436b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he562e4306831dfce4bcc32fb87727d19803714070fdaef1c0c63ff311d6d30060f8c564946a152b671ac9f42b33d7c58771884e333c0db6a9ffc8f9672310e31ef93e60ccdd48fc679bd8a77ea536d1a0635b41457a02e91253b14d14fb826e50163;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbf0b6e5788a4e5c87933adf3d15f4c660eb2e597d1d507a2109f7a006ba6d4d5db9f4912ba4270f086b4eeba49fe0c00939283a5b42e1c16395661d3be4715b0d4567481272865395dfa4cf7b3342ea68a3bec05f6e4e80bfb12b83209b5063bdc06;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6442bd0c7f9bb5e119cc236f6f6bc669bb3e1e363d948d8298b2f86433895949bf647d65d17cef97dd5cf3a066545c0bef052b199ed4fef0ceee85700c4a99aea6101d771114860268abcd69ab8be5d453f3ca79ada5c56820b849ad9b3a2d6c9b71;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haca7025c5261115e360e4b10702936b15d7a47854ff88deb4909671d2b98c604a96bc0c67664951bf24ad189e557c41bd020f0152b284f9f0d3ff963430928f49dd8784901ee0ce4a57212bb5d6eee1190e7ffdc832bee1ebfcae1a4f34fb0ad9160;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a15495c890e9d6ba68f030ef86824456d662754b047dcf4c84eef2dc06b0cbc7f92fc5ed03b958ff51c95081ebaf7def086ef7679e2577cba7d50828216b83cb97fe95a2a9cdcb3abf138f3e89007f0ae382b05286f35fb52f833f17497ba5c87e9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf4f08dfa8ad3ae0d2af2ae593bde6a9745c491eba94423f1b35e89187708b3bc44eac0498461489f56f5c5fb80a7630b3873069add896e1783113674f5a5d34f352dbe104522fbb3098ba21a88afd31a37f392f734eec7dee978762cf58e3933b53;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h43ed551bddd56f05e4b4ab8dfe87ea9a8b5f0e9e5856e53b8b1bdabe0118c9fbe218f7c3244db38b2aa69c1af0e51235d12d1301057017b12c128917d7373af9b9619fc058d928743cd6d6d9cc902446a7a3f07825d2f7b6a49e03485877938033e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h643f3d6fd9418fb6b2d8126a5135ed82a0b14c4c3865bca420a767c714bb6981b9110cfd8353de7d584ce10c15fbfa367e51a67d6cd3f28f569aec1bfb90c4c660ca26b5e064d09a16de6c039dd48ca193ed3d9c6549f210ad8c479b19288c88b6f8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9fc0501169df82f70b94990259a0a077a9ee34c1736caf4917bf00d6981099fc764fe277861ee81616307c9c73444728aef2627fa142aad0f5b303c43c553982232602a24ec6e056f8f165d4353a1c9d9a11ebee75a4c3b9c0c0ad086280268a5f5b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9b86131dbbabb700abc16d714f7eaf5c035ad7919500960f144841cf8c483f5bae94707fedc3c9677e45054f5d2c9dc924bfaa22fb41cfcdc0ec488087110fda11f8c75b0dcf52fd29374f333c090ca4d34a8d3a8a41dad4fef247d692ab9f55434d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1b232cda7ce671c61f084366a7f8e741c94802db6690f4e8bbc6c9bd22815fb694a356b383ff867afb600264b0afee4ed54ece913841a378c1ad8c59d78bfa4f13c953e87fa0400ba2fcff6cf8c29c3172f05828300d046e6961f06049d472df8830;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc9deb1c1f6a4a9a759ead28bb28ffa8915398a123080e4a027aee2bb7af306739a782376c5d2d6a367678aa007dffeece850c28df373e176b193fbcce6be0027bd1bdc236ab81590530a67a3895846babce6714e7bf800903e4ad8ca9d56d0994ef3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3dd714f4b6e8d10aa67eb3a107dbaaf24efc1d75043dd659fbd88052e26dfbd66702a45cc56d0273b016d35dffbb344659a652921280b003153aeb90accdeb5d06544efebaa3d22baca62044297ab7525981d31e662457adbe40de3b021dcbf6a6be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9decf87251efe22558b16a539952cc1ab0dc1b49e8c625b9d46f042f1446a5bdf6b11b0bf4af8f28d3b8321475f83a18a62c0b03ae68f740b68c0a61ad738cc60586053e0045fd1f64326fe4a31f6aebf167515c70cc25f02c27fff39c118c1adca1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2019a783b94210964aa09bb49494487623ff62145af4b418e18e83a7fbfea03da3a7100374e0cdc22d8cbd469d41124f1e8720601192fa075daea6eda4c57e0569f8086a9b16b465e3473fa8b1569d7cba541adabd77731adca7690c3b9ea60a35c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heaa2f247ddc41207dcab2f15f564780f40661271e71d1514115a621d3888a020acf71734b56a0f1232781511f80209c38b08857698ec2bf9785d6b554bbaa8eb964ccd0fe568b3889612c81b6d4808d9323f5f3266fe88e5ab470d4270d1074bafec;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3ddee6ba6d12373170942ded6180d1b3b521ce7bcc67d649826ae312847fc3c86ce33635e0b42055bbf9e0e99f18a3e8ee5d27b3b040d556495450664d3915ea690901adbf998c1093930f4775129628f749bffa822cffe47225c804f91823c555e2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7557a81d806b91bba44e6e533c70b0d17cf8a30b673923ed8a77aa82533a149a5cf138ad9ba445c443cf1d76fc5395f9006b869fd009983f6d49309a055bab695c725905d22b7d32e99f779efed11b28b813c34bc6c036107b1e0c1628ed533a3cdb;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd484dd43747ba47a89c34369b8f6fe684e92d7a1fd1c4c2edc61e1b4ca80839620fb98128fe854f2acd39eb8e4999287f7a963874d5a76f6d3c6c4efc9e529b58f48fa2c08dac66aa0814279db7efc1c1fd0a6298591e027c974c02065404581498;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h354e1a31897fb6197026c8460154e88542e1be24a17263a650d96c2c72ae49d7c94fa6c4fec7ba82a5361a9e5ef077a15289ab87b1ad765d3f3a9df34e0c6b215a80de6d0e3f8c8f99fb40ab299753a8844b72015c84b972f3da05184c50fc09de96;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7bba9d0a0590565bf2ca9a418a9637660c28ab65e1badb457fc6f17bed5c1bba7d272b6f9a6d703a8fc12d013f02367ad291259916f00ab06b307b24999fc5931dbc73a499bbfe9330a9fc56fdc20137661c64a9c1d8c660e933e070fe2e36e38483;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf18bb2c23f7f4e8aea731177983c1424f5c1185dea0521874cd988fcd94d79ac744a0fb0a1a6dd4445043ee2534ed334ef6171d63b29d39bb75a4dc992485ea5f09a3150d6604d66e2f20f4a9b08943b9df628505bf3fef9a2fe32833421ea07e97c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h882bf970292ef08c48990290ff033d2f129f52ef44939e7820dafd5d179c7a249cdcffac05509c3205c773fcbca483dcd2b9d6c649488cc7d2b40a98bdc02958f1d9ecb152c743588953d8b8dd7cde9b1ced119ea002792711354fbf8df808c73d60;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf57fc04a170337ac2caa4204e9ea2eb592577865a2366ccfdfb3684578f1f4d69210af709364fbdec2c09381dda6e400a848236d38083651c220e27900b7253c5ec93f761cbb97158902bf2525eac54d37b13bf4b8c072f541802c68a9bac57ad1a1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32248b393631d826d93987ad097231d77634580d00226381f51ac460d99cc2669b24d88d69cda1854675b27901af1c964f75affd79b08d5b694c3cec1105b7577302042940fcff5270659889addcdd85c276ba6b0b4f131b8a94f864a605b740da1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h55529f424f48299786eee130f9b8042bfbc0b60613885a6c83534b2199e5f0300a70194d0d0a15951e629dfe54a9c831cec49e0ccfeb562dc9d452dc9a63012254eae229af9cbc12ae6a253e5f65c9e4207b34b6ce40bbce80eb73d789042cacf1ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h47d17245553587702b89a3a2e33b90fc355f33bff5906cead8effe6b4733f1044377edaad443a2457e3572e2dc899d20ce71dc81a0180102a4f5f89b96b9d3fe929ec0726a785b241414c5755aea167db6e8148a3fa3c5db1ebd70515e8a7138b946;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7d676e03c574af1200bda09ed6a694ada929d99e426e610d6561b905242401ff11f135c00d3a7220501ebe085b3321bb21d68fea99f04a9b497e244d4e73c68c45fa1dea6409e30ecd5022bc619014b9f43aeb25425899489ffb223e397124a870aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he59243a0ea71a95fd66affd8149ebdf3d34cffe3eeec4af309257a015215ac7dda47273a4e2b055d376ffab53349b531290fce18d541a8cc33886b38f57cc592f8b04ddc1c50a1d944b1e40aa0fa5b9e64a75a9d2ad1b674f1342a1d9434e108d67d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58c5067ec8cfcedd743cad1fb9ee836a7618a062e0b25d514db58af21e1ad2694068e27a84b3bc1258e9cecf680dd98baae52d32d4372f376ebe06306c8ebf4d78a78af47e9b34c1190fb388eb3f481060834df11cd42ef42a50a737a5911d7d0d58;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf2304e0ec1b8d0b367697b30ef0c20d55ad526ad70ad7853eea3cafb496202e8475462730e49589834d6136b03023d743623a1989dbc3d4b0a4b947cd6db0f91bef83278e1b746c8bc9ca60044e7dee2d909480e5c2224d9f4ff3c8e93b3a213ef8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4949f4761f7af10f32b61516fc91452b817010f7e49f442d029732bef3d6eaaf25a97b5c9a98a1f2ca5cda2f78cf9a6e5075198a880548225830c9ec77590c2d4f840f78b57d95a93277d27e8244ad423ffb5d8180169e8a8786c41ea34731fdcc9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c2c1063026df3201556eba6be445cccec2cc08063e523a5101bcb7af5958e19c9389d948c620ced48abbd00a866a186ce413b9c4662ca9bc63f81953303d58f4e909ffcfc0e774942dc21bf9b867fedb91f14a9ff5b231b3a08bbbd96fba882fce9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha257204697c7ec7e51989f0d0677bafc46c1aa42b18664fd6196227d0742b42f0f31986756b562c9a41c5a721580ad182adafbf85bed04d313ee686fff77ceae0ea276f5926e6fe1cbd4082b2855eda60106f174030c0880be3e01a15dd6dd698d3b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbc5a454d16a721f5b19b096f17c6e274f13b4a8fca82a3f89f7e4b899ae4da39aa5bbccf405d8e1641c1dba8080bf9678c3334e2beb8554fa3beaed0c988928b7ec948299b97bd8555d178355b7e5aebf9de67736fb76def5d5ede22d78168190cc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h403c7b123f3e3b19763eb519c3664a5116b0768c58305fbc40255bc3c96a0f7bfc3ac3691a57a969fe774cc933f67bd4517a67e572db42b74d695f299629ca63de6c88047a14c7e2e482d49aa303d4e9143a8e56002cb5a30979e59abe9a6509b7be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc3cff362926216af22697116571bc59dccb64be231d343f87fb935ac2713bc9a8555d887051359cc570131e35b294a90646fb848712ca3394be1169859cbef4d3bc7bbaab9c5c3aafd7e7d0bd10154ac33cb25784951d2c94600e9de881dc966c2c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he09cb44d5006d09f9b19bf9ecaaeb464991630c4474146e2a9c7a63d449a72b4b4b535ad1229893a99dce5c49d1d532529ea40cf2d0269829df261fe89b1eb8e6389da3c359a1cd1af0396884482b6ca52e46d1d174278dc4177efceb11eebbebdb9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4705426a9aa9fcc157ca828772d0887808e03fc706dbe78630a7b5d041ff107c75d4ac9f6eb40a939b5061e65d4a4bd0e32e008c9f68a71f67a84141c9b9811c39f97d9fc5db32ac4740b848678ac7242210cf97f420dc8c064726b78bae686e124e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heefed85eb0d3792ae6a6ac1f2547badefd704bb56d3a7a0c1d448d936dbd738ad572ec2413220d0181aedcb05e6d6b6475d1011fc3f48f548e606d4d43bef7759837c4a035bd6df2674a9f32ccef6088b415e4e66ef75b5e62ebb24414e67627ebd4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h13a91ece66f514c529bf57b58c7ee507b0b6e1d73b860727f174f751bc2d86b05b279284fb241818964e26f2f28110596c43266ba23199451b03555ac58c5a3c22c7ccef188835e1e388235cb655f2c46e779cf6eea29eaf1bc286470b4a40b08345;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h454fed9f59a8bfd7b79300d9d304cc74efeefd3bc201c816ca00e19a3788cd84d67809c97c8bc99a38b3877d91ce8112816f1349a49a4c7a75c16159968cc47f2a5d5968dac0fa2cff6bd767ee7ce45147ab5c963c27f2f59f501d166293113d1e1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h416be2888dd7c29726694b3e2824089b2258bcbd2c575b957529e7268d088388ac35d6fb2b7c497aab77131fd352e11f2a90a1f18a5640c660cbdfc7e529eff73ea069695628ea52dbb32c556f4a900ac911cdd48afc3f8e5b35cc6cea182b266cf7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h940c5de155b67e56cc9d58b39942246f604bba42495ca9d5721eb95465a4181b8ef831432d42c0053f2fc36c1557c30c11b995f186e3831247785effe233f6a2b02167d9ccec19ea3170cd5ac843915ef14623458a47f139e5f0c0ada18fd2bdbd81;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4137db267ec2a142678950b6bc92462a907f7df0bff753df74b61fed6e5362ea29efba21e471d1a02b021870cd68eaaecc402aa2c2b4c03c1af42417eba435af4c30b8066207cba6d28573edee6f1642fad298f45005707fe5febdef3c28f5174f9a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he479d9eca2b89d7d6b4e2b1d091c3eeebdcbb058e107b936b4bc6a46174e3e9abe33fe7163d53accab59dba5e13f755ac11e1db08d4b69cbdb5beea2d5a0c185e69e1c48c7d1d2c858a43dcff9f0a24a276d36b63d38141b85cf05df51c240e6f6fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d555d93c12d180fc8a7544e2c910c0f3c0971d7b1ea8929486090f3f8333909228693fb835772806b83d595083158a73af02d56c7aac28d33d715e0ccb92a645a423895e4f5cf0803e84ebef3f991b9b2d596669134821710530e1328c63b89ef08;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hbb494761fe1f775754315c30a3c39c04e35cd65a7e88aadd1830f5951086c791564f41ff3ce94e0bf27c7a02e18c767e9fb418693789546950fbca0655b3d72c3d9555b39798244fbfc577aba9cdaa3c215a5709035e70af3e8a99151477bd511b89;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha5735f08bfd476e1d49ac870cd07de027f4048418ea1737cc85e37fae50264c6f0202546f44c93228b36a90a193e572c125e7186a3b29fb1348387dd8cf912f469f3f8032afe5413407806b72d938d3768b70e21434e51d83e04e6b3e481264ac219;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heeb4d0b38cc4701fa169b0b9c8d2b19f0762f9703ed0a38a2109c41cd51e3885016969cf72017f9de98071d8d303ccc9c0587faf7816e8fb5da8442d2c33d4341ec44506bd946d9872a4df41016eb7185b8543239f0be7012f751a40760429da858b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf749b6d716bcddb0ec99fd7a5413477085b77abaa1af10425ea2244fc0115da445f228d6fd157b859bd3db2a05bb73317a992ce61bb35b7c6669fa67ebb97cea4b188c7505684d08204ea804b98cc31d5d3172f875c45fb64bb05bdddbaeefe29d98;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9f8378cf8e8143711542db8a6f451e4b8e654bab05d973f2f6ed7af29ffd0177380b097e7080d59fa9c0e28637347f3dabbde73138faab9f9e0b41fc5a693919566717e140aa6a10e361daee896b9d85cabd6c440306537359ab2d636775e0bb1c94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdf9030d5dfc92ef53ec43730660a1dd00252db746de3bc2cf12255c36f39417051b183968b61a2cb42b4e5fd2d6787e1894b1aadbe9478246762779fa5831a8b30293900c83cc935bd694bf19078bebc28ff1ecb5d192e1e47675f71ba4a8effc74e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h76d498791822d7f46db1d523080422d23f6d41269c9a300c2a2a9f400f0f3937b7050f38e260f83d7b238f63468ecf152e42a88302214d08bed34bbbaaad474149e6b37de5baa8885284d0ba9a7aaa5cec6b6ec217d3b4ff7a37c2d429a61546fbd9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h54e2f40e9fd7e966c4b261eeea9ecfd2144d10b3ac5ef2739be66b31170dfcee21a2849d9a845a525439335361e57bb88b33075e565f3d0e0842d728f09a5270c1580e70896072960b7fcf196d4198c233afae8dd0936dface2ae5d01439d82571fe;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d72a1e664a2d4cefddf9c653907b0df0d48675df29a902eabd0f018d5a18c60e602a72eb9fce59f3f176df739450cf1074e8352721d7bf4959012da230a71170116e5f334fcde57fe436fb8d76c83db3447f6e72d8aa92fc1843c7d7cb04cfc67b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58b42c5b7b7ce8639136b2ee2f2a84db2630c017b9366170b77144ff2a0a1e1202dc59b8139af1e8e7431b5df054a5aae826ab58b1afa84e725c214911420344ad2ab0be0b1636e4011049b0bb485505e160c9486a8e705ce7dbccd7e7b29987f6e1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f696875a707ef080cc8a81d4f564de4bc1ed8e8f5125b5ec3eb324c412e97f0e97854667ce92376bc67da710b7fc8d1ab665aa6185f25b126c9b4b2c56781b5c212737b1638c46f76b218391913ee5d457b5918673adb886983b73ee6386d7ac200;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7a0971f0ce5352aacd1b895dcd0301a2bccf34c02a39b1a321f7a4068af52bcd95ebc9ce6f9eb45c6d684b63512c39002f0f30d671c6693778e506ff5ad631d14979fa98e0cf93aa299e925aa7241b7f540efc1a3818ecfcc72d326de27db40a1bc4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h20f1bc267f34c5b4a03c6ec065d0f561745e13a2fccb3ab73a5a7b6a22c80f4153536f7834a8ad09b027b49b6f8f6d90576825a91fa32c2bcf974672d4255e076bdae7dd4acfe33a09dcd12882902b37449696b3bb5024ade5eaed5165a6f746b3d4;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6faf5fac092c575dbf616d056551b958c19fb46c80a22ddb13dc8873adbb285609f003d74650b7b2c1ce0845ab0df6d180b762ab83ff124a409b451f315aaf64bb8b1760832a4df757cf2bdaa10192f695f34d95557810b13457886a7346cdd38bc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2aa0a8aae07b642eab0765e85fbe5e3dc85c7719a86656341274d104b133497d8f682574604db7a4a341e647ff2866cb420cff63d85172a95fab2bf7b6ed7196b60ac4f884acc76ef1339f103946ee1c6244dbaf8b9145f12ab27d56fcd458e80d62;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfe55491edfdf394dcbb419d521fedba795df68c0ef3d722fdec10546c9439649fef9a554bb08d3ab8a27fc73fcf1fa0c6170add3a9183f7f04cbca5c141de0c9ee3757f1362adadf8510aea4c9bd87d24710be4486d266f49486105966038a0fdfdd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h95d4e1b5d76be8c05b0c49826aa0d9def419d4b04d46460af806c4ffadb0d1c0b6cf74a8d5d1e3910c1ea8ea393a459916040751c0b196d0d63681ec621e6ccf2255ece2508c3fa592b0b27d52792b30704bd5811b4be1ab64ba7aaa0ac9d0a83056;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h604740c63452848c9e7f34005c4885bdde6885178dc4c3664077fa4cda388c5017dba327660a3eceaae877f72060f3fe612a3d43e7d3c20716e58699efc8569a38a54651eedad9bbdde512654223016cfd01d48aad195d41568040bf2a998a75022f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h64c16c0921801268521d80e3275a3ac89f3f0b17a46773a0154886f6b4f38eb7e05ee9a51a49d26e8e49d002a62d1432d7eb836e4cc9537f7139b87f1f16fdef1f0712d1de1403fa4af93642d1f613312af940b4825c3af696cfdc3c91e77aef533d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h32ae3734eccfac4730dd49fe803023dbd09845243ff100aca38b043eff4262667c77f14af6d03e50ca05faf34ec9267a1cebe36f887a28cae7acfa6ad56c0c913fe5e9aaf5c5c5d0be74bfc9c4f9aee8e68e83765cf78cec65f7429dfe510b28326e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4953d84a6a595f381d712fe95130d8f143d8adc3935af2dc6f75285a6fd131fca0fb585c6d603a7131e47c6b95127bcd00b8f1fdfd10688ceb02a0d73d9cb36c0a7cc7357644c67523f28a4b5deb6515ef3990e246dda05caedc9fd28ee4d60d3cea;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h23af3c09bb97dc9630128843dcd5b7ff0aab96d2081d60a3b86c292bca71bd1a04cdaf09022ef5119d61e17f5e82eac457b8232ce7cba4d3b2e9fe6d65d71ed5020a25f8d7dd1edeaeaf8ed621c6b7952624613797593b4909460bb0c3d45c83ae62;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdfd0df6f3a62b65426c0ffc8fdde3a4157fc4ce8a86296ff8c8156e27235890d321335993652bae20035e08ce7374358d4886605d5f024f3e463f03084d71778021e07dce3aa4324948f791218f873d2a2cd00af40d820ca1de98de49c8b72001d85;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca2f56b11a9c4d44221a6ee85a2982e19dcaf7ca87e88222663a54b1e02eba4cbbc1407eb476bdf6731bf0fe48c873e5d256d7636da6e84a5afd730bb8b27d16334eefe9b7a845651296fb0a55ab006a0b7cfd9720db01ea1b9f55aa90b73cd84d42;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he269333754dd1a780a20e2ef23dd8e494340ebc72672af1c7706c7c5efc21098279c9cffc1d13402fa38ff49e7983bc7c60113a090fe3e7484472df89a05b207170f30548048ff26e45c520880d7d333b8f505fb863d972a29fd3bdb9aaf5d369650;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he7fd8d9ca81db1870ec2e9ed7c783fa03addc3644469ff35fb608b58ead9f9982952a5c600d1596ffcc8fb61853d474b71ae1bd8f4ed7b44474ef09d51846f3c41abb86739b47af6d1c1e1d9d46a8423d08caf600dc3ab435d16aa84c7e0b39a1945;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc304463ade86c68987097228b2fade58dbb3e2d92c86233ef4e4de5c562840dca7eec5f81aec660da20658dd7d6a645468f05a500544cc1ef451d040051c0ab90d8c33458dbbb72fb940cdcf692b6a5826baaeabf0f2ebaefdaab34549dac23e51ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7c9ed8be3271005261328071b0f759d48f2031a981ccc4f13a2de4e89e1a44a45c982b1fd1eccc3b234fb09516b343d95674215f77a93a565934689262f727e780049eaa673dc0fd4d187cc4aea83d7274f54cf4193d9b184e9f0e8e8043350396e5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h36bc1877c3f9e3332c9cf347bef6ce10a1c7c407a1e260ef21957991b9295ea69ef4285e0e39f8404966e702b3c35c937b5edae03fcabf47fdaeae5b66bd3ea4603cd4106ee49d9571dc2454731f1ee4dfa09d51503bf48f9a30196e91afa00e577a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80e5c11b88cb3278da9feb12aba03c9b3a2d8728af55684bcf7e1703f6487055f8ef23988c7524e67ec56b71c757fa98c8e9b51b994085f276059ed273f596071d66717214ba519b02f3d9eb51dfb4b1bc4a976a06b9f821512401ef30e98c0fd1b6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h146a65460f7bfee935c4d4bfdddd3e876ae0eeeb4d74ab8ef514c2e97a42e51b29cd83e74f72e0171ecfc28b14c48889a2066cbc76b840448262588fc5ca7b9848b92fbece4a987a8dd568828345274aac0ec6de41e213551aa1ace74062ec48b272;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h603a026d6c8413b9fb70ecfc5d1bc6500bf79537e8aaf69bb5b7296d689883c7e719ebdc4f0c4ac0abdf5e8acbc208a1e7ed16f0d1f9a37b3017cae16e8aa53a2c4ad579fc507a0d9c8f09e50968026b54395f50eb4a5882cd53b10f9becf577bced;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he44cdfc630fb28d4a50cb67a3e4315e9a69d0845d52957e1d94a67b9dad192de0df8a3dc0dda1f21acdd5cb292208ea112cd2c610e16fa6ef45a4da008f0901c3b2ef149d05c3e8fbf60cd0f0a5ef9abe716a3c5fd0464835ac6de10e040f84fbca1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4b12e8e8ebf7b9d00d29d849348161751620a39be9b900bd7c9211b7e2d4a1792b5fc8023c005e26e389a5afd80b843a069aaf41cab7b180e2ae471ecb67b8541525044a0fd060dc59034fd92d987e22f420935933f8d6902c5090779026778cff6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd45da5273c3f374a7e0d03ef17b7cc3e06f6369968adee4e32bad20327fef4c297aae67d5704693a8994797049cea50dcab868232eec1f414bd010e964a675284e378e2aae4783bfda09894b8a9c299e07852d7f8a5a0838cc5425378fc30948c142;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h42312cc0e9556b8dcb570208011135b81ceededbd6b4cc9d565cd54256f3f7436fa9a3da64185460b647503669d1131aed869652fd14bf95529653f9803d76d8f6b5674e399a957190841955ed144c46f2dcc9dc76d62770c4e702d123bc4606cdc8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hba6ceeb55061da294480df831e798fa60947ee9c4922793e45dc3a980fc7f0be5ffc92041d959366b2db427fb5d8d623edb27134ec5cc2c9cb3cb9eeebde080f676b3006f8aecc8fcf24f66c633070644c60567e209c19faf40d902a2ae0f39fb5b5;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9192deb56fd1293ae5488ab11b83cb1a004d5124d8cfde9b66053fd49aed05396c10e635aaeb8cfd3421a5443f2441a960334e8c23d81d0afbf855e527dff2648d62267ba38e0abc9da8a0c78d159cfc5023d060256d8a3c3b7e152798aeb2efb68;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he12f53eaaae2b1e472f3c9a7a9b2658297903bf83b73a48c600f3c00419d359c204644490c4d0658c0e23623fcd786046a5bc68bcc94aebb8692dd1572e4e96b3e45dcf018271ede0008b3d91cb1b67c68a3acb9174cdd46e1c5ebc8ab83566a075c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1978ae12a5ce602634f17341f863f1146ebe2739652ced1c85110b44344e4cb8dbab6571d3b8654938a14f7e0b3eedd4b46387bc3f12dfc46c7e4207284dc48fbfaa02e90328cc4eb1bbf411710d72049eb12aec886914769f60f705b76e3d7a0c7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3c03138dcae4a32b43f797d56cba0da3d55a439975ed4e7225414d39077de588fe67e63c604a7c67624e87499fb3eeea6d446541e94a61be4f45a7ef0dd5ad84f2a0d6c7f2a7c70dea30e1573f188da787002effb398a976b30a50ee94002f637bf9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc4ac0c45dca9af6e7b51afd9d621a2d98856520f3ce1b36161c4d63757031662bef054284de9f1b81b6876ef84eb3eccb0038ca2c42c19ef889bbefa527053e9a04d054862ecd6dd3f76e11f2188fb0049eda02e2e1d461d481da949e59f4d2c0769;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9622cfafcadcd4b72f58e22c73349345289170e137b52095791ccfb47894f50f73816fa6f8e2f42e20eb49ce221568e1b7cdbb0a8ac4a4393ad456fa46a5b82416a510ca9d8a38dd81e1cac0281601edc67bb377f13fa7e618ea58bb4be095ca5fb2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75df86354e4c7b5e1367cc4a9d6d5d91c060d25292da227b8917fb8af30ca34bc9b89545a3a102e07a8cfcfa1cd64e590dd8ef661bb9296371b348ce65118b90f1a4baa905f1fd86dd9eab93437651b065e4f6b0915862a1976b6b65373f80c71fb6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h142b0f57c6c2032c5dceccd688b9782fbb5c858370ca6e13e32b1fa5f371f7f0b972fee8e6c6e5ff678f5764cb7ea673708773555912962e40fd375c6348becc7d272a2e8eb32802a421a9785ad6776144751b2bf6e4312c03e8a10f36e04c5a0bcd;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9e23ffc8c85c674f9aafcd59f10807894188d50d2a1dc01f8a113e5388f3017d261187a82b234fedec9bffde3c19dc3ecdf56d371c8f5ab27e8b8b724abb1ee3e336717a1e8f49967f87010d13ce51cd1f21495b5093b77a7d366624105b5c32b94e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7954924bdaca4f0505a3d5495bb785ab024c8c60ba606bd6fd957215a7c44cddd620e4e54ea17fe3b97c8b27068de6deddf577362c0ce01c163dc6a144dbd33d8f4d0f3daaad6bf24df0ddba140b0253558eed9528e7b4a372bc6a17f0c4ed526487;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he3009533ad56a4aa368a009591c2788de3ebec74343ca0cfbbd74b0c139bcf5af35dc95bea2c5b0e0d198a2259023279726981073154e7ba73b0f289edfba55c7a0bf7fbbe6fe040ddbb19e96fbda3254c4fd27f63170d99f01b25ba9c92a86a2427;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heaeb4238b89926049033bfbab5b7947525d7aeb649f01377277eb070ce829a606880df025ae0256a8741b14e401434e9a9d4137529da0b48c8e5155cccbd821e27f2b1701b9465b8067899ffce69df7f4782906884bd314d00ffad7fa56d67449c40;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27862760f734e4a1c23b51c20da8c44f992feacd8a22638b21e541e2ac4ccb6a771e79a26c97d65ef9f080ccaf4a0f6342c1bee80acb7a6cbde6881a3f37458e7d3b725b63f61df89edb7e1ccfcd9a8887ed371043cea477c529aa58de1964c8d35a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfab127f49fc2833135b28a410d1ff60c6214a7590625a9b12e2df6bec5eb5e19a4582e9e3acce0eb6339aa90d82feaf32478ca60e40b360047b52cd0f236f3a4651e85002e0a3c05748e308b49b6097dad498fbc95d2e0887f12d8f28dddc746b13f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8d4ccd47cd8b3f3cd64dbad6dae5e56a89637b8daa2221d73b9971793b514299cc6ba8c516d67ddce110323b4d4a67ab3704a2dd0df79bbea0a4d1a8b3b8fea5111bc6ba62a6697831f1c3620ca45e0f2bb22cf28e475ad94151de13e8babd80215;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h482e341accf7e3f80a56d4d36d98e023d8a1f51e70191d40dfa847ce2d5de95dc5726d55032ac94a24d241ba26ff8c3ad17664e77eeb4c870d60cc70b8268f7d93ce76c3178af7c1106db6f8d63e567b98de0b48c0946d4006ccc4a4144b4b3ae5d7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7421dc8b197c19e14eda592d989bde3344ad43365eb32b688b4e216dad7b9f91915d5c583f44224792e99ce57b4bbbc67678b9a367a0b5ce03fdd341cdec965c6f39f0bfb0bec6a210b2852095dea74cfc2893c8f6f85a329784e75ef309734ccf11;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hac7547cedb4f87d7b103bc310c0c17907aa7a378badccb02b087f79c38a1fb320783774f6fab1502e866f9c2cc812bb6476fc36b98355043f2d1b1a92f65def6b98f11be5c54084045e94a53fc69d6e0e68621f02a74cc8cbbfde65eedb49520d4b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h960337664e31b3a563814e79136c48040c41ef7108929da7bda4718b5d50407c222ca6e78d44bd774a53ab22bd31d1aff61c4fc66bb2f2ab31ea43ec24bdf933ee1885d3c27246cdaeea07813a084b809b229eceea67f5dd5ebfaeab527372673240;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h986d2518788179ec309acca5967b01aa124f5afa1dacb58543cb244e31fd4a8b762347d5e067b8c5f1f333fd9afb82a6fc6593535ecad85ccb51f88cfa128775ce132eabac0c768875188eaba8d8f6c50376178572846d26f3cf5430b1a54a51be63;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h67ac5ec7b5629e907ee51a0e8d2c608e6b78e0c5b08d217b4ca0ea43ce8c24f0e28b08abba4931e8dd774ccc380f77bef61fe1295ed605eba58b6a6fa94429e90649e1afff01210a3b23fb5907078c66f82cff570608fa7cc0c0e38f6fb695f55a94;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd3ec63ab7c644b8f9cb1a79d9a5312b8229a1c33eb34b609faea7180c6e5aba8a63797bbf61d13b7e65d8245012e1fa0f89f1b94542120f49087398712e8626c0c63be9a99ebd50855dfb6dd663cb8754da43d1091697f5ab84c94efe0ee6c55b734;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h40fc759e08739c5509d3248755f9c87b95a502821f3ec6073f119ef0f8bb942ec39b8173d98d6a8f3894d882efe52822e19c6a94ec9dfe10bfce25c13539f5b151298d739b1fb0b57606e5791b2e4dd0d153925a3602355a3b896bcb0757ab548f55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4cee7a3ff3159d29961fba5e77be4716bf40a0080aedac26423a08cc18aaee357f49a1d0eee7da92835eef91e3909e6b575e54106823723c4e58548450b44badaad42622bf69bda581df5050986e61ad546d7178b2000a15231ebe4c6e1fe9e2828a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h41aa83ad9004a801ddf3e6d540bdc1fafd5cf5efd8bd8c21e14e9bae3d2bfc5b21bdd66c8c043427dd5e94281628eb9d9c6ba5087db1b8f2a081ac1372b8ea2e2b8885df146f331a07443c39837ab52f565756d82039608f985d6661a293533f6006;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hec8c08611d96f97f0d6a3a6a0aae5f94b991c5873b96767bedb27781374cbb2384878052dde2bd2a67043933f94d2ad4e072592f79b16250fb45f9e0348dce70981f4dcae76768a995f7dcdf5f30bc9be15fdc0eda585ad70bd000ed0d7ab7f308f3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'heb2967ef5d89d090159b54910b7316ea5dddcc9979a015b4b9bd981746f074a32de77d1a25ac7a792dc14772084d12217d1f2ef55120980cfb0027bd7867d57c2489060684e6fd2f8f051ad72176dbdac4e3e2adb1ae7d75310f7005584d9c27e448;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb040f7de998bdca86127d22d6c53a79ece43853025fc59755092a339ea91654596d5c5683a29e3ef7acef33e2211d1487a22d4b87827caeb28fb0f8f3c440e9c4a2ee3fd3e644467bb9dd66d4e43b21437462d51403d2a648d41931bc50895768ed8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h399d7196b459805484d642027fc4e11ca163997651a15a99aca65b7af3beb3c0c6d1103efdced29ab5e5b98d428838de14c1ea4ab8f9dff07e684ed8fa1dbed25c0f21f888f4cbce810962c2b2be5d665e5bc0049dbb3c5502827fab700dcb7b5371;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he135d00ffff05061b1b2ba890e916e7aeccfb9e71aa105869d4d4c5896d923ceabb7afd69ec724949c4448ce70e6306a8804ab3574661c3acd76004c941f1bb2056f51756f4255384ab64a5d67fa38a0f1f2b4141a239345fcc0d7b2e3043cbcce2f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4add4a7c93990d94e3b3092a695efea13174dd8201268d78190d1599b8c4a203addb85053bdb055ff3167499ebddb76a348864e268b3df68514bad2da715992b30837ba7ce0518fa7b52cf7bdd00d636267d35e1ed2f0619cb9a12ece205a5603b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2b3b72b1dcdb0ac21e1fd2422a22225ec21f048932331b895e6c6c380b735b5f9fa1578264aea6e4b64cb89c3c700f8ea767ebb7039125f95f9ed10b6c5b3eb480b0f1163c71025aaf20de357608ee7a36845337dd36c39fdb0ebc8c260af282b5c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd0fa69e5a5158f32b42237c56062e1a9719566075df79d965dfad9d37c0e3647d0711875e87d3eb5f3dd4a16c3c5d65465fc7dcf3f9f004416fe228bb6b60c3a86a9c398d02fba7a6673b84a0a619f4eb8d6053facf16c7f3e39b0acfdef81ba2c16;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfda70cfee91c67d7cc8e20ea92f504c1b31e8287510dd28e7e217bd41df256e4138ac5f006a3cece593976060bb9108daff29a1e99be3d67d2dffdbc8e694338fb0a0c0c763910b258d3fd923b6b4961dbc7268b89d3ca3dbeb61167fb365bf068d9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb0a89f336f7847bf1c29581fe9b89836a21b426c4bc26e21d599ab7b171cafc1ce165d73a433fff707f899341d0413c8da628563c2d307a457796277d8516f6cddbe40f2c54ee88562a071f22f7de7865257aa968e5501c4577bc557c840d75c0915;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfacc43206b4db1a96885e66778b8e5fbfeb4bca472a8c005a4796abca6ed791f68efe8c611b18a8ba90860e0293bab46ff1891402304f7512eb8abfbad4fa6e419e48faf642b96b85a544434adba1045166c274ccb83e322c553941944940a699f3c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8f9ccd6e6ee2ce7d2f3b759098a56bc2c75645aba7947348ef23d5435853e0d434e67f73b37cae9bfc5a39be378cb92d300642dfffb21972a4f45d68c12a22840a52c8e4d794751e3f4ac7c3978b420850e51f00d8775a2d373492f68817cbb06b4e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf8829ced41520e50cee1e5b4d3493ac9ab3cafbebea079e98a7014b7a7fc0d57ee013fdae9189ef6d4dd7675cd2c7b60c85651ae6c946099ee5037dbe986919b6584c450f24831bfc58cac3ed8b7cf1d4e28b549d301b1ba39fefbd8e37f3224081;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h26d83a2fe5b6ed2fe1a22b6f319f0f2a18ea4d393596e9c38b9512acf9da5bd0f0caddacabf3b49cac53f12c21b8568a2f51b3ee99f2bb0562dc8900504d1a72f033ce89cad1ad134cfd3582045dc9431c2c71eb78da80f15dc3271aa69ff7317d1c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h336eee604277282228122b79cd2805cf4a04cc84170fbdc6964280fdf0ae44dffd73d28604044368b698763db6eb452b8e7cc9938f3a41561b3013f905fa50c003e3c7878e0c4aaeb11ba841ba843315d055b69e5090139e11299e6935b2e015475d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8b103bd04ba153119ab4cc7dee225e357b28559df2cf60debdfd6066535574bb6d3ceb74d505486c84b137cad4f8ae9559dec4d8a50473386720f4b222c7910b16fa678e8f2794797e98cd849ba7cc97b61f4d80ebbb30d0112f8bbd58ff29f43137;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hdd4f0ff24d8e2654de79d5bbd4b740680e3d85eb252066120d2b5de96214b6d1b145fdf489b776c6444f80aabfc7e3fba575804cb4e2cecc1b233dcf2e71ef48eb12bdeea14d9279e119ab14ed05784536d2cb7794102dece257dad4dda0a2439eed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h72f95adecd6bbfed65c17d6fa5f6b5f0b3a26ad00dc1ddda2b08532c46f32e9429c9184d9f3805a7d17e2f8eb07bd259cc0436d54bae220fc49efb094147946c571006e96bd51ed6a91d14793a92491a0897e16a4a1462c7e0251ede04fbdb0b06ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h69a1a72d93ebccd31bc75fecbb0faa9797fc09a7f3d1a7731dce1df42f088c5a6d34f07d5063ff4e1ab9023bc7252942a8679228c9767a4c686105534119cb1d658af089f8f68dedbf47c4dadc12a1b09deba301732fae9d68270201bdc517ce8463;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf7f8ec2f8275158ccbde8c8d019eb33fd52c36cddc7e0846c4e9da94c2557da8544d3b07a7453eb1ae9431f16ade6a9a0f6d94804992ee4c1cb2d68c61378b0d754f97bf69b5805f88afd6553f7ce8b8dd242585c0d797eb6fe9b9e4a2a5d231d4ad;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h58058278d58bec4c451cb5e1a1bafb1dbc15055f289e9347bdfeaa8198f51d635b67cc11ccaad9d58427394601c608deea2b8048060c2d9f8f461957bbbfc496aea87ca3c1eb7eda3397712dcc9b55d51aafdf532a4f70ac0b595d1d05a24604e292;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1eecec247a0c70d13ccc5c94a67642854c3866a8fbae8f044f5e9dd760788c8701bcea74ec8c3ff9b49279e53ecc5e368ff6648e6c4838bb1ec654185dc86859f254b4e8e6a2d0b8f4cf48df23c94817622564cd4b26876b6cefc9dd20c3c6df637b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha048431cce294292a5f7c7914906fe5ffce666bb568d43a4194080d2c0ed9b78c0fc08ebfeb98ce30a7c89686fd121bb16972edb261f6b60d394f17f9cc735844b5c6d60271a5b27f93c5713ad5b62722255c060f49d8ceafaf1473c2ccc42f3752c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc63fee24eb079d3a23adf20bc8a8fdf3e56b40157b10c5f382e0c352a2d2e5a0f5e500bc2957d6f6a7754fb3dfd83975cc8c8d2587cd2954d1f0d9759015c6587d88844bc120626a7bc09eab3df0fd01790d1c107936691bb2d57cc07099816b37ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h769e09ace81560008fd97c63afddc97d7df757a48dbf99d8981b898ce5d343eccac51977286f8f36198942f2baacf0dbf4d073d259186ff0cf6cdc72a47e12f22ace4a822ed33efdd3d1ecccb638d9c9385f3075a5bf5259fbe71f20fbdbc015282f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h51056b02c2477efa9b029f4b78a872cfc77e4ed9f97bed04f91b02db46b2482769b28df76df572834696dcdddd9ecfbf5dd5e1b1848ab85822665c6a2297b4a5bf7b1a77ede7d3a93df615f96ef637eed14624054df078a4a81c9e5569a1be89e579;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4863b8126803b2546e59c00be7ff043628d925ee250005f8778541dc9ed12614743af01873757bb1abc3931b6323de0be3748b18052eb1b0bea1c827348f95a249d372056911880dbf145642516cb7df0ba07d624b85f6d5d21b2b2b9623da2394b2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hab741861e187e114306350c305a06cc29efc30ebd1fda084e40cf979ec519e9a9cffdea67515d677d6755c2c2fa47187fcc56f7be0b1466b729d9683fe2e958d021147c656d643cbb1047f20ca7ed86bbf05c4e0f544d979a97237a47741ccb543ed;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd9acb91d7864f57eb44bb3f010031fcaba1f7ad4da24be1e895178ed79de844191bd521bac149dfc592735067f608f3a9bbea66aa3d7b9c932d88cd450d73d9d284a26879187d2a712f1c8d1e32d28dbbbaf8a5928dc83c4b95816594c13be436f33;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h84f9597eda079e3989e20553be0a84735d34729328df6ff77486e6d5eaee2d644be0e637cb9f981f408dbe1dcfe943f541b6bd3c4165e2e0d5afc778ec33944c46fb56c5c8daee612083cb2ceb3682e280f5ec0c0c63a230e60a8f193b1701a206f7;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h80101ad89a7d294f35bc29fae0ea0a8b484111adfc5cfcd2ee639d3728504761002efca729b38c4062bbde90207c8da0b064bcafb1b3bcf9c1b7f164dcddffeb311f1ad9fc5854f6c62faedb6d646f7d6ef4518365c6d418e4de2dbd9f092d6f330b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d92d531ce019013148f16f1debfc18428b897cf02b0f211099ba52adebab86df42310633eb801d6f15a79d2f83793a97d232a9f619ef8475720f24bdb2ea644173d1837897fbd1050b5062e0a959352c5b090c4e19911875cdd65cc271cf7112d6a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he6860cf4b17a75dcf6fa9503ce90ad334722512f47056ef9c14f4a64d49c2c8da00b01e22487b808c5a93b957ff8865981dc3373c6d60cf9dcd6aa95ed9b83ba443ad688c3b7e9154fe80e146b3940d8b62eb115121fefd777a464f2c1be5060ed34;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3d9fec141634ea7db5a464dadbcb0c66ec0e3abcafc558e232beb5a2d4016286240b59c3ceb03503ae3916e1b8c12d6d662ea735ada01fbe0c6f57762adb85fa1c4d57a9b9b5c481d40ecb5ed8ada7ce2bca4ac09fdf11e5e912f4f967a1addab3ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6fe888f7b3801b17d16bb34a8f5c4c573ac48c4966c4a27d8ce4ed705be59a54e97f6f15e6fd64b0cb240b9f0cdbfaeef1cc78133c8084089855a853e2beb6e5f515d63a6ad422ec34e59f1bda36fc392f45dc4955095b8547d1f147cf04b6b1b569;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf53b8da47d0a905e1f7ef11b73aa905b84206bc08fb7ef11e3cb3d1c2b83b3d648898568f65610be766b7d75ecf8ca1599468a887f1db733a0f2c9a1be0980cedb00be0d1bf842ec82358cf2d6e66e952992af5ec61d9f5769d98236492e21acad97;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6479cd191f0d39d6cfc9592a663b348eecf4841c57a5aea595c005268d124ef9eb80f0d6f006e87bdce9a7ebf8aaa2579d2c6fe826a9d125414b031a8a962f11855f7fdff960f01d58feca7f3e1e569d62a2ed0b134ac1544a6ec92d7544cdf53fc9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hca904957f44cbeb18b7e444a671d5ce44f2bb613cd6eeb6e86b64e2200ed7e723d502cc0e0cdfe15087bcc118dafb8e5a88b1e8324e7970c4ffc68a02bbdeb5386b044fe8a43cc0c7a7902a05ed6cf4d696d0c9a5856811b2702062b344b94088bf6;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he35e5e412d07b30459565c68a3a97d0e351a86ec5e95699e96d959a7998271801c93f66ca8af85a0148967aad738e05d9c714a502109e971a6dff2665e1f30774e4d459a6f5c15be3bf2052aa3853e26ea829cd4bfefa5854bfdc5f16d7d21ec8659;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h75216485eac82891915449ca4e1412e998d2b3a0439dd08b8dbe0c445a185be4d9d97b2ac5498de9ae0784e0fcc0673937408422ffc0902ac00cd0db381518fcf025ff0c374edf337633ced5a0947c85811e6a7175e2ed56b5d4f1e61393a507cf7a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4e000004de57ab4715af45b337fcee2b472b25a5851841acec678abb60b527d994a8b642eb6bd315d25e2d72f0cf9db317cfe3b130987b30ca7bfdf33118af18c7db72916d1311b3db1ed86b1e529cbddb64960504c614e4e9fa0cbc4facc09d7ade;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h408234a646217c1b6f5b70719018c17f0fc84b008df805d19b90d917cb8ffa53dc519a37b5bcacb65b6932139408c94803864d982acf92eaf117a95053ee5c7522b16923590a8c233f75c7cbd4ba0ff88c0d96383db3dc24c4e3ec9287f52c179e2c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc52417d7253338939aabb9e47fa3f4a06e3487c801d88dffa9669524af02dbed8bfcf49e7a96a57367f6b0c9edb3f3aae86b55f95a90d0f98e0829fe0bb5cef873e4fb6c6830cc98edb746229bae05331919401b4924b13d28e8707c22ba0a50a4e8;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h868cc0e9a759a589fa2ac7ca10799eda6d3fee4a317a87a049e362d55c5a97240d43ceae1fb7a9907b799e686e8322be29701a8dce8095866fb74c53866291d8edefa099dbab087879273d6c863fd09daefb0a78c976781a42719bff07c4f6c8120e;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha78abe63220890bc015abd162fd2964541189c363d1ea4a279130e7d2605f9dff2eaa1f4015f84b3f09398ad4e461732c02c81f26df9f069f9ea5850be7f7f89cd01dec38126bc333058486f7d2c13c55ec354f3ccf9d512834680fae82d6fe9694d;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc66fb47a948cf44ef8be88a570f4936f4dee9c6cfa4abaa6aff7e85154a851580a16334319cad7169491cffb828d9c523c916afe75c298828e213d2fa05ee7d1e1941903689331f77505dd0e543cf6d63d6b8b5746c5285eeb2c135ab5abe7d3302b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hce00171dceef2ad6d14dc3dcc3c75f792c601d728546c1ff8f2afa601e068d0343f4576987db509bbb7ee25c9c2092aa896132116a31d3e776ec664a1333b74e2815eb8792c7ebef181093a508163c8c26b6ad293ee47afa71007125474735410fc;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h61aa03b7288f1133a9c18622f86063b9809bfb200d9e64d22ecd71dae1bb46451c7882f403f5a608344697a20ea0e00c3853460309fc28afdaa2551d180361b7c32605353926f329e874d2d0d26c638da870882df9943729972c90caf38ba61bfc78;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7b1c5df66cf121562c15dc4df709b955c43a64e88eb919c58a71768daa82e8496b8d9f678f2b8fc06e3e5505822ab56087f9bf41f6c593eb0ee56dd8e6991990eafd4b768c314275d93276a3a618aa0230591c4f447f321209b52e10f328d4b8f2b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h83952142f270176dc4f379f9818b41e43a3a5efe4fbeaab6bebb56da71893ccc123aad7a120c4c74382967afd159782cf5a4be7605de041159540ae2b79ba9e9507c3eec15c09aeaa8baf4d690e80472e270428afdbdce1602b1263368d27873c3e9;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb00d14ff29f1ac71a19c46fcdb1fff8c0e003c7fbf55f90f28d1bcd2014db2fd402c3cdb486e7fb3fe1ef3e4ac4b854ca1704413dbcac80eba0b02afd82ef01e1b2976ec80b4a0c0ecfe2e9a1c0209798ba260e7a729215360190d3f84b7f05b9780;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h8a31c52ea002bfceea36a501a7844079fe35e928c172534a1ff2728f531be369495be740b976622943c99533a8b705414a8305baf8257a44b118e485e883ed742f72bf86f94f9891ea79f67f9707fd9527a2a08ffb935b8c154125a7a1f125097444;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hda96cccabc672eb0888cae9e491514e2bbfe684b38ffb9db1cc9305563a146ff094984e2ad3ae54f70ef4035f3e057be0a508cfe18d843ee494758f302b9ac2f343079c0b2d100c6f9b1f048d955f8e56a58b49890f3c5fa29d4433cbec4eb7d34cf;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7ac2d6df82c85ff92fd1dd6f9c86d0257cfb693d6452b95c02d26ed94ee90118765d7e2c7ebfc0a02cc13687c70eda5fa4aeaf0e756efe6ffa2ab3af9d4700db1a093602fb9b0eb5d35f4ca12e6358ce4392c59ea679bf773d2f13671844ce26755c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf2af6c43227a8c46c1f9f0ba6b5c9ce5b6f0234daf8ac7d4f15b596efcd4a61b95654bddc80e781345e13b98a2dd58df4c4c1521727001b24dda47b4c9507bc629f4897deee05aa9ef4e842ddb758b9b0fb099ef41d3b9aaa061d6b7392cf3f62c45;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d4c1bf9436f49009004702bcf0b2b3272a02861932c1438a4cee8eaebc93cc214da11c9c864bb243c6a3e6c9006b4a2762154221d1a9526385b910ff26fcdb73c2d8646ed73512ac1c98d43c851ba4505dcff6dbb8bba5f996d3ee55681bcfee6be;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h3336c15afd730a722ae35f0236b7f1114389564bb6e056c585c2aa8f498865458eb24de57024f67642319031fa236fb6205e274c0912d5e08d5ebe7fe572c135e1b3d5a3794ca7c25c00a47b8b6f9ea700a5e7733b274a3bf7ea22f5f228dc44a8b1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1ab69b3d4bab6e795e61e219f6f6ea26cb5ad6db0f4dbb8e914620cfee2c4b7b5cedebced21ddce747d64fcdec6dd13eac3e9ceff5b54c3470d3adb4f9f58def43e93dd6b6300d830309fd2dea658c0291fd582c72912c9ae5fe2cb541b44c2271e3;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha195d9715b8a5ee3836045009fe4091b4699be926f0e27f7990a3527a846eab684b4642db3d2e20f81068433258e93a7efc18eeae93a9db54843b81986587aa20e322e29805e60c850519b5bb547626404bd33896d7d5b04b64cde2878344ace7093;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7778c9be5781cd73e18baf9f61ca62a14768a8e873b4731482f98f0697f4c509826e90379d788c8808837b8b2e64fa0e3f4e864a6cef14800dce1b6198527de50e5ec3c407568f70035a3c0a9ab56c41cdea4b2ab65db38a573683b2c13828a1af0c;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'haf29dbea94e72fb02afe400074aeced601e43ad8fc9420ec0b0b96f99f167e926e68b6f3c0aa1dca160d9e4c01d5f23e708ed215461ada66deb2347f19b3d6d51b551eddc8e03ad679d420cbddbec5c65cd8e633434daa3dfcb9f7086d749ea0a155;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hfa12c4365772821e74d8aeff1e13c6429217fdeda515fa7689e27d024eaf9953a7f167d0fccbfb2170d0b2698997d12c3e3609ff72e63a07034680b9b0d9b726ac88d1d970b11d669b2c07378cbef60c5186baec76665d33b96d8df33366ffb29eae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha661a53fddbce121bdc29fbeecde2d2648405d5ca985c094cead2b8cb3be8dd1cbbbec6cdeadd1250d8616228b3b939e2a8b44f2279351ee18497c9d1cc7d0c3a5532a9a630f0afe83cf1e51b2f5706e4b0446d4510051323ff9418eae8f35883029;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he80f64b01480c9e05ee8ce2a9e8db91e585b7abc4dc2bc7f9b9ad2107a88be28db9f1ad2c9eae4bcdfcebf138c9755e3a73774d9fa1c077ce06cd816b1b470e843dd76c6db38008f3fd0961cd386096371bb521e7f3c50f03ef6e650c22de050aed1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h7099b002a17a6560fd23f1ba95f93a3b5ce6140f2113c7377c0cd3048a2a21b98891a1b54001c570fceaac0c4910c8ae0e218fd7bf34c4b4f957beb6ee51e60e07b90819013d686c4558422c6a81a4d3a2d6603723d81cb1c907c31669b387e1bdb2;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hd5bc7b475e23f5362869ad53bd7cac86ef555b5f4dc193009ee2db5c114ee5e78ff112f4af03b058bb9ebb9c517754ee4205c0dc999d518258dc964fc161b51cc1b58a1aa9f0bed40bedd9e8ab620feed8af15599a0329f34200fa8ac7c1a55cbb14;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h4d12cacc55a2afad9253d383bc0327137bbee190b2ca0c0e658851b2dacd4200f8072ab236b6abf3a371357ebf61749389ca0a70ad506d04eab1b12de53d6701524b4ccc5cb82a2dfc74e08ea1bf26665d08d28e12fbaac60d54ff8ad98823441f;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h511ef98523549e8753ef4e749bb1943ffd5b4f0d6ebd8ebdd73f870de389e763cb06e71bc74f41a123d4722ffbcaa7effb80a0a4bed2691cd9ed4807bc3b491bf2cc11f898447ccc24d366e7c764a75a77f3a44c9cf43f4905d9e751cbffd7f29aae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hcd11ec2fd0e3b8097bb1a0cff7ce87cd4815e69a70620ff2c8c64f6f30fb95f7227b3ce91b1945e402b510c090456e23d4c44002f544431e7dc263d506c015ca4d9633390f38cbf0599d24d080103f659bbbf7beebd7f7c937c11764806ec3776e3a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6af42a2ef4047f64119997ca5a60d75dae842e536ab5a56b0368912f69a2035305d25c9f6c07d63210b966c1cb2c54d192e312c5109fd56148352d9c21229df5ca3e4e22ea92d4341beb9a6149bb20de55508199c3908b2fb8e559e01f0de453f865;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h6902668cedea0f940eacb9f3ab8db8da38a61cf4b982d98d29e22ca139696f78060ca9bf9e527d98ca2294b1ffbdd4705113d7877b6ed94e482011f2123486c2b36098a12db42435d4509a155208c864a7c31c183bf799af0442a2f8b9c78ba48a86;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h27f8dc14537077080d4b2e1ef6d7d4348cc488a4037fa8f28e2fd29d8668df7cfde32c906fc025e35d563cdd129d33e0e2fc8ef815cc33f1ad1caa39f51f99db6338ae0714ae803e549bcc860c8532635a4dd7d917acc3818bc1e11fed0344d567ae;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h96bb8359368fd329c8002949368498f04711e9b3a5ceaf877da728fccb5f70f9df0505eabdcc66cb7972ac4107bb15e318c567aad91cb576d5dfe8604866746a6ced7d483e5b5624ca41e0b1da202aff2b884e42590e21e1d040ac95015090f65441;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf4a3f05c99feef104b34b9824e3fca7f9464e172a9543ab6ab296003027bff03c29aaa928eed4c6cf11fdc0c401bf2dfbe649727a7d8f49d55af99589e634f37b60cccf0a8e0bf32c2d29fc43b1d6ff7917db08f619d86d859fdaf92b9a10e89977b;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'ha0ebec69df614ba2f01cb75a4fad988b7197af01f74abfc0b269fba9aed364b94ebc295e3cb25eff23ee924ad83cc95e1503921f45fc78e0ef260ccf08f78255d92186ea1c6fc01077c1055cec0a9bbc2d00946bc36593aea544c451910bdb3799aa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he97ebedd1676f6fb4ac79a0d52005cbdb8f191f9119e567b3793c1174c8da06f8bd37cafe96f16c95e174cbf834877ecb08acb48084a74e476a586a4d91efbe4350b7be101bebee8a8874c07158d9e377fec8122319d3038597c4621526cbb6741ff;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9da9c713fe1b03507fa8286df5b22411d66bff41a11a74aa2ff5452c77a7d08fbc00fa49703b221e7cf6513327a1a062027b0bed5a5fad3d78052fa044c67c3060100f42ef9a3e00225cad65eeaa3d0ecbc5eb5785ca356f27dc3d9836fec944dd5a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h2f3014c21e7d8e93be80b571b50399f867ca1323ac1c5b9063319385053d474c656a2e47341a579fd9005f552d2508e1cdf675b0a7f57c7b5382747acd54bf31b8bd6db83d7f8c601e917212f976a1f04c6edbc8b190ec8da5a5359e232340703e99;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h38352235570816629ababa24e36968dba1908bed1c0bcf8c4f53a1e97ba446f7552dac593a4c716e90853a3bf1af01977e9d12e720a2f43d18b76a354aed959636f671a2fa7951d385bf795014c4cd78866684f781bfbe5db82b577f57506ae22937;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'he2687dc9d058518eb62555427a7c7edd6d4492e9343f5f40af80b933ff119f1b50be88de14e58bc68d94fd92bb3165c9b16a7a949b3581c6daab5a3e095d1b89fd3552e24ce821b8c592af86ce26251e90f9a8389567797fd5f22abf8a0fa79fccd1;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc1b46ddfe5f433fd6d961bab42714c54ef92b787145e2955148ecbeaa1302c548f586524f45da00ab2dfc4946b037f91b902bf29d1f36b893726dff2bf57a163cc872133099aceb325a6a799e6263b417c1515eef9ad523324fe60baa148c9aa6b55;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hf937cff37b92af2bf2199d6e57eccb011adf1b8f1e03972179122668cbb107dcd109e033e30e4829395876a1de50b715200a154cbd5e577218cf1a564df4ecb872cff869f0247f30caab3724bbe865f347b68f92de110fa7ece94c6bb6fcd08ac187;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h779bda8428e62fbc76260808a8cf7cab4bc30bf535c4babea22f7d9abbbd34ba4c42a268c4d4d5b1373de9b522e236115dba3775c92bd8952e10ef4657592c1e5a8ae1e9f09b91ca017b7f45eeca1f0dc95fc112c8a633095d89fb68d070386d9d61;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h1d2438a8fb5ac96603377ed95b4f9e0e1d585e0a8e8f33005d0e5d561cd72c9b099e2834f147cce37145e113bedbc08215b4682b6638e8f33322e2e5060385e8a45665f8a24c64a5fbc1d18f7d2b4442f194a7606692765799fd70887d87362f819a;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hc011bb56e8ff18e5301e9f6bee276808f8a3e6fd74c5511e50cc969ddda8e87b6fcd317c800325e5ebf22859db24f155b848b3209681f7806a1b9a279a8a156541a8175c357d97d86d5aac017f169d929bea3c1b2f29b959a4056e1524368672c972;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'hb8cf0200b34cafc1c2bdea728278f8d14ed2ed3288d35374cfe1654d3de0d8fb76542697137ac0e6b393b0ebb48f44278c4af5615fb095c818407cf79514535a0a4c97cd779fe1b15655a68cd2e9e32ffd328b5014ecf5b3523fd6899a104fdb37ee;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h719c48b71b0f1d55fa756e22cac070e97fac6157f700a2ddffeb8b91ec7f6c6ce15f2534d38ef05c3b7e27d19d764fb8d83a472746f034ff1c6634e28ff5f4c75bfb8349bbdb1b9dd7b24b4df73d721b9f864742e3c9308d7432a926bb93569a3afa;
        #1
        {src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 784'h9a87d6f8362dbdfffff2806d523d589b802c8cba45d823b6877292c4a111dced84783f7197e8530c34d0e1008c2eb4216b49a6fc3cc2bb097f1c89219616249bfc98d5052ab9705353eba1cd3450f6d4d4e3cbdd70f6702a79a3e96ec591917f75f;
        #1
        $finish();
    end
endmodule
