module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    compressor_CLA256_12 compressor_CLA256_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA256_12(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [0:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], 1'h0, comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], 1'h0, comp_out0[1]}),
        .dst({dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [0:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [47:0] stage1_0;
   wire [89:0] stage1_1;
   wire [84:0] stage1_2;
   wire [96:0] stage1_3;
   wire [126:0] stage1_4;
   wire [128:0] stage1_5;
   wire [88:0] stage1_6;
   wire [90:0] stage1_7;
   wire [154:0] stage1_8;
   wire [119:0] stage1_9;
   wire [121:0] stage1_10;
   wire [82:0] stage1_11;
   wire [71:0] stage1_12;
   wire [41:0] stage1_13;
   wire [18:0] stage2_0;
   wire [24:0] stage2_1;
   wire [25:0] stage2_2;
   wire [41:0] stage2_3;
   wire [49:0] stage2_4;
   wire [41:0] stage2_5;
   wire [53:0] stage2_6;
   wire [47:0] stage2_7;
   wire [70:0] stage2_8;
   wire [42:0] stage2_9;
   wire [49:0] stage2_10;
   wire [46:0] stage2_11;
   wire [35:0] stage2_12;
   wire [35:0] stage2_13;
   wire [15:0] stage2_14;
   wire [4:0] stage2_15;
   wire [18:0] stage3_0;
   wire [4:0] stage3_1;
   wire [12:0] stage3_2;
   wire [10:0] stage3_3;
   wire [18:0] stage3_4;
   wire [17:0] stage3_5;
   wire [22:0] stage3_6;
   wire [20:0] stage3_7;
   wire [23:0] stage3_8;
   wire [27:0] stage3_9;
   wire [19:0] stage3_10;
   wire [21:0] stage3_11;
   wire [18:0] stage3_12;
   wire [12:0] stage3_13;
   wire [11:0] stage3_14;
   wire [12:0] stage3_15;
   wire [2:0] stage3_16;
   wire [13:0] stage4_0;
   wire [5:0] stage4_1;
   wire [3:0] stage4_2;
   wire [3:0] stage4_3;
   wire [6:0] stage4_4;
   wire [6:0] stage4_5;
   wire [12:0] stage4_6;
   wire [6:0] stage4_7;
   wire [11:0] stage4_8;
   wire [10:0] stage4_9;
   wire [8:0] stage4_10;
   wire [11:0] stage4_11;
   wire [8:0] stage4_12;
   wire [8:0] stage4_13;
   wire [4:0] stage4_14;
   wire [11:0] stage4_15;
   wire [3:0] stage4_16;
   wire [1:0] stage4_17;
   wire [5:0] stage5_0;
   wire [1:0] stage5_1;
   wire [3:0] stage5_2;
   wire [1:0] stage5_3;
   wire [4:0] stage5_4;
   wire [1:0] stage5_5;
   wire [4:0] stage5_6;
   wire [2:0] stage5_7;
   wire [3:0] stage5_8;
   wire [5:0] stage5_9;
   wire [4:0] stage5_10;
   wire [2:0] stage5_11;
   wire [3:0] stage5_12;
   wire [5:0] stage5_13;
   wire [5:0] stage5_14;
   wire [1:0] stage5_15;
   wire [5:0] stage5_16;
   wire [3:0] stage5_17;
   wire [1:0] stage6_0;
   wire [0:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [0:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [0:0] stage6_19;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[2]},
      {stage0_3[4]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[13], stage0_0[14], stage0_0[15]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[3]},
      {stage0_3[5]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[16], stage0_0[17], stage0_0[18]},
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[4]},
      {stage0_3[6]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[19], stage0_0[20], stage0_0[21]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[5]},
      {stage0_3[7]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[6]},
      {stage0_3[8]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[145], stage0_0[146], stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[151], stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[163], stage0_0[164], stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[169], stage0_0[170], stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[175], stage0_0[176], stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180]},
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[181], stage0_0[182], stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186]},
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[187], stage0_0[188], stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192]},
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198]},
      {stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204]},
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210]},
      {stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216]},
      {stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222]},
      {stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228]},
      {stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234]},
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240]},
      {stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246]},
      {stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252]},
      {stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[0],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[1],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[2],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[3],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[4],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[5],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[6],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[7],stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[8],stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[9],stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[10],stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[11],stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[12],stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[13],stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[14],stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[15],stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[16],stage1_4[61],stage1_3[61],stage1_2[61],stage1_1[61]}
   );
   gpc606_5 gpc62 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage1_5[17],stage1_4[62],stage1_3[62],stage1_2[62],stage1_1[62]}
   );
   gpc606_5 gpc63 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122]},
      {stage1_5[18],stage1_4[63],stage1_3[63],stage1_2[63],stage1_1[63]}
   );
   gpc606_5 gpc64 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage1_5[19],stage1_4[64],stage1_3[64],stage1_2[64],stage1_1[64]}
   );
   gpc606_5 gpc65 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage1_5[20],stage1_4[65],stage1_3[65],stage1_2[65],stage1_1[65]}
   );
   gpc606_5 gpc66 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140]},
      {stage1_5[21],stage1_4[66],stage1_3[66],stage1_2[66],stage1_1[66]}
   );
   gpc606_5 gpc67 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146]},
      {stage1_5[22],stage1_4[67],stage1_3[67],stage1_2[67],stage1_1[67]}
   );
   gpc606_5 gpc68 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152]},
      {stage1_5[23],stage1_4[68],stage1_3[68],stage1_2[68],stage1_1[68]}
   );
   gpc606_5 gpc69 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage1_5[24],stage1_4[69],stage1_3[69],stage1_2[69],stage1_1[69]}
   );
   gpc606_5 gpc70 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage1_5[25],stage1_4[70],stage1_3[70],stage1_2[70],stage1_1[70]}
   );
   gpc606_5 gpc71 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170]},
      {stage1_5[26],stage1_4[71],stage1_3[71],stage1_2[71],stage1_1[71]}
   );
   gpc606_5 gpc72 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage1_5[27],stage1_4[72],stage1_3[72],stage1_2[72],stage1_1[72]}
   );
   gpc606_5 gpc73 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182]},
      {stage1_5[28],stage1_4[73],stage1_3[73],stage1_2[73],stage1_1[73]}
   );
   gpc606_5 gpc74 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage1_5[29],stage1_4[74],stage1_3[74],stage1_2[74],stage1_1[74]}
   );
   gpc606_5 gpc75 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage1_5[30],stage1_4[75],stage1_3[75],stage1_2[75],stage1_1[75]}
   );
   gpc606_5 gpc76 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200]},
      {stage1_5[31],stage1_4[76],stage1_3[76],stage1_2[76],stage1_1[76]}
   );
   gpc606_5 gpc77 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage1_5[32],stage1_4[77],stage1_3[77],stage1_2[77],stage1_1[77]}
   );
   gpc606_5 gpc78 (
      {stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239]},
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212]},
      {stage1_5[33],stage1_4[78],stage1_3[78],stage1_2[78],stage1_1[78]}
   );
   gpc606_5 gpc79 (
      {stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245]},
      {stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218]},
      {stage1_5[34],stage1_4[79],stage1_3[79],stage1_2[79],stage1_1[79]}
   );
   gpc615_5 gpc80 (
      {stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239]},
      {stage0_3[219]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[35],stage1_4[80],stage1_3[80],stage1_2[80]}
   );
   gpc615_5 gpc81 (
      {stage0_2[240], stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244]},
      {stage0_3[220]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[36],stage1_4[81],stage1_3[81],stage1_2[81]}
   );
   gpc615_5 gpc82 (
      {stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248], stage0_2[249]},
      {stage0_3[221]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[37],stage1_4[82],stage1_3[82],stage1_2[82]}
   );
   gpc615_5 gpc83 (
      {stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage0_3[222]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[38],stage1_4[83],stage1_3[83],stage1_2[83]}
   );
   gpc615_5 gpc84 (
      {stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226], stage0_3[227]},
      {stage0_4[24]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[39],stage1_4[84],stage1_3[84]}
   );
   gpc615_5 gpc85 (
      {stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232]},
      {stage0_4[25]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[5],stage1_5[40],stage1_4[85],stage1_3[85]}
   );
   gpc615_5 gpc86 (
      {stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237]},
      {stage0_4[26]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[6],stage1_5[41],stage1_4[86],stage1_3[86]}
   );
   gpc615_5 gpc87 (
      {stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242]},
      {stage0_4[27]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[7],stage1_5[42],stage1_4[87],stage1_3[87]}
   );
   gpc615_5 gpc88 (
      {stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246], stage0_3[247]},
      {stage0_4[28]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[8],stage1_5[43],stage1_4[88],stage1_3[88]}
   );
   gpc606_5 gpc89 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[5],stage1_6[9],stage1_5[44],stage1_4[89]}
   );
   gpc606_5 gpc90 (
      {stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[6],stage1_6[10],stage1_5[45],stage1_4[90]}
   );
   gpc606_5 gpc91 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[7],stage1_6[11],stage1_5[46],stage1_4[91]}
   );
   gpc606_5 gpc92 (
      {stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[8],stage1_6[12],stage1_5[47],stage1_4[92]}
   );
   gpc606_5 gpc93 (
      {stage0_4[53], stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[9],stage1_6[13],stage1_5[48],stage1_4[93]}
   );
   gpc606_5 gpc94 (
      {stage0_4[59], stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[10],stage1_6[14],stage1_5[49],stage1_4[94]}
   );
   gpc606_5 gpc95 (
      {stage0_4[65], stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[11],stage1_6[15],stage1_5[50],stage1_4[95]}
   );
   gpc606_5 gpc96 (
      {stage0_4[71], stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[12],stage1_6[16],stage1_5[51],stage1_4[96]}
   );
   gpc606_5 gpc97 (
      {stage0_4[77], stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[13],stage1_6[17],stage1_5[52],stage1_4[97]}
   );
   gpc606_5 gpc98 (
      {stage0_4[83], stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[14],stage1_6[18],stage1_5[53],stage1_4[98]}
   );
   gpc606_5 gpc99 (
      {stage0_4[89], stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[15],stage1_6[19],stage1_5[54],stage1_4[99]}
   );
   gpc606_5 gpc100 (
      {stage0_4[95], stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[16],stage1_6[20],stage1_5[55],stage1_4[100]}
   );
   gpc606_5 gpc101 (
      {stage0_4[101], stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[17],stage1_6[21],stage1_5[56],stage1_4[101]}
   );
   gpc606_5 gpc102 (
      {stage0_4[107], stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[18],stage1_6[22],stage1_5[57],stage1_4[102]}
   );
   gpc606_5 gpc103 (
      {stage0_4[113], stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[19],stage1_6[23],stage1_5[58],stage1_4[103]}
   );
   gpc606_5 gpc104 (
      {stage0_4[119], stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[20],stage1_6[24],stage1_5[59],stage1_4[104]}
   );
   gpc606_5 gpc105 (
      {stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[21],stage1_6[25],stage1_5[60],stage1_4[105]}
   );
   gpc606_5 gpc106 (
      {stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[22],stage1_6[26],stage1_5[61],stage1_4[106]}
   );
   gpc606_5 gpc107 (
      {stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[23],stage1_6[27],stage1_5[62],stage1_4[107]}
   );
   gpc606_5 gpc108 (
      {stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[24],stage1_6[28],stage1_5[63],stage1_4[108]}
   );
   gpc606_5 gpc109 (
      {stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[25],stage1_6[29],stage1_5[64],stage1_4[109]}
   );
   gpc606_5 gpc110 (
      {stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[26],stage1_6[30],stage1_5[65],stage1_4[110]}
   );
   gpc606_5 gpc111 (
      {stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[27],stage1_6[31],stage1_5[66],stage1_4[111]}
   );
   gpc606_5 gpc112 (
      {stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[28],stage1_6[32],stage1_5[67],stage1_4[112]}
   );
   gpc606_5 gpc113 (
      {stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[29],stage1_6[33],stage1_5[68],stage1_4[113]}
   );
   gpc606_5 gpc114 (
      {stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[30],stage1_6[34],stage1_5[69],stage1_4[114]}
   );
   gpc606_5 gpc115 (
      {stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189], stage0_4[190]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[31],stage1_6[35],stage1_5[70],stage1_4[115]}
   );
   gpc606_5 gpc116 (
      {stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195], stage0_4[196]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[32],stage1_6[36],stage1_5[71],stage1_4[116]}
   );
   gpc606_5 gpc117 (
      {stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[33],stage1_6[37],stage1_5[72],stage1_4[117]}
   );
   gpc606_5 gpc118 (
      {stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[34],stage1_6[38],stage1_5[73],stage1_4[118]}
   );
   gpc606_5 gpc119 (
      {stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[35],stage1_6[39],stage1_5[74],stage1_4[119]}
   );
   gpc606_5 gpc120 (
      {stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[36],stage1_6[40],stage1_5[75],stage1_4[120]}
   );
   gpc606_5 gpc121 (
      {stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[37],stage1_6[41],stage1_5[76],stage1_4[121]}
   );
   gpc606_5 gpc122 (
      {stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[38],stage1_6[42],stage1_5[77],stage1_4[122]}
   );
   gpc606_5 gpc123 (
      {stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[39],stage1_6[43],stage1_5[78],stage1_4[123]}
   );
   gpc606_5 gpc124 (
      {stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[40],stage1_6[44],stage1_5[79],stage1_4[124]}
   );
   gpc606_5 gpc125 (
      {stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[41],stage1_6[45],stage1_5[80],stage1_4[125]}
   );
   gpc615_5 gpc126 (
      {stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255]},
      {stage0_5[30]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[42],stage1_6[46],stage1_5[81],stage1_4[126]}
   );
   gpc606_5 gpc127 (
      {stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[38],stage1_7[43],stage1_6[47],stage1_5[82]}
   );
   gpc606_5 gpc128 (
      {stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[39],stage1_7[44],stage1_6[48],stage1_5[83]}
   );
   gpc606_5 gpc129 (
      {stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[40],stage1_7[45],stage1_6[49],stage1_5[84]}
   );
   gpc606_5 gpc130 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[41],stage1_7[46],stage1_6[50],stage1_5[85]}
   );
   gpc606_5 gpc131 (
      {stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[42],stage1_7[47],stage1_6[51],stage1_5[86]}
   );
   gpc606_5 gpc132 (
      {stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[43],stage1_7[48],stage1_6[52],stage1_5[87]}
   );
   gpc606_5 gpc133 (
      {stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[44],stage1_7[49],stage1_6[53],stage1_5[88]}
   );
   gpc606_5 gpc134 (
      {stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[45],stage1_7[50],stage1_6[54],stage1_5[89]}
   );
   gpc606_5 gpc135 (
      {stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[46],stage1_7[51],stage1_6[55],stage1_5[90]}
   );
   gpc606_5 gpc136 (
      {stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[47],stage1_7[52],stage1_6[56],stage1_5[91]}
   );
   gpc606_5 gpc137 (
      {stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[48],stage1_7[53],stage1_6[57],stage1_5[92]}
   );
   gpc606_5 gpc138 (
      {stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[49],stage1_7[54],stage1_6[58],stage1_5[93]}
   );
   gpc606_5 gpc139 (
      {stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[50],stage1_7[55],stage1_6[59],stage1_5[94]}
   );
   gpc606_5 gpc140 (
      {stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[51],stage1_7[56],stage1_6[60],stage1_5[95]}
   );
   gpc606_5 gpc141 (
      {stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[52],stage1_7[57],stage1_6[61],stage1_5[96]}
   );
   gpc606_5 gpc142 (
      {stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[53],stage1_7[58],stage1_6[62],stage1_5[97]}
   );
   gpc606_5 gpc143 (
      {stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131], stage0_5[132]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[54],stage1_7[59],stage1_6[63],stage1_5[98]}
   );
   gpc606_5 gpc144 (
      {stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137], stage0_5[138]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[55],stage1_7[60],stage1_6[64],stage1_5[99]}
   );
   gpc606_5 gpc145 (
      {stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[56],stage1_7[61],stage1_6[65],stage1_5[100]}
   );
   gpc606_5 gpc146 (
      {stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[57],stage1_7[62],stage1_6[66],stage1_5[101]}
   );
   gpc606_5 gpc147 (
      {stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[58],stage1_7[63],stage1_6[67],stage1_5[102]}
   );
   gpc606_5 gpc148 (
      {stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[59],stage1_7[64],stage1_6[68],stage1_5[103]}
   );
   gpc606_5 gpc149 (
      {stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[60],stage1_7[65],stage1_6[69],stage1_5[104]}
   );
   gpc606_5 gpc150 (
      {stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[61],stage1_7[66],stage1_6[70],stage1_5[105]}
   );
   gpc606_5 gpc151 (
      {stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[62],stage1_7[67],stage1_6[71],stage1_5[106]}
   );
   gpc606_5 gpc152 (
      {stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[63],stage1_7[68],stage1_6[72],stage1_5[107]}
   );
   gpc606_5 gpc153 (
      {stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[64],stage1_7[69],stage1_6[73],stage1_5[108]}
   );
   gpc606_5 gpc154 (
      {stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[65],stage1_7[70],stage1_6[74],stage1_5[109]}
   );
   gpc606_5 gpc155 (
      {stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[66],stage1_7[71],stage1_6[75],stage1_5[110]}
   );
   gpc606_5 gpc156 (
      {stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[67],stage1_7[72],stage1_6[76],stage1_5[111]}
   );
   gpc606_5 gpc157 (
      {stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[68],stage1_7[73],stage1_6[77],stage1_5[112]}
   );
   gpc606_5 gpc158 (
      {stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[69],stage1_7[74],stage1_6[78],stage1_5[113]}
   );
   gpc606_5 gpc159 (
      {stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[70],stage1_7[75],stage1_6[79],stage1_5[114]}
   );
   gpc606_5 gpc160 (
      {stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[71],stage1_7[76],stage1_6[80],stage1_5[115]}
   );
   gpc615_5 gpc161 (
      {stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_6[228]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[72],stage1_7[77],stage1_6[81],stage1_5[116]}
   );
   gpc615_5 gpc162 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244]},
      {stage0_6[229]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[73],stage1_7[78],stage1_6[82],stage1_5[117]}
   );
   gpc615_5 gpc163 (
      {stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233], stage0_6[234]},
      {stage0_7[216]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[36],stage1_8[74],stage1_7[79],stage1_6[83]}
   );
   gpc615_5 gpc164 (
      {stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage0_7[217]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[37],stage1_8[75],stage1_7[80],stage1_6[84]}
   );
   gpc615_5 gpc165 (
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244]},
      {stage0_7[218]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[38],stage1_8[76],stage1_7[81],stage1_6[85]}
   );
   gpc615_5 gpc166 (
      {stage0_6[245], stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249]},
      {stage0_7[219]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[39],stage1_8[77],stage1_7[82],stage1_6[86]}
   );
   gpc615_5 gpc167 (
      {stage0_6[250], stage0_6[251], stage0_6[252], stage0_6[253], stage0_6[254]},
      {stage0_7[220]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[40],stage1_8[78],stage1_7[83],stage1_6[87]}
   );
   gpc615_5 gpc168 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[30]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[5],stage1_9[41],stage1_8[79],stage1_7[84]}
   );
   gpc615_5 gpc169 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[31]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[6],stage1_9[42],stage1_8[80],stage1_7[85]}
   );
   gpc615_5 gpc170 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[32]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[7],stage1_9[43],stage1_8[81],stage1_7[86]}
   );
   gpc615_5 gpc171 (
      {stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239], stage0_7[240]},
      {stage0_8[33]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[8],stage1_9[44],stage1_8[82],stage1_7[87]}
   );
   gpc615_5 gpc172 (
      {stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage0_8[34]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[9],stage1_9[45],stage1_8[83],stage1_7[88]}
   );
   gpc615_5 gpc173 (
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250]},
      {stage0_8[35]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[10],stage1_9[46],stage1_8[84],stage1_7[89]}
   );
   gpc615_5 gpc174 (
      {stage0_7[251], stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255]},
      {stage0_8[36]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[11],stage1_9[47],stage1_8[85],stage1_7[90]}
   );
   gpc606_5 gpc175 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[7],stage1_10[12],stage1_9[48],stage1_8[86]}
   );
   gpc606_5 gpc176 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[8],stage1_10[13],stage1_9[49],stage1_8[87]}
   );
   gpc606_5 gpc177 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[9],stage1_10[14],stage1_9[50],stage1_8[88]}
   );
   gpc606_5 gpc178 (
      {stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[10],stage1_10[15],stage1_9[51],stage1_8[89]}
   );
   gpc606_5 gpc179 (
      {stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[11],stage1_10[16],stage1_9[52],stage1_8[90]}
   );
   gpc606_5 gpc180 (
      {stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[12],stage1_10[17],stage1_9[53],stage1_8[91]}
   );
   gpc606_5 gpc181 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[13],stage1_10[18],stage1_9[54],stage1_8[92]}
   );
   gpc606_5 gpc182 (
      {stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[14],stage1_10[19],stage1_9[55],stage1_8[93]}
   );
   gpc606_5 gpc183 (
      {stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[15],stage1_10[20],stage1_9[56],stage1_8[94]}
   );
   gpc606_5 gpc184 (
      {stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[16],stage1_10[21],stage1_9[57],stage1_8[95]}
   );
   gpc606_5 gpc185 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[17],stage1_10[22],stage1_9[58],stage1_8[96]}
   );
   gpc606_5 gpc186 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[18],stage1_10[23],stage1_9[59],stage1_8[97]}
   );
   gpc606_5 gpc187 (
      {stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[19],stage1_10[24],stage1_9[60],stage1_8[98]}
   );
   gpc606_5 gpc188 (
      {stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[20],stage1_10[25],stage1_9[61],stage1_8[99]}
   );
   gpc606_5 gpc189 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[21],stage1_10[26],stage1_9[62],stage1_8[100]}
   );
   gpc606_5 gpc190 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[22],stage1_10[27],stage1_9[63],stage1_8[101]}
   );
   gpc606_5 gpc191 (
      {stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[23],stage1_10[28],stage1_9[64],stage1_8[102]}
   );
   gpc606_5 gpc192 (
      {stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[24],stage1_10[29],stage1_9[65],stage1_8[103]}
   );
   gpc606_5 gpc193 (
      {stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[25],stage1_10[30],stage1_9[66],stage1_8[104]}
   );
   gpc606_5 gpc194 (
      {stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[26],stage1_10[31],stage1_9[67],stage1_8[105]}
   );
   gpc606_5 gpc195 (
      {stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[27],stage1_10[32],stage1_9[68],stage1_8[106]}
   );
   gpc606_5 gpc196 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[28],stage1_10[33],stage1_9[69],stage1_8[107]}
   );
   gpc606_5 gpc197 (
      {stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[29],stage1_10[34],stage1_9[70],stage1_8[108]}
   );
   gpc606_5 gpc198 (
      {stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[30],stage1_10[35],stage1_9[71],stage1_8[109]}
   );
   gpc606_5 gpc199 (
      {stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[31],stage1_10[36],stage1_9[72],stage1_8[110]}
   );
   gpc606_5 gpc200 (
      {stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[32],stage1_10[37],stage1_9[73],stage1_8[111]}
   );
   gpc606_5 gpc201 (
      {stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[33],stage1_10[38],stage1_9[74],stage1_8[112]}
   );
   gpc606_5 gpc202 (
      {stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[34],stage1_10[39],stage1_9[75],stage1_8[113]}
   );
   gpc606_5 gpc203 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[35],stage1_10[40],stage1_9[76],stage1_8[114]}
   );
   gpc606_5 gpc204 (
      {stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[36],stage1_10[41],stage1_9[77],stage1_8[115]}
   );
   gpc606_5 gpc205 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[30],stage1_11[37],stage1_10[42],stage1_9[78]}
   );
   gpc606_5 gpc206 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[31],stage1_11[38],stage1_10[43],stage1_9[79]}
   );
   gpc606_5 gpc207 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[32],stage1_11[39],stage1_10[44],stage1_9[80]}
   );
   gpc606_5 gpc208 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[33],stage1_11[40],stage1_10[45],stage1_9[81]}
   );
   gpc615_5 gpc209 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70]},
      {stage0_10[180]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[34],stage1_11[41],stage1_10[46],stage1_9[82]}
   );
   gpc615_5 gpc210 (
      {stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75]},
      {stage0_10[181]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[35],stage1_11[42],stage1_10[47],stage1_9[83]}
   );
   gpc615_5 gpc211 (
      {stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80]},
      {stage0_10[182]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[36],stage1_11[43],stage1_10[48],stage1_9[84]}
   );
   gpc615_5 gpc212 (
      {stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85]},
      {stage0_10[183]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[37],stage1_11[44],stage1_10[49],stage1_9[85]}
   );
   gpc615_5 gpc213 (
      {stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90]},
      {stage0_10[184]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[38],stage1_11[45],stage1_10[50],stage1_9[86]}
   );
   gpc615_5 gpc214 (
      {stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_10[185]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[39],stage1_11[46],stage1_10[51],stage1_9[87]}
   );
   gpc615_5 gpc215 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100]},
      {stage0_10[186]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[40],stage1_11[47],stage1_10[52],stage1_9[88]}
   );
   gpc615_5 gpc216 (
      {stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105]},
      {stage0_10[187]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[41],stage1_11[48],stage1_10[53],stage1_9[89]}
   );
   gpc615_5 gpc217 (
      {stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110]},
      {stage0_10[188]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[42],stage1_11[49],stage1_10[54],stage1_9[90]}
   );
   gpc615_5 gpc218 (
      {stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115]},
      {stage0_10[189]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[43],stage1_11[50],stage1_10[55],stage1_9[91]}
   );
   gpc615_5 gpc219 (
      {stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120]},
      {stage0_10[190]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[44],stage1_11[51],stage1_10[56],stage1_9[92]}
   );
   gpc615_5 gpc220 (
      {stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_10[191]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[45],stage1_11[52],stage1_10[57],stage1_9[93]}
   );
   gpc615_5 gpc221 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130]},
      {stage0_10[192]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[46],stage1_11[53],stage1_10[58],stage1_9[94]}
   );
   gpc615_5 gpc222 (
      {stage0_9[131], stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135]},
      {stage0_10[193]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[47],stage1_11[54],stage1_10[59],stage1_9[95]}
   );
   gpc615_5 gpc223 (
      {stage0_9[136], stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140]},
      {stage0_10[194]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[48],stage1_11[55],stage1_10[60],stage1_9[96]}
   );
   gpc615_5 gpc224 (
      {stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145]},
      {stage0_10[195]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[49],stage1_11[56],stage1_10[61],stage1_9[97]}
   );
   gpc615_5 gpc225 (
      {stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150]},
      {stage0_10[196]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[50],stage1_11[57],stage1_10[62],stage1_9[98]}
   );
   gpc615_5 gpc226 (
      {stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_10[197]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[51],stage1_11[58],stage1_10[63],stage1_9[99]}
   );
   gpc615_5 gpc227 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_10[198]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[52],stage1_11[59],stage1_10[64],stage1_9[100]}
   );
   gpc615_5 gpc228 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165]},
      {stage0_10[199]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[53],stage1_11[60],stage1_10[65],stage1_9[101]}
   );
   gpc615_5 gpc229 (
      {stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_10[200]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[54],stage1_11[61],stage1_10[66],stage1_9[102]}
   );
   gpc615_5 gpc230 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175]},
      {stage0_10[201]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[55],stage1_11[62],stage1_10[67],stage1_9[103]}
   );
   gpc615_5 gpc231 (
      {stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_10[202]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[56],stage1_11[63],stage1_10[68],stage1_9[104]}
   );
   gpc615_5 gpc232 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_10[203]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[57],stage1_11[64],stage1_10[69],stage1_9[105]}
   );
   gpc615_5 gpc233 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190]},
      {stage0_10[204]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[58],stage1_11[65],stage1_10[70],stage1_9[106]}
   );
   gpc615_5 gpc234 (
      {stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_10[205]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[59],stage1_11[66],stage1_10[71],stage1_9[107]}
   );
   gpc615_5 gpc235 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_10[206]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[60],stage1_11[67],stage1_10[72],stage1_9[108]}
   );
   gpc615_5 gpc236 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205]},
      {stage0_10[207]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[61],stage1_11[68],stage1_10[73],stage1_9[109]}
   );
   gpc615_5 gpc237 (
      {stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_10[208]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[62],stage1_11[69],stage1_10[74],stage1_9[110]}
   );
   gpc615_5 gpc238 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_10[209]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[63],stage1_11[70],stage1_10[75],stage1_9[111]}
   );
   gpc615_5 gpc239 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220]},
      {stage0_10[210]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[64],stage1_11[71],stage1_10[76],stage1_9[112]}
   );
   gpc615_5 gpc240 (
      {stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_10[211]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[65],stage1_11[72],stage1_10[77],stage1_9[113]}
   );
   gpc615_5 gpc241 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_10[212]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[66],stage1_11[73],stage1_10[78],stage1_9[114]}
   );
   gpc615_5 gpc242 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235]},
      {stage0_10[213]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[67],stage1_11[74],stage1_10[79],stage1_9[115]}
   );
   gpc615_5 gpc243 (
      {stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_10[214]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[68],stage1_11[75],stage1_10[80],stage1_9[116]}
   );
   gpc615_5 gpc244 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_10[215]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[69],stage1_11[76],stage1_10[81],stage1_9[117]}
   );
   gpc615_5 gpc245 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250]},
      {stage0_10[216]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[70],stage1_11[77],stage1_10[82],stage1_9[118]}
   );
   gpc615_5 gpc246 (
      {stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_10[217]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[71],stage1_11[78],stage1_10[83],stage1_9[119]}
   );
   gpc1_1 gpc247 (
      {stage0_0[253]},
      {stage1_0[45]}
   );
   gpc1_1 gpc248 (
      {stage0_0[254]},
      {stage1_0[46]}
   );
   gpc1_1 gpc249 (
      {stage0_0[255]},
      {stage1_0[47]}
   );
   gpc1_1 gpc250 (
      {stage0_1[246]},
      {stage1_1[80]}
   );
   gpc1_1 gpc251 (
      {stage0_1[247]},
      {stage1_1[81]}
   );
   gpc1_1 gpc252 (
      {stage0_1[248]},
      {stage1_1[82]}
   );
   gpc1_1 gpc253 (
      {stage0_1[249]},
      {stage1_1[83]}
   );
   gpc1_1 gpc254 (
      {stage0_1[250]},
      {stage1_1[84]}
   );
   gpc1_1 gpc255 (
      {stage0_1[251]},
      {stage1_1[85]}
   );
   gpc1_1 gpc256 (
      {stage0_1[252]},
      {stage1_1[86]}
   );
   gpc1_1 gpc257 (
      {stage0_1[253]},
      {stage1_1[87]}
   );
   gpc1_1 gpc258 (
      {stage0_1[254]},
      {stage1_1[88]}
   );
   gpc1_1 gpc259 (
      {stage0_1[255]},
      {stage1_1[89]}
   );
   gpc1_1 gpc260 (
      {stage0_2[255]},
      {stage1_2[84]}
   );
   gpc1_1 gpc261 (
      {stage0_3[248]},
      {stage1_3[89]}
   );
   gpc1_1 gpc262 (
      {stage0_3[249]},
      {stage1_3[90]}
   );
   gpc1_1 gpc263 (
      {stage0_3[250]},
      {stage1_3[91]}
   );
   gpc1_1 gpc264 (
      {stage0_3[251]},
      {stage1_3[92]}
   );
   gpc1_1 gpc265 (
      {stage0_3[252]},
      {stage1_3[93]}
   );
   gpc1_1 gpc266 (
      {stage0_3[253]},
      {stage1_3[94]}
   );
   gpc1_1 gpc267 (
      {stage0_3[254]},
      {stage1_3[95]}
   );
   gpc1_1 gpc268 (
      {stage0_3[255]},
      {stage1_3[96]}
   );
   gpc1_1 gpc269 (
      {stage0_5[245]},
      {stage1_5[118]}
   );
   gpc1_1 gpc270 (
      {stage0_5[246]},
      {stage1_5[119]}
   );
   gpc1_1 gpc271 (
      {stage0_5[247]},
      {stage1_5[120]}
   );
   gpc1_1 gpc272 (
      {stage0_5[248]},
      {stage1_5[121]}
   );
   gpc1_1 gpc273 (
      {stage0_5[249]},
      {stage1_5[122]}
   );
   gpc1_1 gpc274 (
      {stage0_5[250]},
      {stage1_5[123]}
   );
   gpc1_1 gpc275 (
      {stage0_5[251]},
      {stage1_5[124]}
   );
   gpc1_1 gpc276 (
      {stage0_5[252]},
      {stage1_5[125]}
   );
   gpc1_1 gpc277 (
      {stage0_5[253]},
      {stage1_5[126]}
   );
   gpc1_1 gpc278 (
      {stage0_5[254]},
      {stage1_5[127]}
   );
   gpc1_1 gpc279 (
      {stage0_5[255]},
      {stage1_5[128]}
   );
   gpc1_1 gpc280 (
      {stage0_6[255]},
      {stage1_6[88]}
   );
   gpc1_1 gpc281 (
      {stage0_8[217]},
      {stage1_8[116]}
   );
   gpc1_1 gpc282 (
      {stage0_8[218]},
      {stage1_8[117]}
   );
   gpc1_1 gpc283 (
      {stage0_8[219]},
      {stage1_8[118]}
   );
   gpc1_1 gpc284 (
      {stage0_8[220]},
      {stage1_8[119]}
   );
   gpc1_1 gpc285 (
      {stage0_8[221]},
      {stage1_8[120]}
   );
   gpc1_1 gpc286 (
      {stage0_8[222]},
      {stage1_8[121]}
   );
   gpc1_1 gpc287 (
      {stage0_8[223]},
      {stage1_8[122]}
   );
   gpc1_1 gpc288 (
      {stage0_8[224]},
      {stage1_8[123]}
   );
   gpc1_1 gpc289 (
      {stage0_8[225]},
      {stage1_8[124]}
   );
   gpc1_1 gpc290 (
      {stage0_8[226]},
      {stage1_8[125]}
   );
   gpc1_1 gpc291 (
      {stage0_8[227]},
      {stage1_8[126]}
   );
   gpc1_1 gpc292 (
      {stage0_8[228]},
      {stage1_8[127]}
   );
   gpc1_1 gpc293 (
      {stage0_8[229]},
      {stage1_8[128]}
   );
   gpc1_1 gpc294 (
      {stage0_8[230]},
      {stage1_8[129]}
   );
   gpc1_1 gpc295 (
      {stage0_8[231]},
      {stage1_8[130]}
   );
   gpc1_1 gpc296 (
      {stage0_8[232]},
      {stage1_8[131]}
   );
   gpc1_1 gpc297 (
      {stage0_8[233]},
      {stage1_8[132]}
   );
   gpc1_1 gpc298 (
      {stage0_8[234]},
      {stage1_8[133]}
   );
   gpc1_1 gpc299 (
      {stage0_8[235]},
      {stage1_8[134]}
   );
   gpc1_1 gpc300 (
      {stage0_8[236]},
      {stage1_8[135]}
   );
   gpc1_1 gpc301 (
      {stage0_8[237]},
      {stage1_8[136]}
   );
   gpc1_1 gpc302 (
      {stage0_8[238]},
      {stage1_8[137]}
   );
   gpc1_1 gpc303 (
      {stage0_8[239]},
      {stage1_8[138]}
   );
   gpc1_1 gpc304 (
      {stage0_8[240]},
      {stage1_8[139]}
   );
   gpc1_1 gpc305 (
      {stage0_8[241]},
      {stage1_8[140]}
   );
   gpc1_1 gpc306 (
      {stage0_8[242]},
      {stage1_8[141]}
   );
   gpc1_1 gpc307 (
      {stage0_8[243]},
      {stage1_8[142]}
   );
   gpc1_1 gpc308 (
      {stage0_8[244]},
      {stage1_8[143]}
   );
   gpc1_1 gpc309 (
      {stage0_8[245]},
      {stage1_8[144]}
   );
   gpc1_1 gpc310 (
      {stage0_8[246]},
      {stage1_8[145]}
   );
   gpc1_1 gpc311 (
      {stage0_8[247]},
      {stage1_8[146]}
   );
   gpc1_1 gpc312 (
      {stage0_8[248]},
      {stage1_8[147]}
   );
   gpc1_1 gpc313 (
      {stage0_8[249]},
      {stage1_8[148]}
   );
   gpc1_1 gpc314 (
      {stage0_8[250]},
      {stage1_8[149]}
   );
   gpc1_1 gpc315 (
      {stage0_8[251]},
      {stage1_8[150]}
   );
   gpc1_1 gpc316 (
      {stage0_8[252]},
      {stage1_8[151]}
   );
   gpc1_1 gpc317 (
      {stage0_8[253]},
      {stage1_8[152]}
   );
   gpc1_1 gpc318 (
      {stage0_8[254]},
      {stage1_8[153]}
   );
   gpc1_1 gpc319 (
      {stage0_8[255]},
      {stage1_8[154]}
   );
   gpc1_1 gpc320 (
      {stage0_10[218]},
      {stage1_10[84]}
   );
   gpc1_1 gpc321 (
      {stage0_10[219]},
      {stage1_10[85]}
   );
   gpc1_1 gpc322 (
      {stage0_10[220]},
      {stage1_10[86]}
   );
   gpc1_1 gpc323 (
      {stage0_10[221]},
      {stage1_10[87]}
   );
   gpc1_1 gpc324 (
      {stage0_10[222]},
      {stage1_10[88]}
   );
   gpc1_1 gpc325 (
      {stage0_10[223]},
      {stage1_10[89]}
   );
   gpc1_1 gpc326 (
      {stage0_10[224]},
      {stage1_10[90]}
   );
   gpc1_1 gpc327 (
      {stage0_10[225]},
      {stage1_10[91]}
   );
   gpc1_1 gpc328 (
      {stage0_10[226]},
      {stage1_10[92]}
   );
   gpc1_1 gpc329 (
      {stage0_10[227]},
      {stage1_10[93]}
   );
   gpc1_1 gpc330 (
      {stage0_10[228]},
      {stage1_10[94]}
   );
   gpc1_1 gpc331 (
      {stage0_10[229]},
      {stage1_10[95]}
   );
   gpc1_1 gpc332 (
      {stage0_10[230]},
      {stage1_10[96]}
   );
   gpc1_1 gpc333 (
      {stage0_10[231]},
      {stage1_10[97]}
   );
   gpc1_1 gpc334 (
      {stage0_10[232]},
      {stage1_10[98]}
   );
   gpc1_1 gpc335 (
      {stage0_10[233]},
      {stage1_10[99]}
   );
   gpc1_1 gpc336 (
      {stage0_10[234]},
      {stage1_10[100]}
   );
   gpc1_1 gpc337 (
      {stage0_10[235]},
      {stage1_10[101]}
   );
   gpc1_1 gpc338 (
      {stage0_10[236]},
      {stage1_10[102]}
   );
   gpc1_1 gpc339 (
      {stage0_10[237]},
      {stage1_10[103]}
   );
   gpc1_1 gpc340 (
      {stage0_10[238]},
      {stage1_10[104]}
   );
   gpc1_1 gpc341 (
      {stage0_10[239]},
      {stage1_10[105]}
   );
   gpc1_1 gpc342 (
      {stage0_10[240]},
      {stage1_10[106]}
   );
   gpc1_1 gpc343 (
      {stage0_10[241]},
      {stage1_10[107]}
   );
   gpc1_1 gpc344 (
      {stage0_10[242]},
      {stage1_10[108]}
   );
   gpc1_1 gpc345 (
      {stage0_10[243]},
      {stage1_10[109]}
   );
   gpc1_1 gpc346 (
      {stage0_10[244]},
      {stage1_10[110]}
   );
   gpc1_1 gpc347 (
      {stage0_10[245]},
      {stage1_10[111]}
   );
   gpc1_1 gpc348 (
      {stage0_10[246]},
      {stage1_10[112]}
   );
   gpc1_1 gpc349 (
      {stage0_10[247]},
      {stage1_10[113]}
   );
   gpc1_1 gpc350 (
      {stage0_10[248]},
      {stage1_10[114]}
   );
   gpc1_1 gpc351 (
      {stage0_10[249]},
      {stage1_10[115]}
   );
   gpc1_1 gpc352 (
      {stage0_10[250]},
      {stage1_10[116]}
   );
   gpc1_1 gpc353 (
      {stage0_10[251]},
      {stage1_10[117]}
   );
   gpc1_1 gpc354 (
      {stage0_10[252]},
      {stage1_10[118]}
   );
   gpc1_1 gpc355 (
      {stage0_10[253]},
      {stage1_10[119]}
   );
   gpc1_1 gpc356 (
      {stage0_10[254]},
      {stage1_10[120]}
   );
   gpc1_1 gpc357 (
      {stage0_10[255]},
      {stage1_10[121]}
   );
   gpc1_1 gpc358 (
      {stage0_11[252]},
      {stage1_11[79]}
   );
   gpc1_1 gpc359 (
      {stage0_11[253]},
      {stage1_11[80]}
   );
   gpc1_1 gpc360 (
      {stage0_11[254]},
      {stage1_11[81]}
   );
   gpc1_1 gpc361 (
      {stage0_11[255]},
      {stage1_11[82]}
   );
   gpc1163_5 gpc362 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc363 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc364 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc365 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc366 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc367 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc368 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc369 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc370 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc371 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc372 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc373 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc374 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc7_3 gpc375 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77], stage1_1[78]},
      {stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc376 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[13],stage2_3[14],stage2_2[14]}
   );
   gpc606_5 gpc377 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[14],stage2_3[15],stage2_2[15]}
   );
   gpc606_5 gpc378 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[15],stage2_3[16],stage2_2[16]}
   );
   gpc606_5 gpc379 (
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[16],stage2_3[17],stage2_2[17]}
   );
   gpc606_5 gpc380 (
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[17],stage2_3[18],stage2_2[18]}
   );
   gpc606_5 gpc381 (
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[18],stage2_3[19],stage2_2[19]}
   );
   gpc606_5 gpc382 (
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[19],stage2_3[20],stage2_2[20]}
   );
   gpc606_5 gpc383 (
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[20],stage2_3[21],stage2_2[21]}
   );
   gpc606_5 gpc384 (
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[8],stage2_4[21],stage2_3[22],stage2_2[22]}
   );
   gpc606_5 gpc385 (
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[9],stage2_4[22],stage2_3[23],stage2_2[23]}
   );
   gpc606_5 gpc386 (
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[10],stage2_4[23],stage2_3[24],stage2_2[24]}
   );
   gpc615_5 gpc387 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[66]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[11],stage2_5[11],stage2_4[24],stage2_3[25]}
   );
   gpc615_5 gpc388 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[67]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[12],stage2_5[12],stage2_4[25],stage2_3[26]}
   );
   gpc615_5 gpc389 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[68]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[13],stage2_5[13],stage2_4[26],stage2_3[27]}
   );
   gpc615_5 gpc390 (
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_4[69]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[14],stage2_5[14],stage2_4[27],stage2_3[28]}
   );
   gpc615_5 gpc391 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[70]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[15],stage2_5[15],stage2_4[28],stage2_3[29]}
   );
   gpc615_5 gpc392 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[71]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[16],stage2_5[16],stage2_4[29],stage2_3[30]}
   );
   gpc615_5 gpc393 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[72]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[17],stage2_5[17],stage2_4[30],stage2_3[31]}
   );
   gpc615_5 gpc394 (
      {stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage1_4[73]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[18],stage2_5[18],stage2_4[31],stage2_3[32]}
   );
   gpc615_5 gpc395 (
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56]},
      {stage1_4[74]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[19],stage2_5[19],stage2_4[32],stage2_3[33]}
   );
   gpc615_5 gpc396 (
      {stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage1_4[75]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[20],stage2_5[20],stage2_4[33],stage2_3[34]}
   );
   gpc615_5 gpc397 (
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66]},
      {stage1_4[76]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[21],stage2_5[21],stage2_4[34],stage2_3[35]}
   );
   gpc615_5 gpc398 (
      {stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage1_4[77]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[22],stage2_5[22],stage2_4[35],stage2_3[36]}
   );
   gpc615_5 gpc399 (
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_4[78]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[23],stage2_5[23],stage2_4[36],stage2_3[37]}
   );
   gpc615_5 gpc400 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage1_4[79]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[24],stage2_5[24],stage2_4[37],stage2_3[38]}
   );
   gpc615_5 gpc401 (
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86]},
      {stage1_4[80]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[25],stage2_5[25],stage2_4[38],stage2_3[39]}
   );
   gpc615_5 gpc402 (
      {stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91]},
      {stage1_4[81]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[26],stage2_5[26],stage2_4[39],stage2_3[40]}
   );
   gpc615_5 gpc403 (
      {stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95], stage1_3[96]},
      {stage1_4[82]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[27],stage2_5[27],stage2_4[40],stage2_3[41]}
   );
   gpc606_5 gpc404 (
      {stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[17],stage2_6[28],stage2_5[28],stage2_4[41]}
   );
   gpc606_5 gpc405 (
      {stage1_4[89], stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[18],stage2_6[29],stage2_5[29],stage2_4[42]}
   );
   gpc606_5 gpc406 (
      {stage1_4[95], stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[19],stage2_6[30],stage2_5[30],stage2_4[43]}
   );
   gpc606_5 gpc407 (
      {stage1_4[101], stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[20],stage2_6[31],stage2_5[31],stage2_4[44]}
   );
   gpc606_5 gpc408 (
      {stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[21],stage2_6[32],stage2_5[32],stage2_4[45]}
   );
   gpc606_5 gpc409 (
      {stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[22],stage2_6[33],stage2_5[33],stage2_4[46]}
   );
   gpc606_5 gpc410 (
      {stage1_4[119], stage1_4[120], stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[23],stage2_6[34],stage2_5[34],stage2_4[47]}
   );
   gpc606_5 gpc411 (
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[7],stage2_7[24],stage2_6[35],stage2_5[35]}
   );
   gpc606_5 gpc412 (
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[8],stage2_7[25],stage2_6[36],stage2_5[36]}
   );
   gpc606_5 gpc413 (
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[9],stage2_7[26],stage2_6[37],stage2_5[37]}
   );
   gpc606_5 gpc414 (
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[10],stage2_7[27],stage2_6[38],stage2_5[38]}
   );
   gpc615_5 gpc415 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46]},
      {stage1_7[24]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[4],stage2_8[11],stage2_7[28],stage2_6[39]}
   );
   gpc615_5 gpc416 (
      {stage1_6[47], stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51]},
      {stage1_7[25]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[5],stage2_8[12],stage2_7[29],stage2_6[40]}
   );
   gpc615_5 gpc417 (
      {stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55], stage1_6[56]},
      {stage1_7[26]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[6],stage2_8[13],stage2_7[30],stage2_6[41]}
   );
   gpc615_5 gpc418 (
      {stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60], stage1_6[61]},
      {stage1_7[27]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[7],stage2_8[14],stage2_7[31],stage2_6[42]}
   );
   gpc615_5 gpc419 (
      {stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage1_7[28]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[8],stage2_8[15],stage2_7[32],stage2_6[43]}
   );
   gpc615_5 gpc420 (
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage1_7[29]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[9],stage2_8[16],stage2_7[33],stage2_6[44]}
   );
   gpc615_5 gpc421 (
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76]},
      {stage1_7[30]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[10],stage2_8[17],stage2_7[34],stage2_6[45]}
   );
   gpc615_5 gpc422 (
      {stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81]},
      {stage1_7[31]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[11],stage2_8[18],stage2_7[35],stage2_6[46]}
   );
   gpc615_5 gpc423 (
      {stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage1_8[48]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[8],stage2_9[12],stage2_8[19],stage2_7[36]}
   );
   gpc615_5 gpc424 (
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage1_8[49]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[9],stage2_9[13],stage2_8[20],stage2_7[37]}
   );
   gpc615_5 gpc425 (
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46]},
      {stage1_8[50]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[10],stage2_9[14],stage2_8[21],stage2_7[38]}
   );
   gpc615_5 gpc426 (
      {stage1_7[47], stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51]},
      {stage1_8[51]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[11],stage2_9[15],stage2_8[22],stage2_7[39]}
   );
   gpc615_5 gpc427 (
      {stage1_7[52], stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56]},
      {stage1_8[52]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[12],stage2_9[16],stage2_8[23],stage2_7[40]}
   );
   gpc615_5 gpc428 (
      {stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61]},
      {stage1_8[53]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[13],stage2_9[17],stage2_8[24],stage2_7[41]}
   );
   gpc615_5 gpc429 (
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage1_8[54]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[14],stage2_9[18],stage2_8[25],stage2_7[42]}
   );
   gpc615_5 gpc430 (
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage1_8[55]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[15],stage2_9[19],stage2_8[26],stage2_7[43]}
   );
   gpc615_5 gpc431 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[56]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[16],stage2_9[20],stage2_8[27],stage2_7[44]}
   );
   gpc615_5 gpc432 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[57]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[17],stage2_9[21],stage2_8[28],stage2_7[45]}
   );
   gpc615_5 gpc433 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[58]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[18],stage2_9[22],stage2_8[29],stage2_7[46]}
   );
   gpc615_5 gpc434 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], 1'b0},
      {stage1_8[59]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[19],stage2_9[23],stage2_8[30],stage2_7[47]}
   );
   gpc606_5 gpc435 (
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[12],stage2_10[20],stage2_9[24],stage2_8[31]}
   );
   gpc606_5 gpc436 (
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[13],stage2_10[21],stage2_9[25],stage2_8[32]}
   );
   gpc606_5 gpc437 (
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[14],stage2_10[22],stage2_9[26],stage2_8[33]}
   );
   gpc606_5 gpc438 (
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[15],stage2_10[23],stage2_9[27],stage2_8[34]}
   );
   gpc606_5 gpc439 (
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[16],stage2_10[24],stage2_9[28],stage2_8[35]}
   );
   gpc606_5 gpc440 (
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[17],stage2_10[25],stage2_9[29],stage2_8[36]}
   );
   gpc606_5 gpc441 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[18],stage2_10[26],stage2_9[30],stage2_8[37]}
   );
   gpc606_5 gpc442 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[19],stage2_10[27],stage2_9[31],stage2_8[38]}
   );
   gpc606_5 gpc443 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[20],stage2_10[28],stage2_9[32],stage2_8[39]}
   );
   gpc606_5 gpc444 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[21],stage2_10[29],stage2_9[33],stage2_8[40]}
   );
   gpc606_5 gpc445 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[22],stage2_10[30],stage2_9[34],stage2_8[41]}
   );
   gpc606_5 gpc446 (
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[11],stage2_11[23],stage2_10[31],stage2_9[35]}
   );
   gpc606_5 gpc447 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[12],stage2_11[24],stage2_10[32],stage2_9[36]}
   );
   gpc606_5 gpc448 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[13],stage2_11[25],stage2_10[33],stage2_9[37]}
   );
   gpc606_5 gpc449 (
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[14],stage2_11[26],stage2_10[34],stage2_9[38]}
   );
   gpc606_5 gpc450 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[15],stage2_11[27],stage2_10[35],stage2_9[39]}
   );
   gpc606_5 gpc451 (
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[16],stage2_11[28],stage2_10[36],stage2_9[40]}
   );
   gpc606_5 gpc452 (
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[17],stage2_11[29],stage2_10[37],stage2_9[41]}
   );
   gpc606_5 gpc453 (
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[18],stage2_11[30],stage2_10[38],stage2_9[42]}
   );
   gpc606_5 gpc454 (
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[8],stage2_12[19],stage2_11[31],stage2_10[39]}
   );
   gpc615_5 gpc455 (
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76]},
      {stage1_11[48]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[9],stage2_12[20],stage2_11[32],stage2_10[40]}
   );
   gpc615_5 gpc456 (
      {stage1_10[77], stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81]},
      {stage1_11[49]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[10],stage2_12[21],stage2_11[33],stage2_10[41]}
   );
   gpc615_5 gpc457 (
      {stage1_10[82], stage1_10[83], stage1_10[84], stage1_10[85], stage1_10[86]},
      {stage1_11[50]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[11],stage2_12[22],stage2_11[34],stage2_10[42]}
   );
   gpc615_5 gpc458 (
      {stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90], stage1_10[91]},
      {stage1_11[51]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[12],stage2_12[23],stage2_11[35],stage2_10[43]}
   );
   gpc615_5 gpc459 (
      {stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96]},
      {stage1_11[52]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[13],stage2_12[24],stage2_11[36],stage2_10[44]}
   );
   gpc615_5 gpc460 (
      {stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage1_11[53]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[14],stage2_12[25],stage2_11[37],stage2_10[45]}
   );
   gpc615_5 gpc461 (
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_11[54]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[15],stage2_12[26],stage2_11[38],stage2_10[46]}
   );
   gpc615_5 gpc462 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111]},
      {stage1_11[55]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[16],stage2_12[27],stage2_11[39],stage2_10[47]}
   );
   gpc615_5 gpc463 (
      {stage1_10[112], stage1_10[113], stage1_10[114], stage1_10[115], stage1_10[116]},
      {stage1_11[56]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[17],stage2_12[28],stage2_11[40],stage2_10[48]}
   );
   gpc615_5 gpc464 (
      {stage1_10[117], stage1_10[118], stage1_10[119], stage1_10[120], stage1_10[121]},
      {stage1_11[57]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[18],stage2_12[29],stage2_11[41],stage2_10[49]}
   );
   gpc615_5 gpc465 (
      {stage1_11[58], stage1_11[59], stage1_11[60], stage1_11[61], stage1_11[62]},
      {stage1_12[66]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[11],stage2_13[19],stage2_12[30],stage2_11[42]}
   );
   gpc615_5 gpc466 (
      {stage1_11[63], stage1_11[64], stage1_11[65], stage1_11[66], stage1_11[67]},
      {stage1_12[67]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[12],stage2_13[20],stage2_12[31],stage2_11[43]}
   );
   gpc615_5 gpc467 (
      {stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72]},
      {stage1_12[68]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[13],stage2_13[21],stage2_12[32],stage2_11[44]}
   );
   gpc615_5 gpc468 (
      {stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage1_12[69]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[14],stage2_13[22],stage2_12[33],stage2_11[45]}
   );
   gpc615_5 gpc469 (
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82]},
      {stage1_12[70]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[15],stage2_13[23],stage2_12[34],stage2_11[46]}
   );
   gpc1_1 gpc470 (
      {stage1_0[42]},
      {stage2_0[13]}
   );
   gpc1_1 gpc471 (
      {stage1_0[43]},
      {stage2_0[14]}
   );
   gpc1_1 gpc472 (
      {stage1_0[44]},
      {stage2_0[15]}
   );
   gpc1_1 gpc473 (
      {stage1_0[45]},
      {stage2_0[16]}
   );
   gpc1_1 gpc474 (
      {stage1_0[46]},
      {stage2_0[17]}
   );
   gpc1_1 gpc475 (
      {stage1_0[47]},
      {stage2_0[18]}
   );
   gpc1_1 gpc476 (
      {stage1_1[79]},
      {stage2_1[14]}
   );
   gpc1_1 gpc477 (
      {stage1_1[80]},
      {stage2_1[15]}
   );
   gpc1_1 gpc478 (
      {stage1_1[81]},
      {stage2_1[16]}
   );
   gpc1_1 gpc479 (
      {stage1_1[82]},
      {stage2_1[17]}
   );
   gpc1_1 gpc480 (
      {stage1_1[83]},
      {stage2_1[18]}
   );
   gpc1_1 gpc481 (
      {stage1_1[84]},
      {stage2_1[19]}
   );
   gpc1_1 gpc482 (
      {stage1_1[85]},
      {stage2_1[20]}
   );
   gpc1_1 gpc483 (
      {stage1_1[86]},
      {stage2_1[21]}
   );
   gpc1_1 gpc484 (
      {stage1_1[87]},
      {stage2_1[22]}
   );
   gpc1_1 gpc485 (
      {stage1_1[88]},
      {stage2_1[23]}
   );
   gpc1_1 gpc486 (
      {stage1_1[89]},
      {stage2_1[24]}
   );
   gpc1_1 gpc487 (
      {stage1_2[84]},
      {stage2_2[25]}
   );
   gpc1_1 gpc488 (
      {stage1_4[125]},
      {stage2_4[48]}
   );
   gpc1_1 gpc489 (
      {stage1_4[126]},
      {stage2_4[49]}
   );
   gpc1_1 gpc490 (
      {stage1_5[126]},
      {stage2_5[39]}
   );
   gpc1_1 gpc491 (
      {stage1_5[127]},
      {stage2_5[40]}
   );
   gpc1_1 gpc492 (
      {stage1_5[128]},
      {stage2_5[41]}
   );
   gpc1_1 gpc493 (
      {stage1_6[82]},
      {stage2_6[47]}
   );
   gpc1_1 gpc494 (
      {stage1_6[83]},
      {stage2_6[48]}
   );
   gpc1_1 gpc495 (
      {stage1_6[84]},
      {stage2_6[49]}
   );
   gpc1_1 gpc496 (
      {stage1_6[85]},
      {stage2_6[50]}
   );
   gpc1_1 gpc497 (
      {stage1_6[86]},
      {stage2_6[51]}
   );
   gpc1_1 gpc498 (
      {stage1_6[87]},
      {stage2_6[52]}
   );
   gpc1_1 gpc499 (
      {stage1_6[88]},
      {stage2_6[53]}
   );
   gpc1_1 gpc500 (
      {stage1_8[126]},
      {stage2_8[42]}
   );
   gpc1_1 gpc501 (
      {stage1_8[127]},
      {stage2_8[43]}
   );
   gpc1_1 gpc502 (
      {stage1_8[128]},
      {stage2_8[44]}
   );
   gpc1_1 gpc503 (
      {stage1_8[129]},
      {stage2_8[45]}
   );
   gpc1_1 gpc504 (
      {stage1_8[130]},
      {stage2_8[46]}
   );
   gpc1_1 gpc505 (
      {stage1_8[131]},
      {stage2_8[47]}
   );
   gpc1_1 gpc506 (
      {stage1_8[132]},
      {stage2_8[48]}
   );
   gpc1_1 gpc507 (
      {stage1_8[133]},
      {stage2_8[49]}
   );
   gpc1_1 gpc508 (
      {stage1_8[134]},
      {stage2_8[50]}
   );
   gpc1_1 gpc509 (
      {stage1_8[135]},
      {stage2_8[51]}
   );
   gpc1_1 gpc510 (
      {stage1_8[136]},
      {stage2_8[52]}
   );
   gpc1_1 gpc511 (
      {stage1_8[137]},
      {stage2_8[53]}
   );
   gpc1_1 gpc512 (
      {stage1_8[138]},
      {stage2_8[54]}
   );
   gpc1_1 gpc513 (
      {stage1_8[139]},
      {stage2_8[55]}
   );
   gpc1_1 gpc514 (
      {stage1_8[140]},
      {stage2_8[56]}
   );
   gpc1_1 gpc515 (
      {stage1_8[141]},
      {stage2_8[57]}
   );
   gpc1_1 gpc516 (
      {stage1_8[142]},
      {stage2_8[58]}
   );
   gpc1_1 gpc517 (
      {stage1_8[143]},
      {stage2_8[59]}
   );
   gpc1_1 gpc518 (
      {stage1_8[144]},
      {stage2_8[60]}
   );
   gpc1_1 gpc519 (
      {stage1_8[145]},
      {stage2_8[61]}
   );
   gpc1_1 gpc520 (
      {stage1_8[146]},
      {stage2_8[62]}
   );
   gpc1_1 gpc521 (
      {stage1_8[147]},
      {stage2_8[63]}
   );
   gpc1_1 gpc522 (
      {stage1_8[148]},
      {stage2_8[64]}
   );
   gpc1_1 gpc523 (
      {stage1_8[149]},
      {stage2_8[65]}
   );
   gpc1_1 gpc524 (
      {stage1_8[150]},
      {stage2_8[66]}
   );
   gpc1_1 gpc525 (
      {stage1_8[151]},
      {stage2_8[67]}
   );
   gpc1_1 gpc526 (
      {stage1_8[152]},
      {stage2_8[68]}
   );
   gpc1_1 gpc527 (
      {stage1_8[153]},
      {stage2_8[69]}
   );
   gpc1_1 gpc528 (
      {stage1_8[154]},
      {stage2_8[70]}
   );
   gpc1_1 gpc529 (
      {stage1_12[71]},
      {stage2_12[35]}
   );
   gpc1_1 gpc530 (
      {stage1_13[30]},
      {stage2_13[24]}
   );
   gpc1_1 gpc531 (
      {stage1_13[31]},
      {stage2_13[25]}
   );
   gpc1_1 gpc532 (
      {stage1_13[32]},
      {stage2_13[26]}
   );
   gpc1_1 gpc533 (
      {stage1_13[33]},
      {stage2_13[27]}
   );
   gpc1_1 gpc534 (
      {stage1_13[34]},
      {stage2_13[28]}
   );
   gpc1_1 gpc535 (
      {stage1_13[35]},
      {stage2_13[29]}
   );
   gpc1_1 gpc536 (
      {stage1_13[36]},
      {stage2_13[30]}
   );
   gpc1_1 gpc537 (
      {stage1_13[37]},
      {stage2_13[31]}
   );
   gpc1_1 gpc538 (
      {stage1_13[38]},
      {stage2_13[32]}
   );
   gpc1_1 gpc539 (
      {stage1_13[39]},
      {stage2_13[33]}
   );
   gpc1_1 gpc540 (
      {stage1_13[40]},
      {stage2_13[34]}
   );
   gpc1_1 gpc541 (
      {stage1_13[41]},
      {stage2_13[35]}
   );
   gpc606_5 gpc542 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc543 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc606_5 gpc544 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc545 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[3],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc546 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[4],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc547 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[24]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[5],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc615_5 gpc548 (
      {stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15]},
      {stage2_3[25]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[6],stage3_4[6],stage3_3[6],stage3_2[6]}
   );
   gpc615_5 gpc549 (
      {stage2_2[16], stage2_2[17], stage2_2[18], stage2_2[19], stage2_2[20]},
      {stage2_3[26]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[7],stage3_4[7],stage3_3[7],stage3_2[7]}
   );
   gpc615_5 gpc550 (
      {stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31]},
      {stage2_4[24]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[4],stage3_5[8],stage3_4[8],stage3_3[8]}
   );
   gpc615_5 gpc551 (
      {stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage2_4[25]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[5],stage3_5[9],stage3_4[9],stage3_3[9]}
   );
   gpc615_5 gpc552 (
      {stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40], stage2_3[41]},
      {stage2_4[26]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[6],stage3_5[10],stage3_4[10],stage3_3[10]}
   );
   gpc606_5 gpc553 (
      {stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31], stage2_4[32]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[7],stage3_5[11],stage3_4[11]}
   );
   gpc606_5 gpc554 (
      {stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37], stage2_4[38]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[8],stage3_5[12],stage3_4[12]}
   );
   gpc606_5 gpc555 (
      {stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42], stage2_4[43], stage2_4[44]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[9],stage3_5[13],stage3_4[13]}
   );
   gpc606_5 gpc556 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[3],stage3_7[6],stage3_6[10],stage3_5[14]}
   );
   gpc606_5 gpc557 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[4],stage3_7[7],stage3_6[11],stage3_5[15]}
   );
   gpc606_5 gpc558 (
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[5],stage3_7[8],stage3_6[12],stage3_5[16]}
   );
   gpc606_5 gpc559 (
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[6],stage3_7[9],stage3_6[13],stage3_5[17]}
   );
   gpc606_5 gpc560 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[4],stage3_8[7],stage3_7[10],stage3_6[14]}
   );
   gpc606_5 gpc561 (
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[5],stage3_8[8],stage3_7[11],stage3_6[15]}
   );
   gpc606_5 gpc562 (
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[6],stage3_8[9],stage3_7[12],stage3_6[16]}
   );
   gpc615_5 gpc563 (
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40]},
      {stage2_7[24]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[7],stage3_8[10],stage3_7[13],stage3_6[17]}
   );
   gpc615_5 gpc564 (
      {stage2_6[41], stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45]},
      {stage2_7[25]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[8],stage3_8[11],stage3_7[14],stage3_6[18]}
   );
   gpc615_5 gpc565 (
      {stage2_6[46], stage2_6[47], stage2_6[48], stage2_6[49], stage2_6[50]},
      {stage2_7[26]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[9],stage3_8[12],stage3_7[15],stage3_6[19]}
   );
   gpc615_5 gpc566 (
      {stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage2_8[36]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[6],stage3_9[10],stage3_8[13],stage3_7[16]}
   );
   gpc615_5 gpc567 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[37]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[7],stage3_9[11],stage3_8[14],stage3_7[17]}
   );
   gpc615_5 gpc568 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[38]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[8],stage3_9[12],stage3_8[15],stage3_7[18]}
   );
   gpc615_5 gpc569 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[39]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[9],stage3_9[13],stage3_8[16],stage3_7[19]}
   );
   gpc615_5 gpc570 (
      {stage2_8[40], stage2_8[41], stage2_8[42], stage2_8[43], stage2_8[44]},
      {stage2_9[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[10],stage3_9[14],stage3_8[17]}
   );
   gpc615_5 gpc571 (
      {stage2_8[45], stage2_8[46], stage2_8[47], stage2_8[48], stage2_8[49]},
      {stage2_9[25]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[11],stage3_9[15],stage3_8[18]}
   );
   gpc615_5 gpc572 (
      {stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54]},
      {stage2_9[26]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[12],stage3_9[16],stage3_8[19]}
   );
   gpc615_5 gpc573 (
      {stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage2_9[27]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[7],stage3_10[13],stage3_9[17],stage3_8[20]}
   );
   gpc615_5 gpc574 (
      {stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64]},
      {stage2_9[28]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[8],stage3_10[14],stage3_9[18],stage3_8[21]}
   );
   gpc615_5 gpc575 (
      {stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69]},
      {stage2_9[29]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[9],stage3_10[15],stage3_9[19],stage3_8[22]}
   );
   gpc606_5 gpc576 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[6],stage3_11[10],stage3_10[16],stage3_9[20]}
   );
   gpc615_5 gpc577 (
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40]},
      {stage2_11[6]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[7],stage3_11[11],stage3_10[17]}
   );
   gpc615_5 gpc578 (
      {stage2_10[41], stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45]},
      {stage2_11[7]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[2],stage3_12[8],stage3_11[12],stage3_10[18]}
   );
   gpc615_5 gpc579 (
      {stage2_10[46], stage2_10[47], stage2_10[48], stage2_10[49], 1'b0},
      {stage2_11[8]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[3],stage3_12[9],stage3_11[13],stage3_10[19]}
   );
   gpc606_5 gpc580 (
      {stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[4],stage3_12[10],stage3_11[14]}
   );
   gpc606_5 gpc581 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[5],stage3_12[11],stage3_11[15]}
   );
   gpc606_5 gpc582 (
      {stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[6],stage3_12[12],stage3_11[16]}
   );
   gpc606_5 gpc583 (
      {stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[6],stage3_13[7],stage3_12[13],stage3_11[17]}
   );
   gpc606_5 gpc584 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[7],stage3_13[8],stage3_12[14],stage3_11[18]}
   );
   gpc606_5 gpc585 (
      {stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[8],stage3_13[9],stage3_12[15],stage3_11[19]}
   );
   gpc1406_5 gpc586 (
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[6],stage3_14[9],stage3_13[10],stage3_12[16]}
   );
   gpc606_5 gpc587 (
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage2_14[4], stage2_14[5], stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9]},
      {stage3_16[1],stage3_15[7],stage3_14[10],stage3_13[11],stage3_12[17]}
   );
   gpc606_5 gpc588 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[10], stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage3_16[2],stage3_15[8],stage3_14[11],stage3_13[12],stage3_12[18]}
   );
   gpc1_1 gpc589 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc590 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc591 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc592 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc593 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc594 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc595 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc596 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc597 (
      {stage2_0[8]},
      {stage3_0[8]}
   );
   gpc1_1 gpc598 (
      {stage2_0[9]},
      {stage3_0[9]}
   );
   gpc1_1 gpc599 (
      {stage2_0[10]},
      {stage3_0[10]}
   );
   gpc1_1 gpc600 (
      {stage2_0[11]},
      {stage3_0[11]}
   );
   gpc1_1 gpc601 (
      {stage2_0[12]},
      {stage3_0[12]}
   );
   gpc1_1 gpc602 (
      {stage2_0[13]},
      {stage3_0[13]}
   );
   gpc1_1 gpc603 (
      {stage2_0[14]},
      {stage3_0[14]}
   );
   gpc1_1 gpc604 (
      {stage2_0[15]},
      {stage3_0[15]}
   );
   gpc1_1 gpc605 (
      {stage2_0[16]},
      {stage3_0[16]}
   );
   gpc1_1 gpc606 (
      {stage2_0[17]},
      {stage3_0[17]}
   );
   gpc1_1 gpc607 (
      {stage2_0[18]},
      {stage3_0[18]}
   );
   gpc1_1 gpc608 (
      {stage2_1[24]},
      {stage3_1[4]}
   );
   gpc1_1 gpc609 (
      {stage2_2[21]},
      {stage3_2[8]}
   );
   gpc1_1 gpc610 (
      {stage2_2[22]},
      {stage3_2[9]}
   );
   gpc1_1 gpc611 (
      {stage2_2[23]},
      {stage3_2[10]}
   );
   gpc1_1 gpc612 (
      {stage2_2[24]},
      {stage3_2[11]}
   );
   gpc1_1 gpc613 (
      {stage2_2[25]},
      {stage3_2[12]}
   );
   gpc1_1 gpc614 (
      {stage2_4[45]},
      {stage3_4[14]}
   );
   gpc1_1 gpc615 (
      {stage2_4[46]},
      {stage3_4[15]}
   );
   gpc1_1 gpc616 (
      {stage2_4[47]},
      {stage3_4[16]}
   );
   gpc1_1 gpc617 (
      {stage2_4[48]},
      {stage3_4[17]}
   );
   gpc1_1 gpc618 (
      {stage2_4[49]},
      {stage3_4[18]}
   );
   gpc1_1 gpc619 (
      {stage2_6[51]},
      {stage3_6[20]}
   );
   gpc1_1 gpc620 (
      {stage2_6[52]},
      {stage3_6[21]}
   );
   gpc1_1 gpc621 (
      {stage2_6[53]},
      {stage3_6[22]}
   );
   gpc1_1 gpc622 (
      {stage2_7[47]},
      {stage3_7[20]}
   );
   gpc1_1 gpc623 (
      {stage2_8[70]},
      {stage3_8[23]}
   );
   gpc1_1 gpc624 (
      {stage2_9[36]},
      {stage3_9[21]}
   );
   gpc1_1 gpc625 (
      {stage2_9[37]},
      {stage3_9[22]}
   );
   gpc1_1 gpc626 (
      {stage2_9[38]},
      {stage3_9[23]}
   );
   gpc1_1 gpc627 (
      {stage2_9[39]},
      {stage3_9[24]}
   );
   gpc1_1 gpc628 (
      {stage2_9[40]},
      {stage3_9[25]}
   );
   gpc1_1 gpc629 (
      {stage2_9[41]},
      {stage3_9[26]}
   );
   gpc1_1 gpc630 (
      {stage2_9[42]},
      {stage3_9[27]}
   );
   gpc1_1 gpc631 (
      {stage2_11[45]},
      {stage3_11[20]}
   );
   gpc1_1 gpc632 (
      {stage2_11[46]},
      {stage3_11[21]}
   );
   gpc1_1 gpc633 (
      {stage2_15[1]},
      {stage3_15[9]}
   );
   gpc1_1 gpc634 (
      {stage2_15[2]},
      {stage3_15[10]}
   );
   gpc1_1 gpc635 (
      {stage2_15[3]},
      {stage3_15[11]}
   );
   gpc1_1 gpc636 (
      {stage2_15[4]},
      {stage3_15[12]}
   );
   gpc606_5 gpc637 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc638 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc2135_5 gpc639 (
      {stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage3_4[6], stage3_4[7], stage3_4[8]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc2135_5 gpc640 (
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10]},
      {stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_5[1]},
      {stage3_6[2], stage3_6[3]},
      {stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[3],stage4_3[3]}
   );
   gpc615_5 gpc641 (
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16]},
      {stage3_5[2]},
      {stage3_6[4], stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage4_8[0],stage4_7[2],stage4_6[3],stage4_5[3],stage4_4[4]}
   );
   gpc615_5 gpc642 (
      {stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6], stage3_5[7]},
      {stage3_6[10]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[4],stage4_5[4]}
   );
   gpc615_5 gpc643 (
      {stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11], stage3_5[12]},
      {stage3_6[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[4],stage4_6[5],stage4_5[5]}
   );
   gpc615_5 gpc644 (
      {stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_6[12]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[3],stage4_7[5],stage4_6[6],stage4_5[6]}
   );
   gpc2135_5 gpc645 (
      {stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage3_7[18], stage3_7[19], stage3_7[20]},
      {stage3_8[0]},
      {stage3_9[0], stage3_9[1]},
      {stage4_10[0],stage4_9[3],stage4_8[4],stage4_7[6],stage4_6[7]}
   );
   gpc135_4 gpc646 (
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[1],stage4_9[4],stage4_8[5]}
   );
   gpc135_4 gpc647 (
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10]},
      {stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_10[1]},
      {stage4_11[1],stage4_10[2],stage4_9[5],stage4_8[6]}
   );
   gpc615_5 gpc648 (
      {stage3_8[11], stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15]},
      {stage3_9[8]},
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage4_12[0],stage4_11[2],stage4_10[3],stage4_9[6],stage4_8[7]}
   );
   gpc615_5 gpc649 (
      {stage3_8[16], stage3_8[17], stage3_8[18], stage3_8[19], stage3_8[20]},
      {stage3_9[9]},
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage4_12[1],stage4_11[3],stage4_10[4],stage4_9[7],stage4_8[8]}
   );
   gpc606_5 gpc650 (
      {stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[4],stage4_10[5],stage4_9[8]}
   );
   gpc606_5 gpc651 (
      {stage3_9[16], stage3_9[17], stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[3],stage4_11[5],stage4_10[6],stage4_9[9]}
   );
   gpc606_5 gpc652 (
      {stage3_9[22], stage3_9[23], stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[4],stage4_11[6],stage4_10[7],stage4_9[10]}
   );
   gpc606_5 gpc653 (
      {stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[3],stage4_12[5],stage4_11[7],stage4_10[8]}
   );
   gpc606_5 gpc654 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[4],stage4_12[6]}
   );
   gpc606_5 gpc655 (
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[1],stage4_14[2],stage4_13[5],stage4_12[7]}
   );
   gpc1406_5 gpc656 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[2],stage4_15[2],stage4_14[3],stage4_13[6]}
   );
   gpc2116_5 gpc657 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {1'b0},
      {stage3_15[4]},
      {stage3_16[1], stage3_16[2]},
      {stage4_17[1],stage4_16[3],stage4_15[3],stage4_14[4],stage4_13[7]}
   );
   gpc1_1 gpc658 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc659 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc660 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc661 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc662 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc663 (
      {stage3_0[11]},
      {stage4_0[6]}
   );
   gpc1_1 gpc664 (
      {stage3_0[12]},
      {stage4_0[7]}
   );
   gpc1_1 gpc665 (
      {stage3_0[13]},
      {stage4_0[8]}
   );
   gpc1_1 gpc666 (
      {stage3_0[14]},
      {stage4_0[9]}
   );
   gpc1_1 gpc667 (
      {stage3_0[15]},
      {stage4_0[10]}
   );
   gpc1_1 gpc668 (
      {stage3_0[16]},
      {stage4_0[11]}
   );
   gpc1_1 gpc669 (
      {stage3_0[17]},
      {stage4_0[12]}
   );
   gpc1_1 gpc670 (
      {stage3_0[18]},
      {stage4_0[13]}
   );
   gpc1_1 gpc671 (
      {stage3_1[0]},
      {stage4_1[1]}
   );
   gpc1_1 gpc672 (
      {stage3_1[1]},
      {stage4_1[2]}
   );
   gpc1_1 gpc673 (
      {stage3_1[2]},
      {stage4_1[3]}
   );
   gpc1_1 gpc674 (
      {stage3_1[3]},
      {stage4_1[4]}
   );
   gpc1_1 gpc675 (
      {stage3_1[4]},
      {stage4_1[5]}
   );
   gpc1_1 gpc676 (
      {stage3_2[11]},
      {stage4_2[2]}
   );
   gpc1_1 gpc677 (
      {stage3_2[12]},
      {stage4_2[3]}
   );
   gpc1_1 gpc678 (
      {stage3_4[17]},
      {stage4_4[5]}
   );
   gpc1_1 gpc679 (
      {stage3_4[18]},
      {stage4_4[6]}
   );
   gpc1_1 gpc680 (
      {stage3_6[18]},
      {stage4_6[8]}
   );
   gpc1_1 gpc681 (
      {stage3_6[19]},
      {stage4_6[9]}
   );
   gpc1_1 gpc682 (
      {stage3_6[20]},
      {stage4_6[10]}
   );
   gpc1_1 gpc683 (
      {stage3_6[21]},
      {stage4_6[11]}
   );
   gpc1_1 gpc684 (
      {stage3_6[22]},
      {stage4_6[12]}
   );
   gpc1_1 gpc685 (
      {stage3_8[21]},
      {stage4_8[9]}
   );
   gpc1_1 gpc686 (
      {stage3_8[22]},
      {stage4_8[10]}
   );
   gpc1_1 gpc687 (
      {stage3_8[23]},
      {stage4_8[11]}
   );
   gpc1_1 gpc688 (
      {stage3_11[18]},
      {stage4_11[8]}
   );
   gpc1_1 gpc689 (
      {stage3_11[19]},
      {stage4_11[9]}
   );
   gpc1_1 gpc690 (
      {stage3_11[20]},
      {stage4_11[10]}
   );
   gpc1_1 gpc691 (
      {stage3_11[21]},
      {stage4_11[11]}
   );
   gpc1_1 gpc692 (
      {stage3_12[18]},
      {stage4_12[8]}
   );
   gpc1_1 gpc693 (
      {stage3_13[12]},
      {stage4_13[8]}
   );
   gpc1_1 gpc694 (
      {stage3_15[5]},
      {stage4_15[4]}
   );
   gpc1_1 gpc695 (
      {stage3_15[6]},
      {stage4_15[5]}
   );
   gpc1_1 gpc696 (
      {stage3_15[7]},
      {stage4_15[6]}
   );
   gpc1_1 gpc697 (
      {stage3_15[8]},
      {stage4_15[7]}
   );
   gpc1_1 gpc698 (
      {stage3_15[9]},
      {stage4_15[8]}
   );
   gpc1_1 gpc699 (
      {stage3_15[10]},
      {stage4_15[9]}
   );
   gpc1_1 gpc700 (
      {stage3_15[11]},
      {stage4_15[10]}
   );
   gpc1_1 gpc701 (
      {stage3_15[12]},
      {stage4_15[11]}
   );
   gpc2135_5 gpc702 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc2135_5 gpc703 (
      {stage4_0[5], stage4_0[6], stage4_0[7], stage4_0[8], stage4_0[9]},
      {stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_2[1]},
      {stage4_3[2], stage4_3[3]},
      {stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1],stage5_0[1]}
   );
   gpc615_5 gpc704 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4]},
      {stage4_5[0]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[2]}
   );
   gpc606_5 gpc705 (
      {stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[1]}
   );
   gpc615_5 gpc706 (
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10]},
      {stage4_7[6]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[1],stage5_8[2],stage5_7[2],stage5_6[2]}
   );
   gpc7_3 gpc707 (
      {stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], 1'b0},
      {stage5_10[1],stage5_9[2],stage5_8[3]}
   );
   gpc1343_5 gpc708 (
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[3]}
   );
   gpc1343_5 gpc709 (
      {stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage4_12[1]},
      {stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[3],stage5_9[4]}
   );
   gpc615_5 gpc710 (
      {stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10]},
      {stage4_10[8]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[2],stage5_12[2],stage5_11[2],stage5_10[4],stage5_9[5]}
   );
   gpc7_3 gpc711 (
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7], stage4_12[8]},
      {stage5_14[0],stage5_13[3],stage5_12[3]}
   );
   gpc615_5 gpc712 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4]},
      {stage4_14[0]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[1],stage5_13[4]}
   );
   gpc615_5 gpc713 (
      {stage4_13[5], stage4_13[6], stage4_13[7], stage4_13[8], 1'b0},
      {stage4_14[1]},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[2],stage5_13[5]}
   );
   gpc1_1 gpc714 (
      {stage4_0[10]},
      {stage5_0[2]}
   );
   gpc1_1 gpc715 (
      {stage4_0[11]},
      {stage5_0[3]}
   );
   gpc1_1 gpc716 (
      {stage4_0[12]},
      {stage5_0[4]}
   );
   gpc1_1 gpc717 (
      {stage4_0[13]},
      {stage5_0[5]}
   );
   gpc1_1 gpc718 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc719 (
      {stage4_2[3]},
      {stage5_2[3]}
   );
   gpc1_1 gpc720 (
      {stage4_4[5]},
      {stage5_4[3]}
   );
   gpc1_1 gpc721 (
      {stage4_4[6]},
      {stage5_4[4]}
   );
   gpc1_1 gpc722 (
      {stage4_6[11]},
      {stage5_6[3]}
   );
   gpc1_1 gpc723 (
      {stage4_6[12]},
      {stage5_6[4]}
   );
   gpc1_1 gpc724 (
      {stage4_14[2]},
      {stage5_14[3]}
   );
   gpc1_1 gpc725 (
      {stage4_14[3]},
      {stage5_14[4]}
   );
   gpc1_1 gpc726 (
      {stage4_14[4]},
      {stage5_14[5]}
   );
   gpc1_1 gpc727 (
      {stage4_16[0]},
      {stage5_16[2]}
   );
   gpc1_1 gpc728 (
      {stage4_16[1]},
      {stage5_16[3]}
   );
   gpc1_1 gpc729 (
      {stage4_16[2]},
      {stage5_16[4]}
   );
   gpc1_1 gpc730 (
      {stage4_16[3]},
      {stage5_16[5]}
   );
   gpc1_1 gpc731 (
      {stage4_17[0]},
      {stage5_17[2]}
   );
   gpc1_1 gpc732 (
      {stage4_17[1]},
      {stage5_17[3]}
   );
   gpc1325_5 gpc733 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4]},
      {stage5_1[0], stage5_1[1]},
      {stage5_2[0], stage5_2[1], stage5_2[2]},
      {stage5_3[0]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc615_5 gpc734 (
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4]},
      {stage5_5[0]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], 1'b0},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[1]}
   );
   gpc1343_5 gpc735 (
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0], stage5_9[1], stage5_9[2]},
      {stage5_10[0]},
      {stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[1],stage6_7[1]}
   );
   gpc1343_5 gpc736 (
      {stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4]},
      {stage5_11[0], stage5_11[1], stage5_11[2]},
      {stage5_12[0]},
      {stage6_13[0],stage6_12[0],stage6_11[1],stage6_10[1],stage6_9[1]}
   );
   gpc1163_5 gpc737 (
      {stage5_12[1], stage5_12[2], stage5_12[3]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[0]},
      {stage5_15[0]},
      {stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[1],stage6_12[1]}
   );
   gpc615_5 gpc738 (
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[1]},
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage6_18[0],stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[1]}
   );
   gpc117_4 gpc739 (
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], 1'b0, 1'b0, 1'b0},
      {1'b0},
      {1'b0},
      {stage6_19[0],stage6_18[1],stage6_17[1]}
   );
   gpc1_1 gpc740 (
      {stage5_0[5]},
      {stage6_0[1]}
   );
   gpc1_1 gpc741 (
      {stage5_2[3]},
      {stage6_2[1]}
   );
   gpc1_1 gpc742 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc743 (
      {stage5_5[1]},
      {stage6_5[1]}
   );
endmodule

module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor_CLA256_12 compressor_CLA256_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h984bb251b8ee46019253ebfaece327a39866908a4bbd4576c2febf91069a135f5184b84b9a03577ccc7ecb8a7db974738bbb80713b50b8d1b425162a6902aea974f766bb1002160a84f93ba9e00e37f4c6a6488510a68f36660b9a06c91c5b296d9d49c45366d89b95e710d70d028ebd24933d538df541b9e30a9291856ecf131d19e231270c47e8abc2fde49157f51921ec6d214bc38b8afccf0fed9ffd9816eb3bcdfd6a1a7b69245f9ed324a6c3bdd59cf9c10d30b457dca95e8e7cd9b8b365184108782f192e9bf90dc65b6aa5965d274b7b2145fa85c6f35ac75bc7663092e82ea0186f8a8502de3ce79cce732094a53a22fdaf5b10235014f6cc440ff300c047cebcaadd22138a9d7b3553f81b1353d9c95a316badfce1811a00d4d8d8ef64b93507ebd599a246fb389d21bd044a3206648d0cb54b6d3914c2fa20a61bb29489c299ca41d9e6b47c4a3b6b5b38546ef3764766bfacdfbbc06c3690083383eb0ef4ca72860a37bd2c558ec0bf6d12e1dcf1597bbe185bf29cbfc8e67b46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h94dbab931b762dc43c98405e89b98acdd1bae214512cb1ffd33284aeb8e6f5fed05c3da519ae14a739a51e481f858ffdf71258cf2ed1c251e3d6593cef8784314dc09aaf362b6071094423866443dfa28228a121a8fbfc8dd6e770a90cdfcf2f2c4b7816f0dcb1b9604af04d8c75b7d9569a4bf6e68b47be1ed3e7b829f0a41a1d2897b54c58d2ab6bc6e9742287810734318c0720d65dac7846c04de9b8dd578d04d3b85b6fe3c7bbfa049b31fe4fb2ca3c7379bbd366dd42f719f863091ec3faf815d1208629a656515680ed6ee123c4c7897d87e880d701b563839aff59c659b22beeeb0a1495757ee46510e09421ad519ca14256f7ee27f23b53aa1617a570a4c5475ff501f09e809ea29583fca4e2b07e48d44adde78b05ab7ac0d80c60e081d4c717c7b2797709328b7ddd835012ee21863972e8192750321d1d99987243b069e6afaa3a671aaafc5c13640c132844568e52337b9e850b91862c1a1d47de2a2b547478c2f10d76eb4c79cd21de4d86d5fc08cc1b89d9d46ded6d8c144a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h451da7f201f7891b37f71d870a30cb846fbc73b280faac126782d0ef1527c5400dd9d90f53edeeef39735e51c01f28dcdf07b5795cdb579f75ed4483839ff79a4104eef6202c5f53959e3c1227080eb7617a29232c5718a6e11c586a564bf0a7de0cee3d49559acc970b5f33ce940e2e15484ff5cfd7fbb2bc98ba18a61ff93bd1c2a5e9323b86e5c2bebae17ed8a4a02beab893049b22298618f1e9131a96ab21adf662eafb62657bf4e24be835ca961a403adb4b2fc5a846cdb07cd00d013b59392144f8357df5b754344bfab70e50cd716d885af9f8450050a49382faeff85c165dd1e50f95426323463174788ce6ef46a5028234f3afc76c38f8a70535ca4bb62ff5483f694c5891187d08b1a5a3affb1b4a79e96c4ba1326cbe4bbf388fe4b80b0a37f1d5c55aadb5a138b9600f71670fcf8f63f8efca4e74d3b5f3d3a18773cca60774b19c6950d551df269e2638ca199cb15dd9bf0c8dd69289aaf51df0aa10c93e2250cbac022473625926f3a420c3b323fe62b3b02d0906f42bfa6b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha378952a2389194dfb598ffc55a07d6b6703f54ca69ac44e67128d83d12222d4346afa50b9a0908c7598ce55f5e9e64efd8d86f496c426fae4bd72d377253853409bdec05fdc1da16aeb8f0f24f7ca472d72f5af6079f09d7d325997e6090fff833c370104fabebad2bf927a0cfd30394fdd1f1386364bc737204e2f588e699fd1d203d0624c05536c078844dc4da09ba677db193afafe8a098da1f2a54bdb3776bbe5e0201c551af07dfad942ab284ce3a9e30bfc10b9efe651bb168930b0ff8442016572c9a82acfe6e73752ca45eee18ae8124aa3da0965598cfd863ec575bd21614caa32aaf3a8a16610d1a2099752314f983cef7630b36684290094eee0182a3b6351c48da00f5f6aa7cce32afef7a4813b476be7b415c2392e342e8f36b3deff84d82cc59af868e69cf460aab1ff581db173777c3b0ee62fcaacdd443434b2520ac56510a03394e6c72399c1640b794111ff8cac32d167359d134e86c25c7294900b9985aa1cc88600121955e21b75ff1e90d87c4cc00208d18ae375b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hdd35f819548ca648e8045d88ce68b0ab39d4e0bbb7d525c8c512868d429333d5e2c2ade934647901507294862ea07cdb42d7780f11b40c8c033cfd37e0220df3b38d9e7c9e99b64b1e4b72a5aa2964127dd9c51f065a3cb9eca44c0f93a1fd1b3c461f62c30095cfbaef6ce6ac886f10a36073a3063605badfb8a32f0a5ac5ab1ec0e969350ce0fa9617175a2b05937398f8acff82d75e0a1fbcaef6c3c99862ef23cce9c0be5d77eff9ef3010d9ebff8f5bb86d060a270854c32f47074af9cc768411fb3d45fa5204b3920574579b1653a601fef8e5804fcb0d3d8d04b3a53d6a080ade5811cc75a4631c49d10eb9114f54062660b3e39668aaecc2c3c75565bae80bbdbb89f3f20fd7af035614100a46728c1c5f58123fd9161c51e30f894bc1ca39a304c7975edf81797a4b79031efa8071a71fa7261fb9023855619c9196b13b1775587459b81e3332f1d201f1cd054709b9957125814866bb31d28ac702bd4f3fe438d3b8d148fb4410162ca1c5c8096bd273ed246f3eedeb3809f5461b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h57ee30bbc570871608548a255719dcb9dab007b51e99a18ab0cc3d022bcd8bf936eab9d586b33bc13de52cde70a0638d97eee8d96c810b353b5229ea311098599aa041189cebf348c2c674c626831137891068be03da417fc6f4f9ef9194db1c8928b80b0d12cd1af05473c72b29e6c4fb039007f4db1016d7117308723e17ad4e02a8f3976fa560b0f6953c6ec5fb73ed958710484413163df7192cbb5cc7c298caffd7b980be1eb4a3c195d96a05398bc034c3cabfc1cb8ed9a3fdb9eccbf5fc01588373f41e445ae8d62031634c5960a4297c384e754a1f602ef89888e9f232e74cef6e5e8cae6a7ffb8dff9b72f708e7edebcd22d93f8e1ac94acf822799cc539aae2c92dec5d0cd0466cf0b9f508989addfe14c608488b889e1b149848b7bcd293157e147bb1204fa8ad89f7cbd56eaeefbd09d15ab55a876bdbde05fa95fe9c86d6b956058d4e217e97060ab306bf2fafad5d890cdeca99c9912ee2f6fae9c61ef384d68bf49b8080ea3ddc67105262fe796cc74332ef8f4b9cca8160a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h60c8d819803463acb9a0651b00a7a8cb25005ea194f35f40e96105454871f0dfc7413c008ba507c7457a43148086ebfe82f102a3735b19907f420bab8d302e36b649142dc87c7049de870865fe452aa3d8188b0cf2a91d7dd85b6b46d5d2a0b6c5bc44f472078cfd5bec2f01a351bba9aec3a6aa5bf7d5319c685a5cf1c4d44c6d22fef52a48296609ba4d0f84b655d5b4eaec665a75e29bda052e9d9cb7471b718f097d43bf43442cc73dade3dac2c5371078b94562dfa6a96a672317ef8ac604fd3368b31035cd4afef0e2a179cac42412e72c9a0c3e7a9a929541108b2af390d581657c35efd04d38287ad20a2e662fc5f5935b3db1b97549416804963677ebe88b1029d56729b0806fc42932cfdc8942b138a81bf0fa87c56ff9f331db5869909c1c01b30f9170e701c765db6759e0ab6a68bcd88dcd6a25a4b5426a0a62079ebf5d5fa6513f5639ae0791fdea0ce1224ddb736dcf04df4f56f79ffd6e63bfa81a51d8daffece907acbbd886b07e9114e4bf2d096397690f03408a672a89;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4af0ba1a568c8b55e8cb08764ab9937f4a3ac32935e57e7630829bc4c958b28451c090be9bb5f55e640cf966efbf1812154f19e5dfd6b1114c45cff638b1deeb84497cf42db981f86eace3b1feeeca43f9ed03693d70133215f0118ad42c50af5d6e7881543a4003c9324b26c54ac930815084d34d684042dee77f24d4e3b76b958e53275f2a6fe07c19e8c08d5cf67edb6083631883b499becec9f5b379ca434eca09d5fab63791fd55abdbf5259361c984a94cda654ab198ce126adfa443413972c780ac0bc5a6dcd80f75067597f6bafd292bdd1254a12302a92181ed1f45a01f4d80433c3686faf02cdfe0b545672bd0414f3e4bd98f623c7c058c8eecbcf3ec0ebc7db02d5ffa75b1db2f4889a8dcdf5c4271afd4144a11265dba13bbd3587bf65d690368c328d990802671f188bb1d982f11bba81a34eb1598b63eacd10bcbc179c3cd74a04894c1cba8a616189a652c1ac852e0a46f481cbbe404d559d543a308e6d1f4f090b5efdab4560280e7d0ac629aeea2122db86e3709a75e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hfd17036886dcf5b13cd5c450870d3c8d6d064a8d61b7c761ab46ceaf65d287b705b8c8397521b227df6f8ece85bb82fc3d0e9d8b4ce67cc1741f1927d4a3a04b6dd1b878970678d86762267ffd4e907c1549774c6e97f0b2c67e736ccf97acbad14493a3ef0fedf503c4125d6047f727a2c3c8c007317d41433b47eb3e5184b23e6e2ba18a84c3a6767f14f48ff5a1c28b18685b726658e36ed9df20de9173d3164ef1f2e03e20df158eb024ff8c744a3245794745faceb30c3dd3f980c3c96e275124e94584ad9198eb0d2eb21e6bb4cdfb8331d42f7a30ab697373912c9bc32e0a2811fa6652f44bce4f4441cfc25da37cdf6d965534ddf6e346f01871cb952d8afa9a439367b7d8f378cf08a02c8c13120805dc3c29860c802e3e64aeb793cf0899cf6bb3dcc5284bade06756dfd6e721f3360c1cd8a0eb30728c7ee4dbe9f64f24171ff1632f70dab192c2e37399d3fd2f7ef16433208e71cd8276a092063f746d454f0ca4562387eb73cbac37e31db2c63749d22dba856fb55451923b7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hca06c325143d100380742b1368d17e112800c004b169d1e5215d22ac607b0839243f71c0e07b12fd46a6dcd4f4945e47f1fdc4a76ed534da56988c361b542b9e86705627f061bbbb0db215336a1e6c56a0a9f7087693389de17127f5a3525aa4c66f06259287f12d1f147793137979884be8a3c31cc84f941b7acfe54a092ae2aee52393debb69b28be2da610344965975c96ac9ae67f6ef9dc216fefc5a19764bb9531ae9df369a9c150d390710247e542b220a561c9b345eef58f6e6342e91513c91c6b6bc79cb978e69755825b9fc9dfd72edd62d22e20b037dff66ba7077761055142977f28868be9e672430b0664e4e85ea2a3301da6c634d312b9603794c2b7a776eaa4e335180be1ecb5f11115faea8e09b9c2dd4bdfb9556abbf08e5deffa56215ad43a08ae6cb4412cab24f2db2eb5ad53ffcecfdc816159c6f21ebb1eae8c420322743be39462f2a9ec336e94bf6699430de5a3969403a4e086580f529c6cea6a7912d24cdcb2c8e7654fa3ce8e608a5adc1192e89c843c658dd30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h85117a33e24efc2aa3a1fdd5024ed5c53ea6a9779b24f834a517c8a4416ea7fc420a9dd2085bd82a7e959978c534e1095dfd97aa2332f04726776a83f029299c4ab80077ec019571be0c51f4072b9eafebf66e1bca64b075a0e13be5a6c31239a731e898cd200bbba4318d084b209a45639650433ec09e07f880f835135a25dcda0fbcdf190d6395ddc601e9df050ff5babf1027c90e6a0be2ae1cc2a0e1380e9c6beab70216336cbb48cb60a0a5d427227d6bcdb2c3768f599686af1252c08e86ba99209e9b31f550fbd21fb6116e1269b939fb88b85585715e8e5356231339ee0875f899b972a9baa4b1129108f94602efb112008f19bed38697d03ee89c7168b93ba9c711e9b9b852cea98b905228758a9caf9460a693e94b91548f1c278e1072861e46508f85d240f18506ae6a4eac611176ca7bb929ef74ce0ab05a123660f57674d8b3786dcd1a272e86c309701df2bd0b5f7d27ecebc1fa42b2f4801ff56fc81100e8564ba21a4996ef78d89f2efb418ff96babcd375014606c493ef5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9994996c553c5398c1d0226c27dbecfaaa8e78631966b8623e8d56549e92cabb164d65ba3dcf61214ee0e3cfe207a5dc3ca344eea32767364540502d54edc3530cb3ba66e682f0e5aa9bb121ca6d80b81cde9e65f5f1e0de453d37bfa0b440c81e821cdb244000e3ecba51c54dd041f076b1c6846a9beb8b029c4ab8b1cf1a322c43517e3893826ccde65321b72b2b6038239dcfbd5992293ca3c91744e6f039cf0cb6aaa76788e96ecda3fe31d7924a2c43abd5c56934e61c21157f9352b6770e06e9ea2ef140a972bf7698571a5049fd1cb072ad3c896e1db5f167be577e65b0ed0a86babd9aa8029559533d3a0491a631ee1b3ce61399ccf42f84bd33fb3885b69ecea17ea49e0415d8b4981a8c127d1cfb5e249ab43c5529b2efe76b53eebb94df9a954ffa3795a17f9097b7d1699e1285253b284d6dbd91e1e68edc65da7f0479356ad7512760971209fd27621df4637d4e8fc0f7f97f99efaf4ce7eb8db16061e8e9c4fc03beb02bb54a2875a6504e391049a2e7052da5907dbf330fb1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf82ce554b93ee67354442ed41395703474aad34a27defa3594c65222f490b4cef9b3bf39d722a9f126450aac080cb92d7c64cdb924565e193389ffc178864383c233deed3b70d8a728bb89527f1e69860e7a4cc5e66293f12a516c19362e7363848c84b53a45cb195303b217efcbb9895bdb74e8e258be08bc274f283ddbf6f30f51923d9754477d2801b54cfeb6cf1e32245da167a94be0b3953cafeb953db227f00bc61cccfc700e8eca2ede85c8d280f694966dfc6e5a01d4cb3eecdbf7c4e72509abf3ff5e410a5f936b19459983d95266c25d8cf0f213dd183f0e7e566335ec13dfc13838cecae68881f87298dc03d3e6d33bb6b767da793cfec2c6ddc6780fc806bbaee0f0d186d383bdd2ae37722562420c92f8f181283c4c703a835d1374ad0df387f7e01f56244a066d71a9cb0c015767ecf3bf512377701f6510f34ada1b0047c7436c3badad804483d30f052e5c64a7e19c278a16520fa808d465596b1e7ae596801322432736ad11852782b77173401476698de0b604198f8398;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3d96e3e265e092c3819b6011dcb6ee04a3eb307b07234eb0645025577c581bd6df30f0db3f86e0b45f295b0c70872866e78b8dae1739ecbd1cc85f24f1d7780b5e5c8928f2bd78b537f9a329a7e927b2500c94e1d5b7afbde32ad3565d69dce1c5b67790d32635c1178d29c9e70792792f8785b5b7b6287c2f517b5c5ddec384d2eb20caec208846d9323268f75b0711a3be13a8f85eefb93a80bebfc02acfb90cbcbd644eec63e777f12ea80296e19130c3bb65f14865e0929d5e3731e23891501e9920f010fc3d0053fa21f01bc91ac4b907d97a9d03073e4f721f248ddefb78617dafe3c2c0978c4f5ead9d393a4a961f5ce7f7010605abfa4fbcd53cd036d00ba71a13c0cb5de06742ee4143c8905d569daeb28155eaee89526d132a70eb01e0710e29bc1c47c27281c1d1b3310e56337bb84f280822b39c6fd7a07e5e242fc46916ee93c434dbbab8d21a58a3b01c6113939e2658f4eba417306660ca0a52a6e94fa69cf95c1dfe31c5a13412e90b06f24377cb2a59f9458476357bd120;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hfdd78fb89ec2a1523a0ab8e389d7c41d0b798214f5e87e6bc8b27958962bb679d7c42c98575cca3e81be10aa756157c625dd0cecf9c5dc509fdce90e83fec8fe22d953e6569dd1352ba14996327e630f952b4cf281a8841efb7ebbe57231cee0b9174b8b2dbe32fcd260ebcdb90608e2f2f6348b6e9a3e9ae21021397e7015ad49e666e9954b6600205d21252f082eed65992229e555235cfdca4750d806935d5ec18d61c7170f3a69de624dc510d042d620b8837be687e8db627af061ca87d25ba1c8a16ce204e8a119aae92fb50c06616e35824eafefbba0e7f088b7166e24141e75108047a9174e07e9703a824294f0f6e296cd437ed44096913de1f80cad5dabb020e7fd889a3e28ff53804a2842ab5d5d811cf681b9cdca556dae6d54e6aab008d439dcc3c4212f854182a9ea0ee33148da9765c13e220f436089ae0db970e37cc45d92de5034d5f4a7938e7a30900e58db9a7000daedc099b9b63af3b2b10ca790c39dcd55fb5150bd17f20ee04e74d3e8adc3cfbe81da920daf6aa678;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h11642821a0a8615977388c1da123c88f3f89409cc4eb828a1335b5f0922a9845caa371c638d93ea9e41c87c08d595a4a0ad97db9a9d382bbd89eb72be830b763f03c151c3aa4a6b838fe2a5f7f2a5e413edc17750dfefda7c2f186aa68fbb07737239b23da7fd6d71f67fabe503252291c9955ba2badbabdca2b46768b66b8a6936658d1108b576bf33c7778537ae3bec65331869fa9f61f52a9dff3cad80c1f9d7657128acbba361ef5f71e9eef561b4ad8f43c223af48edf227a72f853c03163531a060db1499f38aae97f696336ca20114a8910f09055269050ac3136bb40668bc64e1bddd551811e6432786011121a6bebf47193bb43374301f01d1794d989114bb1eaeb3f04df35dfd9421d7a9ea589e371f95110757bfc7f3d36809db5c8f93270f1e56c22b80c036914f0457eb48e4fa1a088835bf59ee5a7939defe36fcbb8f999a86e7e423f6f7473ec454515b2a6d2cc67902a4fc77c5654ed56b14af487830aa7e3b018d54a974eddc60ac509ee113101e0ed1bf0c48eca1ae6c4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h80033a982ffe786722f1c84a6a640ee09e2019a36873b0f73926a438c9970fdf042b8c0dbd6d4723929b36011669c9ca870b71db4b80a4df9cd40de88f976a6023096cbb578723cfb18e85979554c1d3b4a64a59c7cc6ae7f5127d73e205253541e095fe1f9d3643c75dbb9e025e6efcb3af448861de8ec5a53502cb5829afc90effb0b3dfcb4e9abcd84b24f408ae01c4bc771de07e9e1cfdefb518ccc1e84d4cf75766755b6963286b64bb3afd0cdfa448c82fa1e5ed9411fecb6878c222aa9ea9c54ea4eca5c5afe908d2b9d82ec0a7805c6c03ad328f747626a03d1ee6eff3600dba41f1e78b56bf928555442060c6106e8f67e27cfd3f097330320854ce8feb54d69a5040689f45479e707c8355161d852e103ceed28bcb48c062ddb14629bc0e2ae4620d894af720831d4ffb3f49cf041bd6eeafec981ee119fa350b084b74fc27ddfc261d75988d1abd72d08362037ceb061a75a02f841dd8facb6992e3205861baca0503f43fdd16261c6b77721babf42910c615ed40ddd042da4a55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h25b62656c37271b8700a6c9a6c289249ec4df4bc3ed5a7f4726b637ffadde4d5eb38392f93572aa61acbad361dc35a850471b1aeda5ad9f1efa1738633b021bb2eeaa2e03cc7011e02c34319f5979bb24dc1396faade77c110cb2d95a2b90e8c5977f07f171794e696044ec716902acd3878f29943e2ce2d5a10233a81de41bfdd5eb49d80b6fae2a159f99ed2a8988d084812762907e3563b5aaf6661eec12a56a8dde02d83d03c4d0315b14b6e9398335194547d2e4d451f12f538e8a1ded88d5bedb1ed6b933cdcf83dac9fed9be3c63459f1f5acc91433f30803d85476aff78b7c696d0179cd6bce024ad04bfedd6c026183a79386bf00422ee852231b04d24280bcba99c47c522dc0a3f997654c483b891346188d409c90cbe788fbb88c948f3f21f23b19f3be05c80c37178508fe5058b2d8fecde8d7a3ced580c65525d1ab6c0441eae05234ced1afcfeb7a334b297ad53d85b52696f09365258c084a6dd13928340bee27059f0d6564c8218b7a49d42dbfe9e99abb0041aafa32413a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha458fa85c60f64d08599f32072237e99edd3321d079bbbac80e19cb25521e7a88db57cbc8cefc5526dc53c12248d2be3a5873d9ddff259bdc9aaa66620e1ee6d9a31b0d47fa2f1d2da44922ab9d250e9c39c1fab5142d369453be4ebab6ec0329c6c90ef7c649640de0d99f246648f86879d707ab6212ef5e8d0f98061eb8975021d4cbdbc7b195bdc0b80b21fe2ee9206caa271bfac245f8dac7edb953b92857d2cc5a26bea3224ab17481b1f14136fb1812fb1ad469e535f3cf3f4ffc8ff108626069b1fbaadf329d05e021363d28fea5460947e9c2de297cf06eac624a8f588457ce572110d7c05f401ce1b0f607efbe718fba906f3ba5d7ad6bd25b9543e369f140469a60d4860676942f696109e844cf1cd08916b0f415beffc7366681ae42e408d467fbec4828c2065f9f4c9308c2ff91f9cd712445ce2b609775c545cd67691e5a9c600d4d9df14f9b497b88575575c66bbb07723992d6176ba1a4ac0a86c4568eec1a386d459a0abc10cdcc42ab14aa2b309d290f9f80e7eb75654e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h75a068c25ad07617aed3149eb3b6e0015321b82bf559c927d8a5cc8d41f80ace2a23cb1100f2e1a9bfd801d23b43767fb1350ec2228489a04e5115925f20e4e1093c25bd144604af5eadb94d4146cd1c5d654fe0a0a202a75baaae67269306895300a7d125270358c2edb8adf7ca9a13d64ab06aefe37e3352b84bde09b924c59a2cef51be5257d786210e11c06efa5c8d1160f9473a1f2e5c84c7ad46b73bc730831cf443644a17bc4f3cad0c35863b4c28c70df1e9b59e0cc7f5bdc04ba435d9d0a1cef7465dc2b1f3cb52009d1a5f427a6c2ebfa2458c00a0661f5d4c80dde6536e098bf992fbe41f34aa4962d57927b845959f832973bcb4927e648e5baa4dd19df2d7ce4323617c61e57a68c25fe050e4ff0917735422930c7d0b1759ae554aef1b03c21d03724e4b2842c5cbc5a442417e9ca38775da6da5a11799d8872817b5712a6989f5784b9218b2f491fbe4751a99b21e2e6fad7b962ef208e6b12020f0624bf1a3bffc6c8c4452da95c1eaef2a5b98c580e9ab2f2be40b7864b8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he7a669db89bd2992ff30c7c120760fbebdcb64d407ba2a9084f45d89b5948aedbf76875d9872036875f7a55a425b56e0aceb8e8eca6d54323c9a78eb3ebc190ac306681e9512ef4ecb77c3eb58b05147ff7c35490a6b0a2d6574ea618cc290ab5bf29066ba52b31ba542bb37df5ec32cf107d67dee3eb514054ed739ed5430ae361fc53373ff405a052c1fef83e0b3ff53f5ee9c09717baeb17180d7642fdae3e0bcfed0521ed8359365a095ec5a4461390af0b0f4013c57064449a18a8dd0996cfd363bf6a6295bbf8d7a8eeda0d832c5525f1d32d901e2b6ba6366f9b9b3715350276b0257d9b77dc8e19316ebe0193434b59e857e1787324533956e925da3deb74e9564242c3e9024117a84db3060049339392ea5dd2525e904fcda6062e7b6a0b0c14a1e097d0a25601e8a142506871aeb536203433d79956398b823d5936c28d4fb3fae1fb8bd1f6700648d824d866f53136b7f5ba1851c416d581a0f5e7c2bf86f7b2935f6b586ac2b50e7e476bd1522ecf368c5fc8af02c05fc97ef6f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he71608877f099e5e9da7840f77d8de9e273758b8c7e20c446ae4c2607fca27be35480c5306f07170bc8a8a59b5902fe120259be8e8c738f7b6cbd35534c8c033091fa6b3cbc467809b5e312ac236b60cc7e69fc04cb2a3d1e41352ddd94f83b39f553f1a42ee0c4edbaa169d36961df87f2156f347c89d1e51ae66fceaa51b59c4333e8c673f9e3afc4c2e2a6f7d8c983005f2a6b49fb07fcd09cdfe3a39f3191bc4b8567d52e3c4935bd7f1fec964e8beba98f0c97ed5c7746a5b1c775a8340e39d652f078d1a6c1ecf8cc1e914a05282244f8e5459cf404aec59b8561aa330ef96b9959cddfbb11dda2ac296331e59b42ae3f93803cd0c60b2a11e5fc989a0d446e7f84378d841317fb3e6f5bc03abb9bfdb89e1736fbb15e0fff25c1f3d7cd634af2163f06bfed58832bc68a031449af26b8b2375e156da82e8349c1d37f44d9517d49e2e02ae58a698e23b34093c5470c154d5997830f14b709c815276115241ea4e2850e4b1ae42404613295f232748a3b3842417034a2265403f696cc6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'haf6a3d42b77782b5788bc96621a3b0cf2abc498dcd2ccb8d234158a921f2229102e699acc0d165e981a9bb89e06f8e68f9bad9197ff623cacada15d3cf19d017846346f973922f739bac5a7b5003aaddf2fa7d3e3a5d0b40c3baebfe59ebcae19862316966825b38337cfc59d3c0e680e3e562b87279dcf413ff1c3c323def4717ac47492b692168fb4c4fa63dd984bb90c8dac81b1fba210001c994956921263859655bd1bdd0c5eac0966b0c7d6a7a0c256603f616e20941f0fd111905d49afe238d887c12fc31fb628f3d5e86315662cad80ab08a2723c6feaa003e501581b7aa68222983ec699c5f8e4311e12ac61a75e3c3c1b7c1401fbed527935b7d442e1a0204a65f4cdae759a0509528d153f5a78216f1ebcc3e13e010b24b1bd6259ce58f94eb5d643df9b9ba94ab5daa0aeacbfa80b3d539671914ac9b67a094dc1ada70b145feae6d4eb953f235e225e7fe134a9176056f1c4996434f3a8dfddcdf8d801c0b4536b0c8e638ba3f7984f691bd0a2880523fc4367fe72d8992e43e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc83afd8410675b6bbe3f2a69ed6081e28abb85ed520fdff0ed91014d23ca7fca4e36d2fa48365af16068e10d9116af489654045f69a037f984b3da9401253e5c13c478f257a8efb0dfe24b5dafa2d78b8a54cc04cf311d1d4ea42b48fa297f31872cabe54a64d90292dbc982082c751fd19a9c0a19e9d65f7b285d5be3eeeeb91633e66f174a6fa28c35b7c23c6642ae2f21b28202714d651eb77d64f8759320721e8a9ef1a2cb94b14e0f37dfa1dfee24d7d2aed9cadbf670eb0b5ff8b8aee8ecacd7e6f0e414002cc04be90e42c4d5c69908981149e71e0c6965d370bcd96854f24889c78e8fa4782d834ec31e91e92f3ce11aa94c9991fc36ca078708d474466d40f21dd2e52fda64aa30b4389573b1078977743d0c1d10d4bb2343dd384f5774944e0da80f7bfa9d8de77190fac543ce961ef99a5b7e70aa83064e28b2ecc3c49c32eec5c62eb6acb8c767616d237423e03347fac7842b6daddb4a6e0c86f024cfe08e358afb4e1a03235508ee621cee4847ba1ece88978cf130f02b029b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h763cd8203cc0d31112beb96b8ae8d11fbad8a87dcd5815691c27ba9b8bd550bbd3281634153ab3b1c9bb518cee192ecabd0d5552aad46bf9cea912b43ebccc0bf20aac590a30f7619a1e1c5ff280ffa2acd83b4edb9ff067175f29045efca7d1380ca14f101ac40ec28f20d2905482e79ecc7ee376c52da4c3a9f9dab79c20490be3c11200e5f22efa6e66be46c1be4c630fa84675777e7ea10a469a84119c906c8eddac0f64805dda3e84ac5e2797ac87b76f8c17cf60dc3120af325e28933db6e18c1949a28578f7fb3fffe700adf8b518c00b3bc42454fb6b625acfa5d8b98087b6333d596abcde136ec95a125d99e59c11104a1ff22fe1cb36466eb1e6f548b005ae900ec45b7bbd8c1ada19c24262121951c88133978f331653cf9824ef0a8e8e0fb3dc86606893de19e9b13efb4de17abd2a8bf12c4b2fdb75b515340bd9190b87909b9fee320b4ee7c2bc0487205314b18cb33b2d6a0b287c0313b0ac9ac1c246207b3dbde37eb3ca7d51a99a7ef0fcae3ffc8d816d7eaaf1930ed3be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he516e9cda82955ad7b26ecff0b7395b0435d14dff73224049d03c11edba7ab1d284c00e1bcb65435ec1036e01b45a071a0d1919fcd19044cadec9d0928071387c4b8a0a2567cf70d33ed4ef8642ff92167ef1c686a99b78cf0833a48ce68e5de4c53c245e5b6c23183d97c06097e75dae9efa5c5462c189aa290aeb133c45ca1aeb9de95ea0d75b06f93c5f64d10db82a02fe9a1d80c1a3211306b78959b3230426db9e186685e272a89959406f9bd603c860ee22b16f53e833168509123b076c542523eb9ee12740a6162ad773325e4f81a6f126a5f33ccec06120c2b52b6f2f9e9e2b7d4a0c8596e09e7f6fc4c38c8bc3722032d24759b1f0f630e4786540a9f4b99e718cc05feb381b11ddbc8b00184ec06a8822478a7bd738eef5570d6c00bd0cfc34acbf141f2bbbd28f16fe657eb2b3062350df88bbaec6dfa093bf284b839cbe4eee1dcef08208bacf7abf9b9fe467bac474c5b20f0e4bead56914cb6ba59695c8866bb0104e5a8ac8f9a5e01b10e4b6b13eb307be134b16006d1444;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd32794d65515bf639ba94dcdba7492dd392c3e7dc88e75dd4c27e60bf62e34b482c46fd9c2784ca446d756d5d2ecb835ac8a250f2c95f74e47248dd7b5516ff27e5fc90e2e41793578e0216da7cd71e7ffc1a47f8bdb37bd1f11094e6ba324baa1c086a244f7bf9828ebba7945001ca5d353c1ac25887e8649f373a1173e955c0cc840bdfd172c4d61a6edb26a539fd3770769d3b0572fcad99c8464f11ac35bfbc75f878d2c9897f6028b585ba02f04448a3ebab6cd2fc3c642907eb9252fa4fbecbde8f037b84d0cefd9cdee55ed5c79cda0a1b1a9fc66f2b588b826ba57cd56c0d40620ad396553421d6ad026800b9eb1a0e3ce06b47c2529a3adf3ec73f731550e0005afbda2d2c2bd2c31b114746df4e2c34dde330d736e8ed97158611992b39c6e7f108a4703936b7ca4a52bf8539f93085e5b2e820be9ac7960c68d4dafe9848dfbb8464ca512bcca12ca61b10dffc0d2713f4df9f85b07c8a3e184fdb6ec9405b274f55af905fd09fe2c8744a71502d2d47370365f4cbce986aa312d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h297167a2ff47d3bb59237ec2ee3ebb69209c8bc78308a60879d0deeb0d1cc37fc04491164114cba6163d2eb47f575d96c706a6f27d22859930b8f76f34aada3e956080dbc235c92536fc423410e9ab89d03f44454c1e6528aac94dd33326dddd305131120206bc50814e6c4f5efe47049215f0323b2c636314b84a4b4750094ca2014dd6dd6bb47f0bb633a0d193d7892f229694c05969ffc47e489eb38b27f29699e8369d0c032aecf111fd25f2fec27c6fe8d202ff17ef75e0683656690acf76f7b0f98138ba72dce1cbcdea886a72bd4a5f84eec845a92fa214d965b3591df15f90271d4440639e77cc3e1bdc99895e59e37a45fe4146f176af572f7e2eb0580b45d18506bac9323879b9f94111ecc8622a28ed8fe937f70c0b02164895895562133c2c76121a56279e8048892cff821eb82687e17c90215db2dd18629c4f62d3a5287858da22d219560bc9158357d48f9ff651a628303fcd7962dd14af8f4bcba22a65e88c5c4e2b287f218a1b868d6f3b5518a83ecf862adf3eae967e9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h90d50725450d12b2554dbfb64da9160574aee3ba61ef45a7169f193831b40b713cc4e61e523a8bd244b3c92324e6604306a7cd31c384c4f20f02a04aa346a2913c400f42a2bcd631a6da1d51443273aed30e68a834be7bc9a88502fcc33e0191da0771bf6ab0c4e27f67c264235b448e7763f00bd8549b7c6ca775748330021441992723b2760e91e682c3959e34e473b77e08c45d112a18a1c392a59daccc88e387bc7dbd26763da3844de060eb8c319324e32eb6715ee48acda3fb2e5c5adefa61710d44333a3d445bac191ae75932903031ad9881b76c4ae9e94a13b4def5d4428d4717134e5a2b5f475c8b47dbfccb1b8a30b01676064c84dd3261e33710f3e63bdc6c2d7ed4263b9df53526c632bf2c890dfd9e93ef83a5aec43c4c9cd336d07dddabffd5858feb826931d9ff76bd534801b923d726e2cdd8124d7b47efdea2d72139c856c63ac03c71aee4bf3f1d19cbe4725ee97e89f93f1499f4c0b1c26dc8de54bbb9c2c813b04f93f7084d40413d8eaf69377c4cda852ffe112b8f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9fa9b08ea2af95230aa07e84123417cdbf80a07f21ee00881f9049cd19208119f053f82297e148af79b1fbad891cc04fffd91bf8ac6fae0a85206ba9f0ece8e4b66cfcfacf37cd8b41eced8ac7d2816137385c39edd43bed2b51ff6116e687cd4961733c1a70b5e4e89ac05935b20af2c5e4a8ea5e0c78a240a63942f969d88f4e8d712b78b98d57797daa8dfef80cd1ecd00debd6f7b502a88665ebd4ef8098bb3ad10251cee47f115d320afc074fe560dce746720f3fd845e997b11e2431aa4be3ea879975f393ef69ebb95f97f3d1a55e512a1c6e1156f1b0d34cc6cd3b8c4ada7114ac29e8cb3f9159511cf9c00b0182c0a567b3d9df67fab7feec648dc208a12a4de0596f272b6c8c2aa9efc9ac6b95c9149e3e3ebc331f42daf6825fde5975cac269e96b37388ffbf920c3c3e0efe7dcb07813f0f51d5940bd98814f53c3e027fe9b571a5254041ee3d9652dc0fba7f9fb88eefdc02f74611f783b574a5a995d4d5fef5b6ceb123e559b2b4595e080b3490f61471e4a74849c20c0d245;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h43f71a1fb6806db087df87ffe98d6cb427e47cd421339bee3b173c902f05aa14c895b97143ab7059b34696b79703dc873b9c949980358b46e6cb7f0ae14c7a9db42ccf1db79b2dfd391c0b4d888e50ac8307af3373a1fee289519eca53f518c0fad96e455a36af812d0eaf2bbc3953eebaaaad5d9e4c7548c39b85a0e965d19d65ed76a5095447e23c505147aa221679693c6f4dc9136be8081553322cc4046a1949edf9942c7a96d27495dc35a217e21aceefcf4288cc257b276873161c01181aa1633f7e729cf93a2602e124cc35dac528fbff5d3913394a40fddf85d9ee2bb68a17c0fde32da14dc5afae1cc83c2367c791a3b26196d964b9e4bce7ba87b652277e9c246fcb5c56847b931f5b9e1bf439beb94c9d476e6bc6bd54e6f5d6d2ccf0385790a19ba2e9b39e46dde6dc364c092926f7c7d81fbab05cdd94c2f0bd79827c4e5bf3bfdf1403747eeacbe0d22d8590d7dbf3df0774af093785e9ccc45b5fc9de9fe38733fc4e7910860c5999ef4d350cd087b278bd4bd02c01cd537e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h929a5e5609f0b72dafc8b8756ab2280a3258ed506352271b6c85fff80a12b3ae72e7b95c3c0902bab9c56ec9c2127c159ba51558fd3c6cf5c0774b13161089a552d5c807cac852ea803748dfc8a0f4ec283894bdf52ee8d822a290d6798c7abafc0882d7c5449e1ea60ca30f607e57abc26f511b6d3b164dcc1c4b137afe2ecd9045b08b9d60438ba42f9fc28ada30d39c9a049167af4b9f1b26232edb53c2d5a52ef51ed9938f7d9a1daf330fd8e6e508b60919452cb10217f9134ac447518a38f5db972c0eef76e255fa1b4d5abbe9d05c792e6ec136b378b7313c7ad34f53c346f6012dbe875c53fea9ac166a0fb1d77c4295b7dcba0b53bb113696c0b5944526b0bdc070d127d6bb20cfd9e52f9cc859382053c416ffed75f98704ec8c3a969c5898b45f0c39a7b69da7b461cf1ddf98777344bad66828939538cc8dc11148b17cf4006be3add680f641587bf97fe71aadc6f77609f3366fd9a260ef19b283854ba519602d6f7de35b48d6ab6f3ed1878bb1c63a7ba8160caeef1f802f78;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h73d5786745e92af56b4c0226af10a06177c544730021320648a23eb2234278edad048829566c61875de80a6c06059455585ffb322ea69c88bf977096e191feee00534d3e926891d660228b584f3461ef0ad828ea140e963104f38eb9562b32ccc527ca723d270f43de52103628a965dcd498ed7b6f4645c5b2f7f6d746f219d2f788a270210565b3bc4f4843cac421317c6defb32886f2c27f69024751486c2cb1e06366b98bcb3b2d3ab954997b7ddf2b9b41ec16e0d04e23d85e14f0d5342ccec133d5ee2e152bd4d266a44ee3efa5e2c9a7a74e230e72e42482ef275a7eefff42f9c5d7e132486c205b6fd520821fb80917fa06f20b7376c361bc0bc85b3a8b613ca330a41026e4904ad8064bd33a29a409ee4bf67a0746efb982232ce9d7dcd7261fd86b03b26d37c485b1dcec27e4361a3687643e6975620b6309c2d8dd4a7dd17ec5bf363ea1ee253983ea56e061a91f321d254d3b2449d96c06247c78877e3627691b8604f239d326dc592066721e455c0fdb4dac6e4ab050c2f9ca28;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h31254ccc7515a7468d5a21eb4f6ca8e60063abc9ed3d123756c098a97a4373a91699841f869d41ebd0e50a4204a3e76fa41bcc67b0f2f05376f801c326a8e4549a4b06a8ea2d45efa37d6581d1e1bb269f82ba2e385ea5866a80329466abb87143a73fbf15477ffe4b7490027bddf34d35c6c0b739183e5f1423ce176d2358aca1c9d7b5422f2d9f1264999573bfb7229a8513c6d200d4fdfff28ebc0584070c6b9e7459da4834b3549e735643fd23508fea83b7240fa3c14ece12fa9607de84f894712ac08fddf954c2a1bb2c6c94575a5d6035fc7e9c0850fe77d0a4ddcd2425f8944442f5d1fd5163de626529a50b20b647143900eba576a70113872a7b38cbc775e9961959ca79aac3c5da496fea30c66ec0bb562e4a0d997ce56faa7044c034309f52b9d1d9d0bf716e0af794b29a0fe0317c87d2a1f00257c61e81255ba9b3701b653a6731cbe510e1596e3305431119a940073be5aaa8fd1b75336cbaba88bdc12234c0e6a4026954bfe33c2479addd48e1b32805975d725d05861b54;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9a77e149288c2b50fb626d9568e6738a2e8cc5a743ba30122a526672a1145cd0cc64f4a18c2403954ae87b48bed289ce9d27fc7220032d22b2d5b31c2d9ec8bdd7148eebdc6917296d888c502b9ff2ce0ba8646e1c86416f48fc1fb6fe8af2cf2ce4711f05e46d1af011d6b9b797f753398063fdd390947c3af3fd394cba7510a1feba317be3cad2cbc42c76a5177e566a5efd2c3a7c7c39cabf45f406613120e1997f1b55a6513b19a699d5b0cf4f2f85ef29446b652d8758695724cb3958f611f6514de15aa13b9d5e64d82afa5a70fb95553daf17096fc7c4013910c9a90a45102e9e8d50790e208e7f59ec3d492ac8afb3e1746ed319932a71f44ad2ecbb11bb0293f469e0d1e981ce66791444b6345ce6a16131ae0c7ef160a2fe68d9a4c8274d42e76e443b384940ec923d45100cc8bbef37ea43b30c322a81956e467185582ce997eaa29df67972388fd0870617d9f5c3ce5e9b292a025cd6ee332d0e2e9d3ea563785879b7802f29ccec122d7dca47c00cbeb51dd20765002182fd1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc6267574da485d0c13245ae0a8a2b9a5f3ebc4849e378e8df609c77da160d6afe2df999b3129a5bdbc4b8eb6081062defb0ecf24a1f7f178bb4db99666d206b9a7d3e3fb2d1b4f3a7c291a8ebc35b9143d293471ce269a297b727638970d16f94134f0a0921ec827e94688b2dd8e930b68c79a018abe4a97e9da346b497c6470df5e2dcca9867bd0464677621133c790c37a99d74ca9732493f9ee82d7733b6fc709253e735da42cb90e605ff6544f2ad8becd9db7c3ef91dd9053a6a369ee5d18b2c2d4d49d696039ca760e0b701378230b0745261debb5e46f430f6aa1898583e0c019a2b35ee52f363a88ac8d180db2efe50d1bf21e0f7240cbaba0e95f23ad67c609900e0b58aa324936cf1a8b6e7419ad3a809d479790158165f3ae093991b868e1e9b05abdee7a2c7027bd8287fd52e130a6e1327b4caa1e16c56eb19df126d83b7dda2c1e3be20f9dd6e7897b56a544cb51d89a0f840082c8a8836b0e2a98055bd0f6c352db6c3d7cb60fffff1e241b635f03794bd7284de82b287e2d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5e8c46343e3da12945438aaf138e644c4e859a915dfa7faf77fff7c899bc49864121c2171ea63293ff67ffb9df1f24aad223f973718ba327dba1b1359c4c671648d2cbd311c50c5977e042cd6b6354b7d3cf9b98e47e174e2f738334b388a6771a6698e1d54d4e5b3a4ba2c2797ff784d7999990ef9e260ff7b9e9aaaed11d3d5b0a6ef1575e3eaae51fa064861e6372dddbf59a4abc6a93f9c5fbaba196ba3b6bb2e3aeeb5dbd1b24da34ada3b96c0c8b2c69dc63a13c2a19841901d0456c96a684121e3d473783a786f5d865f2861128c313d00e2738e2272d49e6e86f475817e38bbd1e0f4b8645073fcdd480bd4d4a21b7bf0523a066ab33fc8fb9ceee01b68c60ea81fca1a60e971687e82ac324c9f08099964b7a0b130c2d45ae7fc3e484246e3077a36af024feb533b2d27dffee6dca520e14df9958b707ea6b06c7ef3aae55f9b348e82bbdf851abcb066ea38d424105f912bdee2ffb96af6ebf35224daed8cf66f23f65686a9a181fd4ca5d48f9425aa4b0f0ec3041c983e5876ef1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5479b554f5da4b26dd167ef520763ce227182e94ffcbc7f92ce5a0e2464e913ce70cc3667175d09e8b4e61bc05560c46787641d2e60aebdc12a9af6cb8e550c7dd596cb28bd209665c42b403e7e74e49d79fe96ead174bcfe1d2ae8e9825ad4ad25058276185107674ee4f90055b4a40852d28e9b6888fdfcf2323d4b3e5d7b223b0fceaa47fa3114cf38f9629c8e0a51abafcc696dfc02ca8bd59d5fb459ca8d1e46c140658ed47f067655aa4ba11cbc62aa27fb7a4c2942a9da524d8abb0fb3b4a768c4242337137badfda6f8cbf4eadf274b47c99d17d1a2e0beb70da1d449e6db694aded53817b07c1cfa42cd2f0cba6b14fe3a2e65fbedb0d73ea449f7a39469780b24fb31997f5815932396d6de7f37f9372e46512e6363fdbaa009538ec53e93805255017bd2d0eae1c45d9f65864fec5a54d9fcad5a2a814bf72c05cbaa2bcc6d39a3d18469997389559196a4ba173eb60dc1b13901871b6174153d54b1ca58afab8db6476c725026d7f3abf0d3c82a3c2257f638eb368a39cde51fb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc777a6709314db64f1feb7694b29eaf3bc03356f240af71fc632dc91d4c18fe981c9b51ee1886de5165c7022c87be02271261cbb315b82414bb4fec24398d1a257ed0326069764b9546f87979485cd7c96ca0fbc02a0bc148f3a25103a5ec5c2dbe93632bb3063cf1655aae4b6ca6b2377ccb845ffb99329e4c672b38b2a62a32f2a7c52f728e7ffa10215dd20e2210b421d673a8867a66725016fa124f93454e47c0722d974bb35975eccb5c16ed23b51bc25401fe5dda1023dbcca1e9dbcca333e9dedce6a181dae3053d171babc7e33654e1aa0c799d89bd969f8cd2db651af08551ca3a5d5b3ca535997ded2dcceb1b81b4c67506b084d9ce98b0becea9b1713ac28504d345e538270295bf707bd5c485f3466b54f44fe3802fbcb69b337feb6f03b6a9d5a70a92efeb7c0b376811afc234c7a3c3af0b11daebc4eb1f8114fcc1b2bc86ee40dd4c1540b2e8edc3e81a3e21321621e2646377c553efacab0e21b44ec0322b568a093dede89e15554b249fd46305e4a3d49859410afc38c14;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hb9dfc3dee84ea58537f820f5c9976d4c29ba1bade48e4c9685febe1360ddd6cd32c7b98f67f397ba293539106124415cdd797e62e35233cf51dd068b37a39417a9f382423071a94bf47b6b16bf0c517a47af42a8602f21c5373c2d411a1c554abb1a5a2f1f9c6514f3488b22761de4b873776e449b450ec6d62e0f42a66433b70bdbf26a16af45467ea2799e7217e5d27fbf4e00e88cef098f4d533b19b380ef0d8050a6861faf34e7e6fb3273a9d1ae239f2744ccc4ea41ca91314a268046b599ddf1edd3c66eec82fc9d498d8db5de72459f13f1380f6ce40400f38ffac7a533b12582b96739a86dca5f44b2f17b36f974ecc868231337f5b584b1cb856b0ece7752c96efadddd5cc964f165f7f20251561e624088837e4c6936b096f53d22f0469505f5f27953d099efcf013f6738ac9f320635345094c382c9a85918000057808b93c269835e5bbc4c89ee441a5b7457e4dbbc266a2b9ecc564cfd713f57a852e570e5a379d553fff7969400c157f758f6029ed62cfc69b9c651f5f1378a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9a6d2f9a7c2ac54e5bffeb045e09e557390d6601647beec44db38a5111e3e3da90624532d7235e96b8d31d2c184324cb7d03fc4e9560b7330bd15cda662b81447e3f40d29cc3fd147e624340ba7c20be71e49ccaf7149617ad9dc240959f445cb542aa538ac68e5c1a7aa4094ec8ccafbeca61477c32ceb8adec10f4b8286e264fe02f8429c1f14556ee0b2718452206686ff2839c6e8e8297d9026bd478513269e0576729592a52678c605de09cf002f8925db84be45f1a26d5b88d7a4efa0042bf809a847bd0c5b80d54b36b1aa6655f473ebbabc86d53d806f26ce8141ead25ae92680f3d758bff936098981db46ed47fc351851738f2a36050f997d7091233627b496665db5d6f7271716fc5f86fec9918ba8ddf5dbfbc643067a187e9b3ae8892e5a7387b1a02adab4aed37d32eac69e2ae7bfce733257a2bc884951be4815da0ad5323aeb45f357d1806737c5d2c643d9b8e5ef2300df1f72cc239ea3ac5ac4c0d8b9562f95f747761c9485ce39377b23c0688f2c0f21bda439573a98b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h409532e012c46baf8d7e0a73e02f7d5e4671ce481ede3517296a5bf196f25fd57f010d8a688ebcf2d866a04bf153995a6ee61124d593bd731ebec1caa69a577b2ec9041b3613cb3c005a62df5ed0692c79a99a9a87574d4c660f22a487941023bf05423ced21842c4b9dad5c854c6931ec2b4620cd6b9c2da4934317037854d590351f41f37e86ae7786002d14f49b2d66b580b43688eeffce51e98260f6e19e26c034e0d81fde68579ce18e8f903fcd0ac4c2b395354f94d4b1a9286ca07af426e26d506a39d071394bc76874470860b256b6c26d5eaeef27bf03829821a5b7bf17a17ed7911154da8043639ca2f8618c57aeceedc9c9fc570843b87163f4fd3adb0a0b28d8d8153511adb2167a926a1f261b8e12651ff48bdc9e613f6217dc7519b4014fffd041447e7a4c2b83a15136cf85d12f8a4099256d023f527897a8add8b17cfb16d1172d49a02e238dd83b1542a6a66256fed6242e2ffa4f7d831d9b064d227ef4cc4b4f2610f389664a4098d277cd6bfc12d1ca9b8678c5e8aa9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he0eed66d5690f3279b0c364191d4cc2739395474720dd47b41855ed53e761bc0b728ccc79193eb9d85223694bcb491cdb5fce8de48ce0975d59337126dcb659e318b5476c8f7d4cd4c211653fb51aba6db07f07d89396be12a44603bce585c4c6a19bb1aa37790a4eb9187554b0303c7430bd15c719de4ae3e06f09eb299ce28eaf367812cbe6fd1b1f439f32a526f7eb8f6762d2427ed19eee2f830b517ef4a9b3e8c3dd342ebb28fdf1186ca16c3061e332cf4b8174a4b55f73e7301e16f4b31891ac49fae72356d3fb418bb31ff073ecc8a648b2c252d07f040b47019d4b6c0cc23ce1074fdaaa316ed26b6efcd05ef22d2d016ae548da497164bb2660068651973b6d174fe8899eae501a157c8797d5e1a98d82d9788007910a75b6f37432156c9541ddebc7bd47818e1596c8cd45e23fb3d56ab536bd9ba63937fb34fdbbd13a9065c8e6f71909221b13c59442af7517f11fd37a7a7e80125eed07b7b236bef0faa11739a9375202fa52f132cfb6aaf28dbb8907c354819bdd0ff78c09a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h76bcda63102480cfb6c17aa0cca4f5e1f64ac5f8a9f9305aa721ef7f5b8912d706f10751e0bc3e4013990b59a10fa28c2b4797eabeb87d4b57df4f3c0df06f450ec982ce16b51db38e8b9962ed1d1048d7438cdd550c2dbe689ea77ff54cc55527a53252ab1c2e8a13da4d089a37bf5504e95d477a4c709384cc4f616749576b3095d0b9b81bd94da0956a1a3af7fa2949aae1c6f93bd8fc648fedb84d9842c6ee26aa0dfac4e4f8dca1976bee194143b245a1f0ea5d9d7a95d0ffa4c0edd1608572c2590f79b3be4b08abaf1662276064a1670dc649b6232b63abcb68e19f2c390d590ad9820dd6852213ab64d7fb49c4e51fb36f1a297a960ea9ac6a63fd2fe3fffb8b0c1e04560ab392ad0aaada905bcd4c23e38a43c55a04d59641babafd21bd95fd5a179eedc2471eee35b41347d39411974943eba3005467f8d0d2f1dc7f7e29397986b396c85f944ce78a8c1da57a8ebaf8becdbc44f543f5031c79479fdd7b89ca7318a9b0aeeed31d00e72af98559bd8d829eed8a9842af5ac1ec9d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5ccf79422feb67d9ce59f4ddaf93904a5eae8a9aac460a612e0a29dddc222e929cbec6dc706d4eeca8eb68590023817a0605d2d6ce177f01ffdc0b185b38dd5614a6e259959b96d93b96966758b4bc47231f0c31afb33edecb5becfe08899165bc2bbeef53410b56b0b5f8fbef02e2c54a05c6a697e867f271f09fb62170ec9040344435c49ace6aa920692e79e4995ed0f1739dc89bf083234cc720583371dda2cdc68638c6e40e366fcc67f69db10e109ef3a43ac328e07003bb8848f91426fea09de4c1ac362f2b1adb28bc8335fb24e23a2a245d6e42c71c2a3ee21f38bdc3bb7c195b0810cf5dffbda042bd8ccf2068938fb27f86649552352d2610b40e2fc2616037fdbc5fe9bb65bbbdfeb953f1327421ba31455d22926884b447d4c30661dd9beb6ed8a64e91d33e12bc7479a8662ef233647f55bd7ae8c6076464f46090ba19545d423ff1e4077b96c9d13ad791b6d3b307c4afd703d49f7c49ce02965a1d13ea4c7b4dc1858698cd481d4117c75c8999fd58f39c924ab1befb8f58;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4c1c94dff5bd9c8333fb3e941f94b2a40417112307c17eb4f127a0512ef9d14a76b49c3a00f4b94405524995c2222e938bb8744647c1b7a77f3d3bccc7410a637c93aad9149cf8d3d31c848d352e203dcd33172ca033a073b8a04e0b211e90be9a54c4ebae6991ba23898b14eb90e55a12912b06edd5a9b671350829ec94de200b9ad08a1e03c92500bcea92d2b6d745fdccf06a3fa3f60e7c490b110080ba0e96025c5b47daa0faa87b2e931606dd8d02db372b1011daf77496768eef36769d627bc061e5d3ca3520acb1ca3422edf05d4311a865862a2e2cec701aa369db3d73976f187f517b663231fc4bd9d0426675cb7c8e0dd41c4e5839c2fefd6822ee29157fdac7ed4df6820776d2519b27675a56a803d62948891f402fa8eef2a8099dc0358784d1ffab841b5f9631f02469b12408a5982383167302db7af12193bb1fbbf92f384a0a0faaf60fefa575127d8fb86fef138f98804a5655d8a695512276ca6a0bb1fc5c77783a268591241f4c564886ac4f9be0de47761e03366e3ae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hb265aa7856d28aea2b56e72fdfc11820a1350dd67f297273a656c64f6bb7eb9fbe3283a5671108c3532c3a31c145cf8280fa5389888e1d575f1c434642fab9b9baf3f0926f061ac5d0fdca2642346a1115120df594f4590342d205a7ad8b814ad59d56df9a464d2b4506701b979896fbea00ac54b443a2943a33b447775b27ec381a0721e5a13044da8528f41b8995e240bb9c067a4274a3500c1f856d6a2c0cd06416622f2d9487172b0dfe5995e43c9306949208e3447a54b9d0b490b1af25b84c04248447243eeaddbcbd1d759f38898a2fdabe04e9f71bb66076de141f5390df0898d8572f37d8f95b4f95a11a76bd2ec4cd6788c50da4a328c4a59b435c06d7c38cbc0c33b601d2797a38ea27c667d84cdd1decf20b1d8b044b6dac1ac397604d3fd29e1160c68ad6cf77fb88d63891185673e173b81f90b960a50f0ac167362bfb4ebed013428aef8bf2d33c1f02ee71821418b71983957194510f644e991c89a82e9d7153c253c017bf408e8d135c96d6906beb1f2e7e0899be79184c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4aba96143b3f8d648b52aa892524be600b383a9ceb0a57c9228d6db0ea1558d840f29d5257f8d9f461a5a6d4832418da3bc08e5874865c4ea77a2e4a68f15ef99445d731c5ed77de8896b9393ab90b9ca4fd26f48a837047b34e3a40660ff12d2cb1a2debd0c6dd1e7609199df3cc13f2739e1c0eb720320f1e10b62f812e7b54f16430e5b497e58c846c34fc794ab323a7fa32932b20849c0176a7bd482f4d0a43f3a15c03a8a62619f570bc9bb5d0e030e577d796bf0f847884ba1e1b8175a43fd862cf04c0406f3bedac4269b8823ff5ac6c6dcfcc08dcea3aa5696240bab46adf2df3645aca241d69c4b2c7c08cb6e63cd55ffa7e281ee2cb8204492196ec656ae41ce4f58819820f071a7d2bcd9150d66659b13fab671d876b96591b058288a8f01c1fbc529d9e10eefef1df7ad9c4bbccad969696c08ebac36a70be9914b744eb013a1e7cd4a3f9fe3f13b9109a4ea1795454004a2f793b9376a3775916d55e621e0804de62c02c332223c623042bd3b032781425f8dcf6264a0c2a885;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc64437c8907e8789a0573270ba9b7f460fe84337c05cb7c78de973bd8bab8e1c6ac30108073172e298ca042f638433627ee3e5f95001f9c5ad3de0b079c385223c0f9dde9886fb0ab12ef12a21459e56a2c7f537a5cc655d8bdde0dbe60bf92027d088b87dee24325b4d8d12cef353728146827aeb5cb58172337277957e3aa1acc5e5650e842ab89aa16ef7486b5f89d65ff665869c068f86043bf2ae029c6bfaed28110cc78197317a2ba7ac09338f1bc4f78df725be6c02253710be7e98beeda573a7d6f561835d6ea4084c65a5702d32f791737be25982ce8e3d13a7aad3de4fbb0a70b90acfe546f7c950e4516ebf5e38c06b20bb22f762c352b9da1b6a5feebd23490eeceff3e348f3773cae2621cd64ca5c89fdd9e54e0077e62dc93581dda3e61011811c183d443410ea6315301715003d9bf60bfc038c955450d139da6779051f4a3ddc7b7dea64c61646db5fee09d0e68fb1d0537a30a8ac3ac24063935d40f627addcabcf339adc1bae488adf8abad09753b351cb95803df6d2ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hec439fa2830f23fa70ce3d406c2c6b39b53e306dd4229baba4c5449c4707248f31b56302a5d4fb4cdc37ed7d1b54224e2c56fc030be907c9e461ebae5bbb6abe5e6aa89a7a60d441e4763f4af147553dce420b2a30cc713c001160f45eb31e2ae67500302cdc37fed497c57f089095bb21f1d4e552051298aa417f7b6e1c93b20de6ed8ec0a78cf7c60d27c495d53d6f44cc209fb8ba799e1fd95fc5fe6222cb603a6b7ba398c739447e76b30ae7f93312b95561bac07dddf1f2c50d52397118e0ba06ecf6c017301893fb402b9db116ad571579a1f136aa9fc9a51032b5dea0b70357053bb10d09848bec8d7f45b910f4ea1fa77f3eecaac96d5d6c06c0e7d5df319ad4e548403540afd0b86e0891f9a37eebd7a0f55e4fae9fe060d1e4156c2867e862a73946c5898eb7b4bc4fab1cc5ecd0c5b21a260d7e9a9bb24e2a98d49749edf5ff22133e2560719e6e030b7509421798a918a2e7427b2ff1bbc4b52656a376d132dbfa09ddfc009ed9d5f77deaefc0a4d47cf00c7bac2a0bdfc6108;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hde84fcbf16b6d9faed999cf2e62104c3d388fcb72d6b3ff97a3f7d976dacc137c63415d54bbff017c71256e8921c0f9626ef81da086f45a9618ae251d67e8e991eba52a7b5631ac7d47318c3d2093d32b161d85be50a1914d8ef262a44f5a012ee4a4cd10a8b1605645d52e6ce19ade5e80404cb27fe91070d109a4a9052f95d67933d0652a1f489916b237b8baaef3a025e6481732de716b4ebcb136e8886084b56a1410da30f73c66c50cde2d737c8a52f2680efa286c75bd509fc50b591c13a5fcf481e733de6e0c00f9f406e8caec89fb51d6d97ff94d38c758c2c038004c6f7addf6700236f51f0ce68053c51e862705a421b552294815a4c2db770aeff548b05d446cd6613a5491a493b95fb7c0510706a44254470d0c6a6021ed4edbcec435811ab0b46e74b040efe0ccf90c237f7cabf3afb1f1b07ead6a6d0a8d3e84349a568714e69a72e6830109b1c2481e0179633276b67e2c38b061bac7d6299bf11cc6c64846946b720b55556745df2d4c1ad06dd7260ef36213e32416ca6bb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hec2833280aed938c8b2c7b6f42a4561309bdfdfc9472db9b778c8df2cee5551c0ac34b1a4ddec7c15cb044af4358e316d9db49fb5c303b16e856b9a70f871f9a138df25a70643c7edeb1e3555a816901d91fa1547e83833171af2d9f48b7e8dde305eaacb672c84157a1c7335be2f68426a6096efd5cfd397c1d9cfc0138232c50fac08bf87909a8b022d3720c335c8562e5b47e2e3ab5701efe61a63ad8540a5136532a837fca568bda976ae5ad93ac60cf051dd3b8a91eaa7bc624ca2e65774c93a59127301b88ce751f7c8c027f1cdf90cce56e4e212f62f4ba6964069332f826d9ceaefb3d0283ade14d1984e90a9117deaee6a636a1d4af09231d5a2da83ec1e5287e0f8d3c2ead53306596e8cf03011d3983c046ddc4afa02a97bda3920a5823e449e937b6352aef4d5ebb0ce46c473a8a95ffde0e8b821b9e0e9749389a2729df0611e95ff0e6027e6314b7edca657a2bac02e48f4c08fe9285b9b5ad536907cd9e98054d135c1db2ea33478405f8f0be0021a257898a258f31c771c7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc52b3c64cdb5c1cf1741f4194a8eca5230e2062445bc8bf00bccd19bc08c35cb6e87820db6667bdb2b45488b20b49d1d55213929ce8cda27862abebf022e04aca39e24ef3b07e19b7ae184ea3a35850000b949a781c89a1235eceee3b324516fd8f63138cebcc2a98e3b11d1304e7d7e6adfeb536a872a2653e89ef8ab703913d8b6b477ed3259dbe7c32527e03029d31e3b9ee749932167c81709f4b1f1cbc88bacdf6c4a5512710069e3e73aa99f81f710c93315ab811b8754e98545f7f39045aacd2525b47a5dfbcc176295c925f7b2ad3d1b471142f341f9df71c6b39618f7ac46bf5afee94a400380278a2c34dd3e71afc772261142c3b3b2b2b370909dcb62af87419d0956319cb3a313522ba143f352cdc8fabed142deecc97f141863a2ac423d9acbb59a2b10483bfb1658dc21e76a558c459b2cbdeb3ed58b249ad4146556b8a6e9bd4decf577c02cfcf681719fb7c4ad8b7fbb2379f9c1e68881d5713d53757142a1f18111a2ec33658731444f5d658559f4c38b9ec0d5132dd802;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h51878f3dad871d5f1b8a003ed9d73c9e42b8ea8c54c7aaa118ac1f6a474fc0394fda1c85ef59c8b4c0bdbe2313369437b78679b5783452c76e4910266855518e0cbc4228864aee98e7f0c87860c47a5137a621badca88f50dd42f68db8f6f50f23813cd8e3ab1dca00028648bc4b7267e12e9c36de241d13ef5dd2eae048e85072975d28830036bbdcd6400a3e20a1067e83b85720485a19f5eb94dae0c8bfb2a6f451b7c4cf81208738316b26b1be547b17ba051ae37ba3745b5fde07d038c9673c671e74cdf070e1dc1d90db0cc225690f26833c68c6244a908ff11c92ab2f7e7bf5731edc51e3ac7459fe84bfe84e3f1cc95532748236424726f34435cbd90c37173f3e9fbade1f619f10db2ae7dbe4b4cdb75b754b86da33c8bd4899a5336b5d74671d0578f04b09a6a4da51817de0c56e50dedcc17271dfb3f1a0fbed6170aa151dad3436f0d86551e668e629c38a0b7aa8cd8024fe75a663cc97f0116b9a8993f4daf531e01e43c3bbae7a603edfee01bc6d4d492bd41ba8485cacd1f3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3ee1dd8a891d2643fe5d732d489899b5f040237ab3f8e97b4c21118a35e50c8d0a2dbfd5a33998f5e50145ce73013a9fad05fdc23d749ae08bbfd219b7a4b325f24bc0bac60565d3c244d5341ed849d76ce4b6d2ebfeae367a0df4bf8993210d76857b5ec41ac4d82b68dc3beb6c5000fdfa0de7e08915f2e42a854a33168adaeca2f07426f81387cf2145a563085c02e1a2175a64c1c6ee6af2553e8a9e6bf1ec8bc468a685547751042f3acdd19c7ee93601d6205a0b86b7b667085be14a225ee759cb3d25ea3aeaf63b96b823779bbdedfd8126d657ad1810ddc8315de056b49709c7e4ee40dbd9f8ef386e66b657baf61a49dab32d1040e82a35553170fd6c3aa2a8c37a813f7bf7e68651323d6b2e7be50a21a7f9b956a14a89a2759616bf7e54333a10de169cf681759e2620843b4bcc88d8ebd20b09809c2985f65dff2214f22693ecac78148b153c1a3b34c1ef62c72cd96360a919230eef51dad3f4c2d19e0f0f9e69427a16ebd940dcb41670c8ee8746aab566057bdf597a400ca5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hfe2252a69429294a66abe8bf1d638be69607968df7ba333c2c73635cb9ba622f47abeb3fed18ada4369c26c4cce7a65b39ce45a8a97bd155d101c4ed944886b228bcba4d417b86599cff40f0b65d5e1a97ea7ab1020d898e070e5542dd9857d538780f51c7bf8d05f9f751653806075808a39a8a8765cf40ea244ed39125b193d4a9d737190008cbd4447f96f2c2bbb2b6100d48f7f3e2995620bc4076b91a6475cbeb19eabba47eec06590a45190ba0b7f65eed0a0474927ddbad32cec1216b29b4f2e29bec5697ff51ecc09ddccac592c32eb09c9b5e51c577194c16641f44d52dd04db7873e51aa91adca8fc54af36bf78b45f6c5488a8b5dc80ae0e7054e51e15ad4c1f0516c1f2ccc481f6502e0b0558502fa9709d3aa2e552eb924b15b703cb9735801b220333dba775ecff58dd61e01aca4b9bc75bab5a23154582257e16ec8f00b9cfdaf94eb7ad37aa6ff227d051ae5d3ef4f027444505c67bcbeabeeaea39f45e872ff2da22b78cd4edef5c5a6f426dff7adac2dc832b219727c00;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h72812c2c48bed8e6ef7043fd7098b3d70cf63a7d8cf387aa2b0eb1907e2c7dd4adba1382ae335d1257ac2f6545a798efa805467da2e3db93ae8c0a77d74a68f523f61f3799123954df82c365cd5915a3dafb9d20d507c959c93764e964834c8cc8546ed95ad90876abdf8e015dcda16dbf5669a66ff12890c6df8eb5692623bcf942f26d78d9f1db0951d9a2a0a80a40be5540b9422853d8722474883975091568f14ab4e3c7a6a077080f2fd8b4a0bfc7905a6fe1ba3e0f3b570d88848030e14b45896e70d24ae2f876a913902c22f181714d63b8eacbe9511818649109c9a012354ad104b06ce30106cfa693dec56c0b5c0a7b623c134c79c914768e27521193e56f18e014d039206b82395afe922445b08cb04b8e229d62dab14c5eb2d137a417c735b6cde90c1b1ed33716681b7f826fae642d03c00a205b12de9502c870818a77d7dd02f989fa5c408ac5583d161ee9c109dc92926cac2f6a1848c6a66bf64dcc0065596255407275ad0f48b3cd7bf7f6106241f52448c9bce080cc97ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hee25fe69db981d1c2c401b17c5f29df40362ba7539d74ec6b9b066029266694bffd2fa14aba520b74261373ef5449bbc98f97b21dbd09856a6da38649e98a091a5aec8be7ed6f18231ab13f6c8051f7b437d897683cfe16cd0c0d07598e3f66d0e25c5c06e13895e8c8f37729fdab14dfd0513db9107094cfa97dc57036adfc9e623c118fb606336ce70812a5e9b9e559c46ce3f60d418f41fa2537217f3005897bdc54e7eb5249a6c9c84b74cbfb1372c23fc225b58c2900e75379d884009267e7f098c995d5610c7f0aa2727ebad0d59bcdbb94d8545a64c89903c65f33221fe1311e6f5ac8be463a1166966af4151df460d5895aa722b793e18f390068b39830ec33d2a75fa2c690adbb72804bb290feb99361bdf7acb1bfe239b284c073b11725bd35ba91a90316fe7f58c6fb1c683b5edc1541528164c8c3c42ed61d2aa653101ca93aca86d84ed0e9ce13bda17cf74ab1153e303b9730eed334fc5e1f9e9bf9be30d5ab90bc2f203bb5bb125afae6a4892e9cd35a9c08078a50d6c51f4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd8df4eb0b57c9930f9beae0f0306d522541579b1580fbfcc7cccc53fe7095b045ebf3b07b122195bb7e6c66b311eb3794d9fcefe13cbe0b044a41fe4c8d3785ad7ef5354252b4765240b2762585439ebdbd85e515d3ef7d7a51f46f99d3fe6b84a15910f6eaf7c4aa21e6783378ba01d8c2bc9a316d0ba38d2a308f9ee4effd287656e78660ca0628fbb5f7c762d2a5d8901b8970da1293bf072844c3e333c0f2639b0b937a406a797e86c4e68ae1b730f0747c564d06c33ff48dc6a51d5d6c9aeaa79165efb715af3239588fe12c1fdcafcec3d0daeac70306d2a65503e950242ca5b6107fde74cdd9fd8ec946219b5a22b920b19bb5e774c33d05a8b688d33a2c41bf9b25601411e4069421929f95243d54878759ac16316fe7d4d7d732d7bb43c21ce974e0d981238c1363416525eecfe7ed1aa935ec20dafde91c186bf7c97833b3d3a2442a82dc4cac7169d5787dc2ca005c3775b38ca26fd613871dd298e01c728fe42776fb5f91559f93df03faf233d3a37ddac48d420d35ad6220430;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'heb87d4169295cfcd8d9e1af9aafd931fb3a948b883f1faf8657875e2f4ca6bad9adf1e05f2d82a941dd26ca7f4268af27e826503a5b98d1e84033fddfbe4391e6320c0819f6cae1fb01df8e6ee3608c93eee5f830ab34ed2b53c479a5f93c1a2d298ebd13e833da7fd8db185824cb6a3917c932849d8f7f4e76cefaf75440e1399e94b4e3def1a17fc7feae7484b7525474254a732611a904d3cfc90de8bbd4005404c8a7b97b8eab0a62303976e9cf5dae15a39a5827873a372066e18f5d12b3fc84104b21a97a34d9f123d7432ef0af188117c873d8d7f1e4bb09c0e74a6747994c8375fce34f6f3c7e0316efbc34962f4880b108295afff3ace21aa6bf6746239448ba5032019d740c586ae68e02b24c1966f338b3dd76994462a11a91a19bc80350cac9065f5293adf5dfd461fd37780988dc02ab3476d5f32e984fa3ca0110a1721af0e04919da2baed84884d1e1f5ea0609aa4b5b79639caf73b695b132821788b508124a3dcd21c547ae1130d26379b48d225546ec1e46a51c8555dff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h2ceaee0d3827f039e6b88b9528a3fc4a2d23b3aaaf998b7027e4db00eda3d97bf27813723f1019c33cc1acecde7848748c39c8be2453a3a9a20cca32399c1a69d48dd481d7f266ef0a83605bd581057a4bff30e60efe4fa6954e4e6f604917762b7f088beddfda0d12d9ccd5570dac5a14fa27af3dd360600b4f90a9d873041e7c0e59ae0cabba621845c4c768b7ffadb1dfe70babc8194decc078731d6bb0b5331d25d5032f0bcba2e0181fa1b6052f134b7c7fcbcbcafdd7b7043ea5d35e98458b8317420af544f59f6d73d96c3521b9a39b528dd53c471539a55983b9692fcc6f6f978d88a86f7accd21f17e249cc62dc34f04948bfb1fb24784a14508dc562d140c12ac2f0d6fd5d6f5ca1a2a8c6b5c82327cf20bba47fd78654b58a3a87102fd77d5b029908a15d0e3e5a35bbc9bed33839c25ac452453af20e745e5dee5de3d04fe1a66cfff2c43b0159ab6c2a611079cd158e9eb190b7d0217ac7d62afc4c5e8881a2b7b3e584b3f2b8a154581326aeeca7b61bbe66425147fbc74dd4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he874a13a821a8de0ba92dccc1b4e9d5b99563c06397e04ad878c89b5ae1234ad935abaf325bd39b887cb7189aafffdde001e827ac58b97d0953c30596f41ee00b60f8fd70a160276e5a1868f8f10e367f7229e153cc0384b0d2616db68f42086d6def961c82199586ea820093a91ea7667fbc2bd904349b026363bca1d2b8520d931af38d312d59bbc6f59e2d9f7e3fb4a43b122235f40e138d15e90dcf061e14b6085ce3752402266b58149da14b31ceba6a372521099086f46dcb842a8893e8a558e90bd26f8291cfe01f8cc14641001ec18a6ad89d51b335f742feb3b778bb13e0617a943c3340fd629b5bf75b7c9859b886fc311287d009a1f054c7035c98a86b21c36aa43057bf6cf9edb88e4fb49a79033dfba67c0663079778482772b44d24b7854dd59fed08cf34c70d58f568b5b7e08665dffdd69f41da7026e830cddd44684e91f5b1ede98085184cccd1a6e44f11d0c28229080733252468057ea256a91f7e7012676afb5901674205fcc16a449ba1535fa7c5ac07872a29c8fb0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h7f64d9fac72c961608f5eebd59fe2f0e71d0301feae7714476e24b62a616ea1325888968627a0dfb5f440b56a3c80f1183a202b6d99fdb4c024398c7bb5eebf2b6a7d0b25bf34ba49145b2ba3d88741893ca896c78b5a1cf508ab0b7b5bd79fbe477d9b0ce8288c6ef7dbac7e665a738ed8fda0014c469f9d41998b77d578eddd5ab914e50df30ca761cf166e890e486b5c661c44960b0ca8a76091e65d91e6e622269a771d3e5510a5e9a07464da1f65f753d25f0f3c0226324345562053a8745c4a6294824738dfbf53922b9a41e4985c0a9b89680b10909c91f3dbcaed18d958188de9e2f00ef281bbeb6d6949775753677a32863d7bf1adc694590da7642178d1baf7b704ad10aefef9b7fb01397c546f916ddadb7e6bd97d80ea1103c0fe0d0e1c6d145f5239adc31beafe7f48935087a6e108c570cd8f29dfea1248131ac2b1dedb6b3d63e10c51433d032029d331c0d8deb05ed5a6c4e653a98c04ee43399495f138f7fdf2815f9ddab91f9c2127703b548a2cb9ca7a074ac0d996201;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd66bf0147396392a2468da267e11c74ab9dca36bfd77a62270f5e5855d710ae80ba45715b5ea6ad22071cd3008a920dc243f32a98efe57c56c2fc92f61e379b77902ad3dd7c130e1128e89d4cea1e5d31199b7b7862af3dcaeb76aebe664ba981051017527d4984d3e32fa50fb1b1ab292b10c5a94b560b6be0fd24f00c1c91f7653860542fd60b3a89f4e2b7f4f3e6e914df2ef90e2b688bb4603878683cf3f600be03f4d7a28447f083417e66434019038b6355908eae511abecf6a1aba88b98c5ad44c55c146434be461153d2b073967351d136ed98bc369598d7faec8055d80c72cd2cfa801b96a18fc1538c7252412a6f57e163891edf9d98973d5a2c1c537aea6917a97e54478582a0139998531172fed7ad8eefa9a7b5cedc861eb1d478e8dc7bfa87eedd50d5b67e7a65815aa56a5a72669ad1e2b502cd355a7919ed262cb9a46511743d833c61db65854b938ee9a61ca66c0ca14d32a5ad97819333b5351a0192c8891d281ba759b47117956c979f1d60ec2bd6db68f3fb2bb47576;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h7a92040ecf5d15d5e94fc5deb99f2ef0926e60f8c0a8140ebb50125689ecd9e12a1ac108bb43feeef9cb218a7857624da46a6625e40bb5fad7c5dc68d234975aa38c7e624a69af36acb032983fe1757b247d307413bd7b18bec5b64fc864b7dd14f8afcf438e08cd85479a6a1b33fb0634260b683f352d02b4c8fcb85eb30c6660db31f3e3d48dc28e4a704a4704276f24e46d8c30a91fe797e7d183e494adf45dadd5d04c492f2675a320f44f05453fe3927c9c2da80d650ca5051dfb41fef8cc7b9ba3e425b65c9cc8a935e6915c531faeb2d87cb6abeeb81396701fb25b0d5b0be566da9574d4aaf8970c5e8baf36a6f616b818b6bf80a41a5d8941edc11257312da63b944db7aec3197278ee84200e3b6e0312ca8d28c4209d194abbe76ec5ad6edff1847430e4bd3bffbd15e449890fa07c6ecd639b06e51934029d47173757a610cf5d3868e946f0a3b41ac6462a930ecb5a4a321ccfdd3c975858f809626ae17d9291f020f852181a8bde83d2f60944f0bb71e1aa3ce138c5e7b6da27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3f0534c4a50b8fe8180a36209e669e68e9b20e674ee4fc37b6d790ae7a23fe382b62055c4eaae9dca295e5d868434746ab4aefa1fe336c8db1573b9feff54725d73f17288fa1a8cfa90c86beb3d12d037187fdf79f8cf8c68138afcc88cd94893facb644feeb92791af4262c48c1f898a0bab01456764dafeefb345b3fcb0bbe8ac8d7c4407bede279fc3515abee09d09d0b98341ea6dcd510d620b722ece6fe8f187a32c009a5a0c8c6722059b1155ceb3ae3e2e38a6d81788d6a366361f60b0fa2ea0cf745a357f8bc1044778f1b45eefe8ce94d40ce981af40ba0ceb67f6da6608bc9ea11f1153da9129dce6ac3f84396a14cee7eedc0cedf5190867508f2b55b5012ef76a788c4da132ae48d98d2a572b66190f48a8c1294f83a097876ecd2f76cf0a20e903523c9f69cea6f240705792866f32e6282806168c4443d7161566da78efc99fba9251e4a0c67c7063a4dedf0f3c451ffca974d429549e3f37b52d722079854ef6676e2bed7ccba09bb14e3c586bef66178d51547d694a9305c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h43c0a449b9f05eb0fd146c73ece2717d901ee49b12378139e723356ebf9b718648c7c376308394c4af2cfd13cc643900c675fc1d92c018374d7af1190dea9826bd140ea1f4f0278f9ce0158a97808230cdc3826ae722f22ee9186012b1c3ff2e07efd113bfccbf8e2303c14b7de288ce8efd5c969b1a5e15fe72235ba7bfb4fd5fc0b9d0d009e26d455a24b519113eec9788384cdc1cad9f8bbea3c1ab22e2aa02c4460a7ad2fe8c36f7feedbdc9a2d5e66411dd56911a8c67e4013bd94066c0de8b0a638729864dd02f32d9fdd961ffb4956518155cc211f1255fac5612a3a5fd6129ee32b3c1a526bcbdd769b74098a47eb84b57ed1000f8b1880e3212b0261f4ea639af5f94304c0724fc5154b2839d0dacb1f693d40246ef8010297a3c191cffaae1215293b81e1c33fe191bdc47418eea91f8d1f261367b21570fd3004e435ae4977b637647a4c04e697176321feb312d74983cb0a959e0cc330e96a220703715cd8afb6a7c956ecb2918ed595ace12d17f069ced2dc7e983ad7d9780fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf8ca9f45a6b5180655c5e041ae39c6ffa98637c1566adeb789cc09b8e29e73ee79bcc5ddcbfbee5b2960f8655869e53c74a4d9ac2316a68076b95b5e1b8f5e4aefa0e8ae490312e02283e3d1a9d672dc6c8e828a5b83edd69ce4a926025ff983e3285be0e3cb4dcd68f5cc70faef587897917b07c6332968aeca81c94729f80f268fc79fdf90e6aedd4bee83e1bf6b01128ef2616667cc159b35b93d2cf45aa91c4f7f784ccca3668512246019786d683a21c57b601303a783cab309e5cd7aebe5b89cc12c40443ef61bde87b08df6449ff487797e1e784528877c9fd03d38b0f48ade4fee70dfb325670ed76f1e0116abdb55bda37f8df6f30d268cc25b6ae12815b6b5e60f771bf2e0197fd633a9c369e2ff427388218323c5144e7999f87fac6889d2362c79dd2392e555068b82e3187a5a97933f46d74e03e89a7961e77de0afa53b4433bfa22edea76fa1fcc491caf0087f5d6f2b0ba2e43c22a126ccbe27981d3aaedb67eebd27fc53757e988919540cecba2ff8baf97ad963fa3efa43;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf5f6e9b6994c0a882aaea45110d6e5e7d26156b92cdb2981ae7e984dcc48a471ed6c29e3fa42bd45f011902fb6c122b2ecec1a79d65d0896fab488004028c6f1ef74df5be6dc0f0dd77b6892b84b1e055881c06c7ad057c70cb6998f8396d8d3179dbb46360f9f27b90199023b5b508905eeea9050d3b507a08c927c8cd686c75aa9990fcbe59b60dc5429404cca7943538e616b584948a6cea2af3e8ea100712e8b269a7653fa5f4cdcc79f2c426803ccc6605a8b3fcb22f71848834c66c487d9c8a93fc4c9797cd01423068dea16d1df5d4c28661b19ba2953fa8787272560b05310d24a87fdea89975d7a7bdc6068e6f4998f9df2c4e7c721506580e678bccd5d3465b5cde84d5179dc967114ad2b2f57d530e531a071d578c29d23d009b1f2b9655a102030bf563a5d21477e13b46bec97796f2d219ebeb4eaabc1d85cf72716e87f2c479783e421cafb137dab12e3e71c378acfc9ccb7cea9150b3097fd1c69258091e1e2b22ab78e1354cdfbd0df081f999569b87efbe910fc8e7d2da6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5d90fe1cd6fa280b2700f875074ecd232990e49293d8972e40ed67e1c6d597bf114052c7a4226d2783fde898f618eb2f286b4d946613ce8a524b896bb7068ed70f1467ab073c5a6ad6e904992d5bc77d257dc1fb5daabe5587c6dc082db571fd2720f8e0e1cbcd7ab32c47f140fd4d22437605e9bd149b35a7b1ecc5c04d6b599847416b5698ec355b45df227562664cb4116a0319c8389c555759cd17ff63292ac8e7bb95057ee04848dbc1c2396acb1cfaa96df7a8d40f1be4581a431408cd32f8fc97cfec8db908e26c499f5dac539542880e1b7716cae22bdb916ee4c29ecdad00798cad404e1ba76bcd8681a7302a6388098e46d9bec35f0bcadbc58472314907c81d83d13b782486bcc8963446d4894fb140feebe3b244c8a26478a1469e551dc761ba324b72f4353ee37cb68f03df64e0510181ec5396cc9b8fde0847db75d659431bd7951f2547da9bfd84f98486bedb069c765fc807a281bd1fb90704d7c9586965057cea27aaaf72cfb161467714ad7b8033afb287341e97d9e19;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha5f46e4c9f07432d1d844f5f529ac9c7c8df5e98fb76df072d65b6389ea8180616b8a077bb2d48decf822b65066c533bffb0c160d81bd0bd84b0722f114e447de44982f068218ea169022dc651687626203cd7e7b8cb09a495ad8d8492c7c6d3c09245116d1730f06053d5de4ddc32afa828e222c0c2cc73b1476fc9293a3e429f390588e63609605e8fed1ce0bc66f28ce77713fa8941c9b8a0864ed3e110a81516886997a7c7c396edfdeb76f4851fbc48bddc5b055bd0ce04b0413858736886fa48a3d988a9d15939d9dc656765f4d11bec4efb9dc34fa60561140b697dac0c01b1a5e84699f2bc041f995ec5b223863fda13990e2ca3bace68beb252236e9e0cbc0c2ad511dc6b9b315dc3c2f5a1bfe186d4e09a9a1ebb28b86a3368f35d3b4949274c6750610b64c4592d6069c060c2b385573feaae401326ba5aac31ec6ad95261bcca39a855d142e2dcea9dc5d56e29ea6b577993d97081bd40a1b549d052ddfaf8657c0c72dafefe07376922a862823e50a32fab97c3164e2282fb5c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hea73efe6e2c31b461d5210927a22fcd8e092b9cbba7fd356fd27d3bd4d1b201d1dd1b184424c83b2f6cd5896b5891cfdbad0c3f45ce2700dfdc989304e178bb8a23677ac9aff0ed69624e7f4b71f06cbe4c0709f3e85da1585e761b0231183fda0b74d61e3325b33735c5b7a1e56fbc9d54792bd7e534fe5d147c03a2e5fe24f439c9eb783e03cf370c07c2ac4f7c0ad635b7f7bd0c8800f6102283edb76b8cc287a8566fd4decdf3cd1aa7365486ff4a8c0f1bf0b528d499a44ccf68986e352fa09baab5e02347bd51c3f252ae14a05e73103a1ef5fb061e09c1fa08169548d5c22c916436a5b7531ada14befc04bca3488a2a619370214d996bf4a7a086c0f0f87c81d68a7fc504f377d12d42c1b222e85aea0370b90d778af1a2e22d262a9c94c6aa20978c2c8afd6a11070feb66879218412558a7dd9cdea5d72a994d58f176a67143fbdebfa4c56beffafef1e1a248b69f848167be0a3e350c69260ffc87eeb6d34bae59b8558c4d8163b4cc5cd7e788b62c98e120ffc1e01c3fc430e4b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h35d80c86802125f87e8695f05b8e1f84e170eba71a497882c00125c034450cf8c3ffcdb3cf51b0e9e9c517d3bba80d9abcaa35a48caf3c9542bf3d3fddbe648accf1965786fe36b518cc878d8e0ecd4b14d483f8e9c48b759dc571651f3890cde8a9ef1e465d0e070dd90cd40a2a62b1c326135dd6a65e1db0de1577519ef4d8114245a7fa7f7ee1171862f864144f05efdc6751aa686af1f05fecdec57f0e46c64e244c6c863fda0385a9c46b8d12df69d22681bc18eac6d9f86657c7e534fdb1f62bdda2e7dd6d7de012065b6c2c48f089709bf3352e97decded6784a5c006f8bbc7313244874eb350b5f9ae9269e5ec1fbfe3e5be7eb91d13fa3dc0377256cd2ac8e295eb807ba16b82a46e0200a4aeaf300411672e61d018a3b2d26c0ba04ac4b67b7349a2d3c0b522dfbdf11d2a271ebb91c1aa85ee48f499a658d414e41382f107e8600792e5e304e4b58b236e496726c4ad5e028d9e457c3320961ee437b683533b043dd9e09f30598905e3227f80192e07254f7e375feffc392ee69a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3575997f529a3018c6eb22261124182367663a1d1261862b36fe779a938caa50804a8a2b5266c81e4bcd7cda5226d30dce63738255008ddbabe9f90fcb76652af8409b8fa28c164ec5ec7c9a0b42ac629c0d00e758c69e6bcdf56e31c0cfa28eaec3c18e3a9670699aae93018ccf49cced97f2ffe4cc8df32775301dc5f550d6f916477f1e247dfab81c8e14f83957063c7714fd2ca808d4e28937bc6f2f21b889aa7a6d421f8111843ac6ac1a75b3e8a35749d93e50ca8c96679d1135456d521fb81ad560272e20b76a8644edd2158f278be835d6ae85d771c794642aa32a3a9d41aa9a603a1eeafdf28ea4f7353019477a88ca61a1913916bbff9024056f1aea89612beae178a688b52504b86974df4a4730f10de82206fff57e4ee0181461381625a2e111dde0b03504db53801e304d4a74a5826d0d4fd3d43b9f4f3bfacb4a7ba1c36c3342dbe9c75cffbfd8e078579c9129dd9394ec594fc2c6c3a987466fa98f5043d79e7da156b7322ed3e77bbe17b05aaa3984838dfa757e270abd9e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h7c8b6bec97e53838346f3844cf312b16623bdcd9c9753d17434b3c6ab6e11e6f22e116c4868d9d3ebdad8397a3b236b5cf8e6b565999a3cd33e120e5590a9236164a2394246652181884ecf3768ad24ef3030f9e0de809932eeb6b8c155e9d491077b0391107882fdb20aac75d519f1ef0942c68f03d35a2cefaf3b18bbb1b8234e8652d490c75da8c432037da2558422f3bc439b8c96e8c79c1f276550e1dd7c1cc7edb90e42268755144cb1bcb2b428babba1ad20b2bf044d0e3114477c89fd9bd32342cd0214c7aad9c1d0bb2618ce4e1e5620e080ec2a1372a807bba39c3278de41f70c26f2c8a8bb40ed5b2cf9be5b18e56215ff0f3d91e4961dcdb83c02e49b0e7ad70447a86dac4bc720b44c55c32a94bd5777a87f018f38587070556da50992e28e5ba268bd7a55f1b849794bc0e16f370228eefb38a66303fd61b339bdb1bbcd5ab63b91821b2db527b32ffddbf4c2d4a02b3875a5b01b19f1a1c8dcffc3afb2403badfb03767fb1e6c33bb236b9a61fe1564e136d27c9673972ce2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h63475d9fd5349e87610b5bee601fcc6a202e9ab0643a2b35e8a122973f7cdfe3dadf44da3b589637df505791d20e991c99e53ec16506ac8f83fa6a520f4319c813eaac333ed62b8e445e8995ec669ea391d7f3dd20cd442f013042f958be3bc32241d53d5ab81b1cb87ec32bf9aa3a90f7217865126562e5de1b2c9c7d5af599e212fa8b0e19fdf3200c7578ae6a95b2553bcdb13a5460ac4e77731e2c7f0da2c136926902be5bffd5bf5c231c0617b8f765e1ed0fa2d8c8109028ff5818465c5d64055c1eb38609dbb8a93f0d71da5d44a9adea1d0bb43de2cea618e5565e51a3e8d1893331a48656cf59bba4930a7d6b3a23cbbaf119a66e5aee1dba6e2cee353136c840079861a2e4103daef47a6f2dc80471e5c9599eab17a22896eadbbb1542051c5f4e5518a1fe6b09d2a3b4487697dad0645c4d471e81af165e05be7ebc292d0f590b162e98e551c0af0c4ce5fcbcb948df3ae74e211819aaa6ddc69560085a4e73e30ac26e7fd02a6dd55a8af28d27a33cb8a31b795d0afa224347be;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h63be2c4b6ef246fcd5bf0fb29e7d5205a6c466a182128eee5de5a3c3ba652fcae69e8f8cead425973d37e26057545e52032837f2fbf4599f971d59f949563a7ecc03a9b0aa0360334b3425c5bcd825d104e267bbbfeb6d52c29344a8e166648938ac0410e11edeb234940df46aba71dd4058a2bab4f42f666063a8bdb4c1a7a97c1e6e0d9cb36dc16a7870175239883f29777634e31cf3bd3cf0f13a3ef3d158f01c3ce0be53ad55427e305a5c1a4f42203dfeaea280bdea217258cb4ca634febbc3da8a397328065a2957e19ad1510f92da98e957431e5d2a8c2cc13213509cdf9c66c6ca5286b4e36598a1b7a5bc63b434c4a3312dacc2fda90423fe72743f6dff6ebe22f00b48756bcd7ee0a15a8648c0b08951e1a8b3e3ab8611d1269af2791bc06f64edb7df055194c355f3b17885c448698fcc58dbd804104544bca8cb4212b09ad7a39092938385fb012d9bec2a05962fd989ee4538c53175e0db330da77ff8b2a4d1c5eb8045af20554bd3d5e31581da09b08196a90e3d99d832d181;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd2d331731d45efe967ad8ad032320ee7295f304f0bace8f136880b8a4d5ce20daa1b63d03e98312ca105539785212832cec53d5bb99683185749ce9b4c91cc248bf1253615e514f69339b255e7f2468b033cc09b6caaf4a57c1809f5f7e477139f6e8d9bd72015d83bc9199292fdbc351cd67365f260b225c1d530d78a9cf9c98312f1390593da6a42ab1271b147126346aceada57eaa666d03e46d689d85573bb0cf685f71f814b26bb056c9a2a226cba5de75e54dc5d0c29dab7d54269744c61a8f314711c8e419025406b121ccdcbd1ba21c422ac92ff873f0bf0d46e3f4c719865b52aac058b2c094a86bfd6dca16cd96bf69a396415409445eb97b2c73e39de6e4c442462a3dd159c2f083e78e09aff2baa2c4b26c5f459e893fef7941b30dd5e5937ab23eee0ff32f8cdcef3ccd96aeb3fed0d1885f5ab92f7cf2740c6edf98cada9a23e77d8e0f3f5268d8e8c8e2df9aef5ccb9980ae4d0fb1e6babe588b089639fd3d0813f9d0d6add493a53d01e42057f6af2b863473a1ab5240961;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf0fe0ed0be328b1dec3600462ada5210659f21d886c6f6ba291144619b96445f7c4ffbcf0b8bc7216e1d487e972d76410972d228b5b149f8b9946832e3a6afbf2b48c3b3c1445dd61f74838c06c8b4670ca5b84c03b9035a40c20eacf07555f106e8c45cfbb0a00936aa20023c00bad73a4b36eccdb831778f2d479bb580d1fbc6ee7cd4bb065f0e525747536207014a0e7f89f7f10bdd8c0d10383deb934823c19cb2e1e95b3d0606cb76b88ec4ec07a20237259da93b6d60eec640de05a40b8d45b426814c6272069f7da7b656fe5d06ae2fca8437e000b0f36829aca308ac62847b385f865762e82357e32360a363d4c3e379a24ff7c98b408061bf6e50a1fcd196cf7e12cd16579bd44446dff44e73513ddc69698012ace56999242ac33b4d5cb74c869bc878325c7d1da92d85fa8cbd6b04e29bbf5e0a2983068db63782b4103b3f848315f2aa6d3ec97e395640aa04fa9b7e29490bcb464f6a86d1cedb7f8c8bc39c61056187d43ecbeba1171a530120eed3573a61cd2dab6c64be8e89;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h72ec14a13a23ddafa261b300d68f40bb3e499a703b538401a4d4a193774cbefa1e6f6da035923c439ada07fc42bc0de4d102460e6247ab515f39801e61cd9eba1678f0b8384e22de3a7b3f81052c1e893c3ea595606202a6ab56e6728df61f117eaa401759565e0653065b69ed8229f6f4a2930b5a3542ee39ebe3807efc0a247154659e17f6a7a7f74924731e176061d8caa7d40f391e895bdd075c4e9b1d1a59a1ad9558190725d37a21f1d0edc5606409897db0f4468f2b5417eba9771183d77623c779edc68b6e090f5417abad13ad51ea0e616f0890996b6fb428e093faae9ecb0ab3b2c4f75d89f6adaf519e2aed60b6d814ac3f309e47c2a2c18c4ebe07ba995f111a368503c470312878a80f7cb621f90643323e8a93f7ed5ab4b48c4b6c66b69626e9d4e7fbaa6325b4ec7ac2883821487925d19efca42793231db4579d77c8b0eb68ef4224c09de948980a95e7c3b7089d2aef898c6fc603737150056eae343842e91cdb79978f96236f36484e8006e34293bd4ff7b41ec7881a82;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h96a02b13109a2d6882b8435661476aadc7c5dc6f3f6cc9943dcb3d63a402babfe1c1a0c13f3fd4010fe8ab28d7474bce651b02c2ddf16dd7c8daae239d7be4745e88debe86fc936d5ce18f647157a0cdbbcc347ced019de2aa428f284f3d0fa0a384c983fc5f36d30547e8c6b6411218b7699eb7ead8d7fafdc4cba5aa0d765d9adaf0998279f92ca526a661c4cf445441eec8b4d88c1ab1fe6ec1cc69fe1b19b32a79a1e72a98a2cb63addc4f30b4f59dfb8db88bde05d0e83fbc62fc886d2ba0493e13c784496f9d40ad7ef234c28a59fe45ed099c199d748182bb796dc8d37979a7fcfaa9415b3ec9aa63f7a017107025b5c6d6074547d20c70f6ec825e8b7f89bf339ce48defa5fff94ab3954f2f3878c2f2114a414c54693d3879b623ed973c06d901a55d2320111a1484e36c44d13e2814fb6f477bdeab192fbaeef0620445ce2bbcbb4857b49fc6b170027d70046156527013076fa45e764cadb4527e6f4c1ab73302e5a9065ac46deefffc84fc96682946b99e68bab6bd7ecfb0ee3d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h199668fbc6bee08e54e9bca1d2bf0d4482ee69d78ae32ba865c535648230450f5beafb3d7a4b176f64a44b3e34f1d068dad791ecf2ef4e8092ed0847c51e1c23d9877d11cb99a50413ffb93d32fe669244f619da90924a25ab747abf18e4c1818ad0cf42f8ac466ae84185e0da6b2d3d71073cea4aa31352461ea79250d43383a4ce62467225244162dc09b88e85c71d4a435b0f5f22c3efe883c6dc92a9ecf726011f5db9ab0f74ca7c1410952d94270bfc889c3ebfd99d81aaaacd2719ec86a61397896ce0234b4697bc62ad3104198e35ced7636756ba352cd2a255fc093658c85ecdb7174ce1f41973a727913b2bdba489347576540f364dae3b8c713aead90abe2ee88dbd34cdc0a98a78d0ad6acb1ad231059e759ccb15637c206b223f51183a59f6253273c2b8a86c1c5b2400a961dbc2773e0d01df9c8c2df829d735f34b6e62666c5f0fc8fb38bbdc92c352a497682957d2743d180ad6e1a18070ab64ddd3048f7da9f6b246214460155d87287780c8b08eb655b9bfa65d14f94bf2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he4651fed298133a92fb49030a7d2459f0b33f3cac549d914dcafb1a68b168ad85acdff58502121bdc39a7730784903c86e38b1ca247f37ad74f7aa96056caa3a0c4fe144d3faaa5bf2f53b597fbac41c85f49f0a843530b88eef6593af528eab0e4cf87ecdb6cec00edbd8b0b752b29861cdab9e26a6331783b52c5c1721c0e7722df516db6b724c7d30c45001f10e2b2e2a7bbe68a475cc5a7b2610bd1b56306a36bd418fefd704894b1030800bf80bf756cb89ee3eb9e25db3f703a46ec246d5ffd4fcbd7844ce1323563131be60a4ea5c0fcd2b8201577d267c4eba3f2be4a3f3278e9eb99cf56918801a89c4ab3033c5e0bfc7ca38dd2f1e20cb2bdb69ed2b40eaebd9a0cbb0dffb9e7249ed0c68a3cf98d1436cc588a9b36775de673f275aaaf99e7c3f2d47f217c107cf03ca7bef2e42ed6689deab4a069592af0ef86b7527df7259c6335460a16a3ad989c667dfb986ae9c1ef5a5c034f029e266efbfa0b26eb90454e2cd6ca01874fbac9110e62bb3c9dee68b34f60babf0bf5d6b03;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h6ba86b64635ca09c4beb90c02fcc5b71922787fcf8964db436c849e22fde76ff1188f5acdea56f6963c7dd8d341d9a3fa8fee5bed77add8f21d30a010e299b1ffe4f04cedab6c573c14bfbe6c761f70b6a8a28d89be1dba66751e3d80f3799ee46dca34dbbd2bcc8c5c4cd789929e06e6d1ae23e6f607f797326d3cbccf7d070cd1c9df1f114cc0edac5eaa0af7e4a35fca6f51442d17861cbe62eb0d3ba9644066051b38230b00410146ddb711ca78671fd7f12906c19d3551e1f2978f4273852c9d658fd21e9b2567f6d45a82bf700e19b137bba98b0fada3f7950ce978e5dc4550733ad3d7e1b6a65d8079a327c550b59fa8d538089d7fcd6f5b3e8c2c44ab73c843f2da368688fd37fd383d60512727df58024814233d8d5d982da064d295dfb33002292765a302a28752b0f0d743cb60c863f99444e8cacf0d0b49818fd62ba48add1dd20eef410fe125cb3722acd1cba1f09cd9c77f9f6c83730e564457efb787647d600933a8b69312a15184e6b9ae779eb706f086688ce4ba7e4a6ec;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h73491ada0e8c82deeb6fd47c9ed9a6d9349f7d452f6110fe4467eee9ff8fd38735f2e66355543e92c74bb3191e2517e42e3aa0d6b0ec3f61d525b2a15c47d7a1abda810c6a9a85dca16067e9b5d423b7a65606a251fa6acf5c81255aecc3098139f28a018ae4abf2365e54b30e815e2395f281a700f31712d2a925e4715eb862198674c4b098889a78f4c9a685a670099eebf40c9847f094c3568483ea1621db2a67585d9e49a89bb7ff47016ffb04c644a18cbf990fb1571f8db249cfa7aaa27624d639a8126226d8c4a827ce067d07453d16bfe218c855d9bce4e4a728228cc63058dad2170bbc88c5ea817b8241832030e76751b6a16e83808dd11fe25f3c3f155b0f9ee2a2b1ecf2336127d2dd47b44faefe29815f86ea4d02684e4f1041ad5362f0e6a95af1002e1ffbfcfd006207cefaf4d4b0a49cad3aa75299e4aaf42be1ce45e257f171a15b7023f3575900c095a72c5e07a2b23c4597ad69fbb66e7511997504678116ad3f987d10c911f4cfef29902756e4394a672be4402ad983;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h6fced19258e1dac30caa360aa87b090ac0f023c33aee683325c31d5226d67352576d68ba33b02ca76a2d4ed1d1b68af8cdc61f79110f1c6b8179d25bcdf9fe29614e8a333c46d7411d4f8fef85ce80559ac61056fab382b9b68b77a24a93c6d8eb4385d66dc83f0db74e1a57a1da62da98f4ae72d369aefc97c1c7ef4b7d9ae47c972bcb999d34d9196b20dc54e3ef91418d78f4f25e9bc3599877d4fafbd2b159e24ab6ea68a94903f2661300086532360fab3bbc4d86de1ce3025ac5dcedbd8283c17174d37be947eab2a6b7374de079640d51cfe8c29d0396cd8ffa71f8f74414ac66cda45ccd0f18edadd65b3a8814810d9b573a5b6776f3e74333bf89e9614f92acdb14b74a7a759e9926e0312014fb2904216170db89780c546f51c1c3f35c50799741354cfe567778ea6d6cfb42cdec2adc66c390618793d962f7b17881d595b9692444879c5255717a89cc981af8dc6f1f04990e17f46854688195480e3ec6915f220f770dec290314dae0a6c7d1003c23f68dfc1fde04fd91679273;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h926abb0f97f08e527be38c5665f09a658e807a0adb56b8f13aaaed469e37fd9827138228619839f6fae8a528a2e8d23ae5dfcf83cbc1f62a6d62ce57db80256e0632884ebdaf8ba4b97be6e87bc7894195ccd835bbed0c4f55a2b696e3b709a792fd35376d5c6908e8ea335b84078a0c2ba3241f2261eb997bd38a19eb5267e79dfe16237f4fa57236cc8a9cb33b7fc7e74e43ec18c5f69b35dc5f06876c2936a95a6cf0aeb9cdc0d0cd50c50ee3fb87639f0a2c03f70c0c55b6420e576fa07f11e95887d55a9a460ef3044c5ebee688cd173c33f48a6a86ece586ac37d723305ef39646d2e93c258b93c9f41314e04588f7a22ae36af8fd3e358b0714d035bfd0f5493b081e2c1890737674c58f0c65802d18ee3cfdcb22ed4e661131c58ea690eb099ed42e6c1d102162a0e64d933606f1f14fdf5441428277e82ee4420cc015d78fa723f3f70745e0f6b7e5b8ed3336f405ebd7b952792e91683071b26a2dde9d60dea0ce8d1b39f462951c9f8dbb3697002f0d28f212fc0f7c5ebad819fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4de658b06b94d1f12f8c9ec01dd511ba51ac1f21c09890553ef1a5decf708dffc091fb1ef6464c82d5b5be0def4da159d3f4cd90ae5211646d0d777d34df4b5e40e9999a40ba7e1b01648f36e98e22be1807abeccd74aff43086d07f237abe79c6e61a9e1d50ee856f3b4a1a6a843556ba8ab206bb545f6d60a9d4dda18224502391368542bb5ed4b394f98c4926f57be79b2c292559785af2987765df476a1ebb701b2b39ab3bb998aa708e9a8444f390e9bbb3124136394b0a599f4a2b33690432040db73ca71de4f0c27c415c2e2737d19c881580de6c771c4b08071496661b9651a023f343bff59418f4dced6bbca8328aae1b33afef800f282f1c3fce406ddbfc5b96a74387c3367d11419cf42ab3852671434648b97a9f4c661316525761868f21e129dbd822770f7f4e5fb833df31308cf281a0e064944bbe550b270d669c2884915a9053b0a382d468eb67d79ca849e74a75421162f6c3b64b272671089de8a928e331f15ce24d339562601cf99e81fa0ad1c0771abf324de2b5facb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf8c6f61d044bdb8b70408c854ace36cef7e743d9bad51bd88f459759324643ef97fd3a49e8c0144d6d0be5be00a23852f0a75c717d3021aa912f1085ff39d75113cf583fe40823e39ebd81f96f6d1bd8093ebae38413a649591af0a8f58ef335282020535de2184f2cb65c7d40c6ddd96154de488a7526aa1a03c3620f6866473099321dacd20aa476791f3f91bed580da2e0307c1ebfb7f7c34dadcaa913d57a11939ebf39c1e7c12cc9cf53e1481fbe13c2dc8e1ddc4d38d19c49e51f4a5be31311270ba9b5c70c1a51f57f04654fb4d0eae6b42aa478909aa85e65a901bb530fc59f2989f07dfcba55a2e1f4b2beedf8a169b83e56139ca2b19a23a5358de6013c8ba905c950fdd20185ec150cc710af7ea89098d349d6750af45ba5bf3849e4a99b74f9b4a7a852829a73216102efe659a92c063a45d5e7e85fa95d6ff8ae594b6879dfce0edb982d10d0287b00ca880397aae303680b724a520a67c37d5cadb05c9c751f596d3358930c017295aa56518bffe6c692dd562df5032937a58;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h235c8ecd5b033c57b336b5679c9718ffdc7cc3b57cbe5b94de74e1fedca5a6762ee84d0eb06dab58a509070f24c40a7517d4362f4facb3ca3c7bf508824203e0bfc5fbf1b31e98725ab6ead2d760f9704030315d9aba90de39221ae824f686c73a3044c86718281cb9349fcffc81051f14f1109e1af11915d06fe0d633812153983aed6e23ae7801852da37fcdf5c3e1897ad57bfbc2c5edc6eee28b477d2d79dad0cbc128d70da5e26776a0095b7c3ed8d7219b545c391871fe64cd157e1373d2b3547fe5539e941a0a6da758709035ae3659c1e14e7714a1eb1a1e16a52be6fcd052b08f0e917fb80695d68f8b2508c74653a33c44ffe0089f96f0f7cc112418e35cab5d31f8c1e919ac04d864d13f47a49ca607f307bc10bf897e65900f29eab74d7542acf74f1f6ef7d1caef2a9370b445cbfa8ac960046e51a999d275abc77ec763fb307b2f40cfbd17a16284a06666773bf4ca08d855b76fb440ad5e3b9387057bd092ec6cda53c5b17b44c56c90138ea8074cdd99b502234f8909f217;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9e43ebb8818235b79786083fdad3c37485d459f11b5673778e212653355f813e51ecac9a95e2e32fff17cc41e479a07dbf85de1936cd2d73efd9750a688b87159f69bc407ad93b70269d718782f4b7258c4ae277dbf135fe350a1fdc375a7cef68fd5a780576b525f8864e44795a69283aed26a7588fabd3fe6141d451413882f0980cdae74807ccc354d792c047af04b5636d4034dfb6af94a6f95971680886e0c8f296655e763360b8a829f0d57689e5892681cc3d828a8075a1cd1f5600c0816edeb78f293a7d5ee4d0d9cabb66692b2e5ff9de473af4e2e28c0e40d0790cc4ecb2e22f128c494fc0c4e7b262b776e188e6c610964b34770280638c787ba032a435198f8d48e79a96a8dff779de62e0f44c3840f421f5f496a9768973ed9296f3137edf22aab6dfbec5121a240133c9ce315b90ca135d9b6dda7ff6e3613900879081b73fa41e1f2f698bcfcf1f848748261f18bb0e1d43f442edbb97617e13a7d7bb2a8cd97ce09d1260ab86487da23c95cc83d7cb956d891795aebb8c65;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd8c3462e3d3e1772298ca92bb8b57fc233fb945c75f6d9311e86b12a23f4f5acae1b323d0eb8d00f358aebe2aeafdfc737b58e01973ebd3eed204c962d832b98025917b3d3b965888c02531830c5c11234c4d4e70e961e272c7a56e7af3068cf77734b67ba430d74e84ddd7266dec542d53593687656fa93ac9e6290ce6854e37aa9aef2c75df024ac753dd319af653ee3c42a9720da143a8fc20b5e62e761493db14daa06d1788390afd6dbd4efaf62448d05341526bd6c25a48d98a84249a5bcecddb1fa2a2390e82ac35d702647a0799e954ad2435309d7719b81f4010764d3565777fd6c05cbfadfcd4d45701be5c4bf9d994ac69de625e0e69ca8b54d6330e2bc44936d6d452de96e5d96b8e8e23792a5dfb556acc6596f7d5623b01ff1aa1debff6a30c6813a49162871864965be9284a39575438990fac424896838b7b85e1c97436715b7053271cfb94626bb82948692787749c3f09600499c8a894a7c2ff83c0062da9467f3ae242035406a30c1ff0b59a58756d6c0eb944511c2b1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h13829623c878e62ca15328c50093d8d24d4248004236677dd2d37031209b4ab34141ab336864a6c7803ebb1c265b9f995390b3664fb879014183f2e0f830f8f22c8e1cf8412347b6da3d9039e3fcecd4d465a1c04a367a0e731fbb21d9b146b0c7b5917bef4a62381e2c705eea54a2c7336f08578c11eb989745ba4a8239c4b92d5997bf3dde837e90987885e007f30d0ad44ba49c53fb380d79011b32ff57290aa87c29ca6e778678bf58e68583849e9808cee5e31e8c15d352e7851827489967cf51460572f1088849f48d4968d9e7172d151ff5be01a52fe9833f6256a3b556f58f9c9d281a1c855ea701deef6997aecf398143b4ee894a2db207f0b94e595d24c826f449c617412ec54636ebce470707ab6c28cd65e8d16a09fac8033f91c97d7b2827614c9b9451f1ea62ac3718fc5e8c0ca0e81663202309d2c18a77e9fe6aed7abdce5bd7af72a10f8b52658d993b3cd03d69b40b67c851e200bc11903ed9c9e46b2941b0025266a2cd4295dce3d7a8786d9915e8607a16488ab0877e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h38aca6f9679d82c8c86f8ba91aa8d4cc72b0088245ae45fb616ba9403df5b3f8173930713e17570e1fe7b819429b59e62802d864cb9fb35c43c9af35416b782d3333e27682b4adddd3165e3ec5e9a1b710bd1b5999625197412873a00022d392c11bb98a6fd44901fb6019a7289e79b66dbaa52e6d5910ebc132de0be1205f55ed494fd8848ab7379cfef51b280130b0c6d769324c90cfd25acf798c19ac04022dc2d25182fadedb05e1c41dcc086e6404e51239c3c285ab1a88b5164581c96c983d8bcb5a64f25149a3ef33ba2638446dafa958572452967c381bb9cbf8be6ebb3766852f0af9d808746e2f0b7c1a89a9d3e99eea63ca21234388d4c962f8f04820ec65147186214ec60f6b0ce9494de1deaadf59d537f275573933f7ecd82744d330f075f8d7c33ac904c9fcf6fb3472c2e55bba7bd2d1df2ac4d78889bd51b711d530e165109569e30c34af6763ac522c47ee74a336557b1dccf78199363935a0d88be85c6b52bfa9ee319083868292bb4d596824f30d02d4725a3a954e2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hefe2d943d222c4a1f3ddaaec7ded5412474c547d6657af384ac92fee670bf47e020251cf826288a8e82f2456384b80ec08319c65e8f69eb714513318932aac9a6772eb0e0bc4da25021d2a0420ea5ebccf734cde5f3d4c520e9a6c10b591c79d5e620b05bb64267b9e56e56795bc2c1f41f686fd87052aedf2540dcc94a551a74fa02e9baa6c9ba8f51244ad69f72c0d97712870b84811a924c8aaa3e23944e0baef2e19f3c39a67e90b6b43aa4c1e676b638c583a52f70fc52840858e4d4c5a82dd683c196f286baaabacf4e85f0ee81a38106ff4f43bdfa021ba92cad11519d90e00427fe6c92fea1bf6e1f56f7d40daa7e02cd7626e641398a46d8b0643fb6471e8dfb2383279588a7324b99e599aa5d2a0b49aedc993c0028b421c38a185f0c4676b76e8000998a8c9f5fdeb2efc7709db2b7e5834ff08f03212dd763497d04bdf12cb7b8e22646b3744bccec75ca2ac9a1f4b2168716b92fbe8f8c3f6052613dab25d2750018285072dffe533bedd536aeef0181d1cf0e2834e4b2c6d95;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h40b6ad9f4c49ceb41d1ead9d423c3f3e684d9ffca84da60105aeb3bfd3142b1dfe40a6287a3bfa8878621b20db1077a067889aad01de622cf020e5eefc6d6e7a630c7656351b2fb49be05f80e8ea4348f18582b17346ae7154e27286ac73139dee7a186199b5aba8f00e9d830d4fa729f33940ae83d0240c4d1a9a64333edea15ae826940b97de2d5716e3c66aef7d48ca713c7da92bf893ddde077456a49c399e266b9f8630df9091b56eab418b40f7293d7f17d48efc021748ffeb6b60d84e181bf9e83d5adfa5b5b43a01c1766ec02c126bac4498cf2a90aa717b7f3758df099d0c51b39185f157b4bb9a49b2e49261d63e6f1a7000378130bf15d1b6c56363ffe581560655fa3dcb8aaac66ff8c42abc4ce79f39776ca7b4cec5f9dc9fcf2791f1d49e702205714ef087cd92055651f6dc7115777b6ada06c2d2c6965c6ec530f1b87dab3c0a3e3e14ca0a94483c480c12f42edae7f2627e8fc37690ef8b5ca9e31b33877d55b20b19fb19499b5585377e32560c0a6ba0d9c00c49904d01;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf4061f20fe6a8daf8e57f6ebdbc79e98a1ebb5e274f5be73e37982ac5be337b1a03514cd81e4344e0fcf76619a259822f2be3430fa7d65b78c83c8d676e4e6a7fb19d7e2b14fdbaaa24125826587eb2aaddc499f1a9def293d962fcad48c1a05c5c3bb8692023e1e42a2115059454f83b56fdca5fb42a9f8eeca56bfd24c5edcab5fe748ec03038e7818cc4af8a1008e87f77007fa9994d03bbefb17c3abcecd529c45647b9cdc2c6efb4bc10bb4170fec419bd8b533e4353e6107c7a8d4e71f07865c65db0deba24a42e83ea318b84c66dfa3da246f66c9446da2dda16f083dc878a4a041f1e8e479f7dcbb1d5cf0503344866a6ab24189767ae4b81fd68098759124904914e57fbb5fa847079ba005a832db07da69a04c5d06291f8b84d37749305f454ae85f377850f9a253261babb90aa5b13210463a3da872899cadc23ccaeb4f2c19a955cb7e29b6e07c68da238daf88bb8f343f9812b72784846d8ba317044dde650ecba4d41f4e6f919ce2cce047eec8f2061ec2ba245ee003404933;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha51d78a24d5249d23a7c52e050ed51fcd731cbcd7d0cb4d97238526acd2281067b0038a53b07b9b001c93247d15e25f1d9f6d9d7cd7e230f1c61ead3d176dd40ab6b84a68d42c47cff82a79520afa8aaa8053a612d875aeb3444a8c21253608ed3efe72eb93bc1eecd6efbadb358e30fc840c3d1a56ff5d3c8c79e1c01c72b184835055219221f090a9b87cc0f216b064ac1aa7c0b89c53160aefed8e97420226fb43d03fa133c0b121e9ea395fb6146d2812726d2f2060939341251cf5213ec86f7e92accabb2ec3d09e7d63118dd1fa6578c4fdf22996eb78ebac92fe74712c80b67269c7f87f028b9c4b6ebe74a8b36c9aa98f46d192dbebcfb7e6a5ae00406fff4815c04dcf89ba9812d3b878761ad53c6fe27fe26ac23d63ca4c20e4d78316aeb475607ce47dd2dbe2dcb4f8017283005e1bfaacbac77e86a306dae3871e10764839d88c4e12aac69c69e7ca85c6034e08c8e1e029788ec4477658eb5c22e071bb2ec659a84b5fb99dd127bec1400ff5c42d645f14252f576a62c1d8d75;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9db1b5763c27813664a1b125bad562bffdb0ce70934d4b2e6e868085063780384dcdce35a882b0478d0646027e38396b7e6abc8cd5dfa7fde3a6fa5d77fa7b9e066127da00bee63ebe5397073be9866ffef7b3069463b0729c3490ae03412baee869fa71b2aaa764b56a98750490bee8f715b46f4f4f91b20f6e9b4e540bae1738fc0691433fc65c235079228db81cad59ae8560cfb8b491ea05d3edbd62a39da44ebbf89a1310b88dce037fdcb70e3f5add671f6dcb7eb9f72f5bdc0c7bcce4310224cff50b70d095e313384b9c97548d46c2dfdf425e643add4dae709cd77d22e92351e242a67d66941851f40a7fac30cfc5c6105ca788d715b8b3f0c40bfea877de9bf8fc74a4049f99378b7e58051301f33b77fcf80ad3a239aff9c20e73d21e4a1e457e38b91dd59dfaac537530bb6b0d30f54f92ffae1469b8e4dec68f46d8d23bd752451c11a82e36a93daab6a8601126e8e4040aa22f9ac53f09f7da7c19f4d437c945d22d198c6c3e2babc9e4230065f082f72366f07940f921ea2b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he54395c5d2c727c5bcc1bf20864be20a9a46558a93be18d13219e7015f583e84fe31a1504a24377d270746f4c20242f947574ebe92e5c9b426837edfc71b6d09b78a25783e3f3faf439e22ede51985138a9b1df227afd4c1b30029eb927a016a83d8ad98c75c7d4edf418c6a43d58c2c30a22b59f7ba9c184fd8d42f23c39fc39ff56429ecf7c342869f504a5676176e043faa714502acb9ffc75d257ee3dc55cf515c727b32b32cd0ce01817598f2ef958c841482bb3ceab9e833e75681ddc66d1ac4ac3acdce639dc16ed61ee7481030376b8c1972633ee68546f30cb1159dcc945bab932fa9e654d1bf3fe9697e2f5d8c2b7217775f04ceb9896324ff0e6da295d515e60805c2b887f720e7999dfb16a79901d5b6a4c6a51f08b9d5c3afd2add77e4b69a8393f007fc7e55b2ccc6c81b137a48c36d99f3b6ebff315567b396686292b7699cefca8d812545ac34205ca1c51bed24eb635c15b271dc0f26f810da3f2f7e4c594df410966517ca082ad3aaf29867013440ecc5acc0f69351bcb;
        #1
        $finish();
    end
endmodule
