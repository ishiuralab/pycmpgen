module testbench();
    reg [8:0] src0;
    reg [8:0] src1;
    reg [8:0] src2;
    reg [8:0] src3;
    reg [8:0] src4;
    reg [8:0] src5;
    reg [8:0] src6;
    reg [8:0] src7;
    reg [8:0] src8;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [12:0] srcsum;
    wire [12:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128696760387cc0ae02f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4203661d1e4ecae2874c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bfbc834a3cf17582c21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde4dde0b17f7d8e1298a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ed0d9e8a273af6334a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e848dc20e9150a83c327;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68da1fdd300f9be24e5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h734dd23ad1bfbdfbe653;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41f01662bbe13eadb338;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f34452483b6198c0f12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19cf0ffee2b8280f4ed25;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f1e0ab095097fef1e72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a9247966736bdb8bb28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10224bcb0b9961ab7c7c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de9936297fd33746c272;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfe4d68a4ab53447c519;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b70c9d300261987758f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac03572236567299c393;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179bfd21db1f0c4983fd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18330bd97e06b92fbbd85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd512dbefa1857dc0c713;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9f810fcb4240c6dc514;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc623a63bbebeb31ecf5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44b60c3cb94106d79299;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h29752919e0ca253a56ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52d36ef8ab35f3d062fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d61447a135435f896c7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d2f1d35d304f62655fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90fe20ffe1c60bc0ec39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70c86f719b8692eace9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d17c01c55da0d2b3a42e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c48ae7ca92d9b56b6d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84e7e19e869fef088c42;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12be15d93067ba0e54028;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11943df995e5bdad16936;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ef00b49dfbedd6d12d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d3c016edad47d3ee7de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1caac54d0847294b96327;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a10fcbf443b05a6839d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158c1ad35c39074cfbb4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18db83e90a71035c0ca87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10cf9de75e4067345f747;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h934d60222cce57d87956;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bac4c3ce6698d3b43c36;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc68b1cd2a24d5c9ac26b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e529f4c74ef1b1a5451;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5102df1dcd276d43811;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3443f072252937cac9e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb8675a1467b58a23585;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d69259e6f3ad674a8c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb13f8a3686ec96f428;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h644a58e4f210070e80b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b22e812ddaa023ccc5f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19def7f607b536505ce88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123bac6ed42770a77e122;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6dcdc8ce1a42d97b366c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4dd32f0e734218591bea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h184d6ab750097e7d7689a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h77e6ab9525d24bbdb46e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26453493b44db15c2a6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1624b9c9b6b4be9f6d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2120fe05d21cf72d1208;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68ed49a28b1d2b261837;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e54e209a7cc4fb6bb890;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbae7017e9d4064b7fbbc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h173ab392c137ac2423ffc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd5846187bb972b3e8a6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h574900643d9d1812a883;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3db2899226e6f5967ec6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h659ca7104cf262edf567;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h359b55d2d2583784544;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc6cce4a046e081af5deb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0aab72ee3303304446f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb9cf49d45657d74865;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h194f17d9115d8028d9cb7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habc652d6adc9b53cc6e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185037e956299392d2c3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0808158d02e86daa499;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14dd2ca87dd4d72c48b8f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aac4331d57541c209953;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7db962e69043d004b29;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42c6afc8e4d50789b3db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164d8541786b18ca3e080;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7765b1914b5e84eef6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16cc7dafd15fea9cd341;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0ca04e994a678b8d99e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a7996c2625bd160b748;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he85a6c5b5a036f7cd5ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42ef5549967153369804;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f402a8aa3d13819e2116;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13183151e98c9ef57eb10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8930e67888a6904ac8ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb692713d0b28a1989b0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58f35b7bae6c843104d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4eb0f46f9cf2486bd855;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc86f95b243a34a0dc73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d465a7b55a2b88cda90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h307cc4cb69fb70ce80ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf038bf0bfcbec448622;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f23c8ef6d1b46f0708cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d72dd052364ea302181;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1823af7e6912f6d587e49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ea17856184dff48e049;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5029a492c25ddbb473d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10bd0ad07128d65c90190;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ccb9834f4a8d4dc4deb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1d3f52fb15873e174d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda0064160ea61e3174e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb36a48861e94a923c906;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd347314a6799b3ef0f62;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168c23c7f2cde5b1e9c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1525e0c73793c9addd4f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0518b8285ecda87d12f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h130a727f32694e8596ba7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee8d832714e4252616af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e8492686d6ef534995;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd2440be98a80aa51e982;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h867a4de19a8cafb39499;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39560e6e5e653fd6e28b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a2ca3b6995d44d6b2ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h910f97f6feefdd4fa051;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3b7bde3a47b8f7612a71;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed0fbcfb2f60489d05d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8710d28e72a9f8de289;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7eb71fc4d0621c2a199;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a224b89519bac9792e1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132e6c44bfed150bf3f08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d144eead099c6d308c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h129f70d3e46bafea0545c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c33c31d7951e8d27a5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd452f4563572681f55aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf833b4fa880fdf0a8dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h363eee18d03426c3d019;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc99c4c8943702a2edf45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81a38d4b5047edffeb92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0ce40484397e3c0340c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9367369d8684a78686;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d165ed79806466d854b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1630dd662a30aa642ff0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h206310ed7c4eb5f6aa83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b42b9e9c8eb6efd3baa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14538213bd82641e77f9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5697af68bfdf1c1ad3c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddb6a1f61107d957fda2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1835f2062a6e841b49543;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c83dac24ab63e3a342d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15293fa2a99e81fe4a134;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19abef0e44588cc70213a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1130a446a5e5569a9b457;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2ed5cdc57878eb53791;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6d4131a9b600bf70699;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4aae38e678cca9b3f842;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b8aa4b59a2ae4479d7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f5f07c3173b3fac4fd2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb8e0ff12ffb31205f187;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb794e874383072fc79b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4f0e3ef47d726d8c304;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he66eb9447eaa357e2fff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a3c6395c7dd10576743;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h66aadddba03177be1a1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175f46f1bf61e770cd40c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb45ac361208e04f25bc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49c78b98972f2af6d36;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38844cc3eacfdef1f762;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d01b577197906e152cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ce78f4a0d8e51f65a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ee5fd3a2a6ee20cbe0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h544635eae07f9a1419af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3558e45c467dfa3bd93;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfdadb9475dcf4488aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb26443e590dcd690eaca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9fcd2e226b9688e21e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h65fe218d82934e60d827;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec8f2b6c6019c9189832;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bd0c89e09148d3fa5e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd70e4d787eaa876ae49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he264c10f55da2f4849ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bf87989892d29b50b43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c2c2133246309607e7b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21041b48f99c53165a0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41f49b41bef15bf1e043;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0361ab82a469e773579;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14dc068554e91f0ddf94b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7cc6ccb4de09618b089b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c064ec9addbe4993c1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aba9e688413da0769d23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fdd16711fc5af33edb25;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148ed5e1440ea992103fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9e9ab3e990330d469f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h63488d5cc485e21b7e64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef84f28a230ba1062ff0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bafbf04d1d118b8e8da6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1ede7e2dbd056dafb7a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha639137480ec2be30b6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1283563bb2be9ac4498c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h180b7952cea849d4a444e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a36ac2620248bb277327;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1071cbb008ad9be4dd67f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac936813b1236303030a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d71112aaffe7b74c6eb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c6e90cd13f73fefcc18;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h170a77b4d7634951e4ab4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c51a234af35cbd1b0e5b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc1876648f91d39846c8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b4664c46f3f23b42131;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h379a50a90209d1992b75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb0673e1a1a33cbd2dd21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd8b6b911f328e19b9d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a38f5f8795050ec9b713;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11a3f73ea481c2b67315a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e94d68e671667966c9d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb600f5d4ec6af114e47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc94282070e82b191e679;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd7ec7478c518a5ffda3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127092193279c7e1030cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce27b8e6b51d62556dfd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1497cc575f8afa832e252;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b9ba5c3e56a2fec55b47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h78ff08544faa088d561b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d94a6487242c2d738de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bdb529b684519df01958;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104dabeb425f883c51cd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13226ae2b0f563c7ced37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2fd4822f301e0367eaa3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c671052280cc38144973;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f8e28d7b0ac33dc7fca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf05a95578f9f53da728d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d5a3c8a019998ba46d51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11b07d6bc7ac6c092a251;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ca77bd6cd48f7c6225b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1782eeb2458cb8aaada6f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7598f72bc15ed34482b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h912f14794d9eeaa6a632;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f7bc95ee8264299064a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe72807aa77135e5836;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc102995acd24be2574d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144caeb14865b80095395;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h299da486b39516bc2244;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd590fb6fe1a02dfb21e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1680d6de329fbc529b481;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7018874977128e31788;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108d57b117aaf11634f76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d0d8f619117b93bdcaf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff47ad7d341600ff4da9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c993f4222691d4e50790;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4fbfcae5c98a17decef4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14621271d68d959bd31b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21cac19596bbb8d762ca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb60860fbd111b5e5525d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117ce1e3cc8aafcae6f70;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8eb2cfc3899241fdbb0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51fea750dca0161661c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddae06ca3b9bcd67a1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106ca3c8109dc3416f8f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h174a4cb980018c9704d0b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ed88ff8a52eb01d804c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha63f499b81285bd5f5c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70e068eeabcfffa259bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60e6066335970cae43b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha78a8bcc59ea2749425b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7914debb21655d20340a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d15c63a2e7a9d7daabd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1acb3778f4b548514ca33;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e77d71d6af2018ff6a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ec683ca6bd16182e58a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he68ea0a7bd8a04592ec0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1328f1ca9abc9f6b7ce9c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d5ebd66fbc693228559;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12866a251d7cc678dd424;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ebbd7cd2478d1a98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18939c67f440a635ea94b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h82cc199b3653e39612b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15948fce0794c9a8e9637;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haaca4f67c02742775960;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183bf6db29b6be3cfdc2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5da39825016670c1367;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf91180cc95b4ae319d7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b26fdb2b41e641505db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119d75256bc30c8d4a4c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152ef5767fcbd0e3c4d79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf1deb2d1ea468aeda366;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda00c69c215c1873fda0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce90fb0c26351a6ffe92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h27f4f31fed2cc4672dc0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha1a82c6601cf91fd0cab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habb10cdff89b21a8859f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3cfd04fa5c8ddb294ff4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a990672d68a51a340f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b11ce8b6d44e5b80925;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee202770f7600f79ce14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dc60c28522a5b5c200bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae2fca1a23920ccc1fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e4cea59023aaf5c0c54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1037c498e717cabef98bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d930e76ff189d7ac242;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef0d3e70a11cd4eb9283;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5bfb322599fd3af84367;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h624f58794d63e544a8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d9edb4bc512629c927c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4a0a87c9f64ec0734c16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a490c5b7782e730012b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c73d43a20e950ca12cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h145485d1150aed5c57fcd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he353d3378e09bad38eab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141e66d27148ec8a167e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h172b91757764b1744875f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8b268f0d76c3dbb242c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d45d7f1d88e9ee726995;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21070943c76715e7f500;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h639795763756be379421;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8c4954f1e01d9c361b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f1ac9fdc6d04fc60bdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee2cd993658826bc5eb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105bd62130a800bc3e650;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd996acfa43a87b298f83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha5e9e48a4b62f4118679;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7920425284ba4a2eff9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8682c1ba0366b314ce21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h723889dee49cfee7d95c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13dfd2a8e1011a394de7d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17888df29724b366ca18b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22100d4af18c29be9f93;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1948b49bae5bd3ca8e477;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h410f5065afa538fa53da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c66d5420b5d913a06ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d0be0118261237c8bfd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4849e63380cc12a606ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17135a6fb13af5883bb4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e4e3beb09d16d0a14ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12aff74608bcf93a3fdf5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3aef7c80fee86b634788;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd3c19ff35c40cb832a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1981027e0084523165676;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dfc3f958f4099d11ad7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f04b44a0d76b06050830;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15923de72ba83aa201698;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e325baf080e0c54fcf11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed5977ac838ca4d57438;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6d6d1d5a3da11d478d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11aa3cf90b3b96df7268;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c2798a82bcb2c83cd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ac2cf67591d670b5c58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8e5b5fc0516e396d352;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c18c3e20a2f588e333d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e619538c13a2e723e1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108ef224f9c81bffe1ee1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3bd72c1827295db1c42d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1617c9caa7c5f97ff9e15;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd052c51359d62242a1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f81a19978ab519681f2d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf3c6bc51d7f3a6a46cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h121d17f30076568fff9ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd0f627c79b80f9cc159;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9df2ce53681a526d64d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed91bcc1c9bb179f6ea6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h155042faaca54af7fcde1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1226c6e2b6779fcf4d998;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haca8b02883e4552a0445;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d19d4673a0385850c43d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19614f72289ef37f1d6df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8daa46474d80b4e7bd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aec5651409d511f37fd1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb69332cdd09de8ad3ac4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b75d4784d4716ac246b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57476a0083c136fd1e0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cea21ebe1fb2625e9863;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a683752e02f9eefdbce1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ddda19b5ae2a86ab4aa4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11914d5dea0751271f632;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac0ee8e475896c801592;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151b1959982e4b5d0e81b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114d6226a5c2b3fc824e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f1468c413cffac5cf293;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73a5bf9be9b77dad68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he44be65f8074122b4681;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160378383087940cf0ee6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112b13a8ff2b2264cefb0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c04e73a6f446d1145b08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8930325db4128476406;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hecd6ecf220c7fc739036;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcecdfe8a76de2e1afb4f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1736f37aced51fc12bc84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc8b142fc113daf6683c9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ea9b9fe5f697af1a06b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149339aab9fdcab2255de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e9249bc881f78b6ae49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31e457d788658467386;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152bc1ac2251795d662b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135119d862d0bc864c8fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23030fd5db04bd120986;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a08e56e77984c4ebbe0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b450d103eff91ca9a864;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a07a3d15ab668c0088d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad9bdb59f9c758825089;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h114c8429be4671288cba7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h737688284770ad355072;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h896eea2b28ca9bab5e39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1992cf3cb2d30603821a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e27c8977632211f81c38;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e181a9b1fa6f799b3148;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf908caab47fec8ea011;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1efb5f6fb853ed693e0b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h25b6f622e79c309d1b9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c8e9d7aa9f31b6cdbc5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1570bb918eeab45dfa65c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc78cb10d9b505daf586f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h978becc8237fcd8ce385;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ddc1231b4929c188939f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf046a40af535830b3498;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed4e8fd0bfcd6bc06e2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1929e9112054ea3629977;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha19c7337a2511a98536;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11aa290e2bca50e601b1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a07131fbadae70330d1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5dda0fcab1b1802a9dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c8b23a0664c92224973;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc1fc50d0dc167feb1ccc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a13d5f8b90063137312c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9f2f7b02c77fdd08de2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156691958ab5f99a3dd8f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11de31e9c28a8c62204e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b1a80e8e7d30f37dd0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0b9955bf67b5f73ecb3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc7cadae08af4bce7af52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c187b292c9c414bfad1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1459029fcd2044d7282ca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf5648c404b1d00e667a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17a47051f06b02f3fcf0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1994ee8abce242933aa73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1189e364f495ab591ae6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h510857768b6d1305eb9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc0ee7f81dfc03458ecb9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9ca0e5a45181e5a21f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h770960c7a050d5307a3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c439fe7e4e22e6adc581;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1412fbc5096b6ff9108e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e32b5b0fcdc00c2eea8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h48ddb430fda3d1623d7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d5f5069888456548495;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5bc26bba2afaecf662d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he5153ad4438d0444755d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c87872cdfbd772c95e18;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddecd2d8deb3227e8acf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13de97aa6e64e099f6e92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68c9d0742c6e7a67275b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17353f8b03e4cd934ca40;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5722e2937498933fb284;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb7d6f1344c7bef80997;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160470d82464ed4caaaf1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8b2791c2b3053cf1404;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1efde07e28de726e4ef9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b8ea69371d0e00abf12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h608a9630ae122bc69e63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3810bb0999b4ab91bfa0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc0f611b151f709b3e890;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he70df8b14732eadf654e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18851c089ec144aa64410;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he614fd74b33e4dd24afc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12367bd089e2712e8b24b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9c8b5c42c0b5122dedf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1304d2f598b58bd4fce76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef5c157d5474dfd43cce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7eab2aa6112687f1847c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42eb831f01d7554018ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h193bd33ba3bb3c1fc96a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf28a7b44f889f02c7a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc373053cf9f3a3ef849;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15fdee53514c505056132;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104ad7ee632c1bde2a622;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137ab65a497fe30989cca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9e2b8ce9902036fdc9b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b36dba7af2b6aa218a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10875dab0e18c7541c2c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5fcc8b21fe26563e34;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28612cde941bedf4842b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9da35e85fbcfe8e7a43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf1edb6a64874616d5e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f66f8b816d932b30e90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1809a1d33af2488d0b83f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149853d4a50bfcc7fcc24;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcaba1146c913b042a44e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h166da5a4a9541b81346a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1260a759460523d9b7134;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a43030ce6dcd5829d60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h78c0b269038fdce4470b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h375557b6c0a2afdd469e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e06da8b38c83f4417e60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2ef70fd0d6464e14eb46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104d7cf051461cc30491c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c1cd8833c73b3f7d5da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6218bd5cddb28fcad06d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198f7db23560db84f9d2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h303f7be40fbfee6673c9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1218bdb3cdab6ab31b37e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28d24018b14f24887579;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf9e8762ef0ed98900b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2893dcf51865fd9e3ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e67a3df33086a7602e72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16a696e2645b5cb73c373;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198fea0cda85a48c17b1e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18812d9bcac49602fcf1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151e41a9b2f1727286814;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb66357656bfb235c6723;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9a80c5fbaaf629f82dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc23076d7eb67b6d2010a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he35bf61335d04941b5fc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d9fe9fffe8f81b7db6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb96eb8570c3dcb4a2a20;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9238c16c52dee22f41c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf709e6c52120e1bd697f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha55995f99bd7e6e3f7a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc51ad0a4954d03f71ddc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8f69b958aa7d863cceb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h837a5e0bbbbfd0a25233;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf2c390d4c026b4e0b4a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd841f964167702bf942;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd153cd59aa64c5ce777e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bf5cd2704bd5df16f8e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d2b320577860b880c92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6df324c6a78a92743e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcbabfab05276e2be3e72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfdd2ea14070bcb82599e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12fd2f198f81d16b63ec7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f7000fdb11b367f2c86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2332d59a15b7d523df0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104ddb0d4893a1e11bcbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f6b2ff372d19ce8156b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e3f4464ade1adc3f4e9b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcdd073b4a148bbbad972;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0614d29a4be9cb61d2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138b7cec355d52eb6f115;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f6c5fcabaf162793066;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2d7afffca58a6d826;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd76ca2373c35fb03c949;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2289a33e04cbb2d28c81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h726ce5618b5f3372633;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b2c2a6aed44c3917040;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c8107c56dbcba88a1bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138de83627feab3433f42;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e3b67ecc0eacb6fd18f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186f74f5dc2769084cae4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb95215d93d80d53c747;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e69e2001fcb629ac151;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1651537c1122ee44c40a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h559850f3f9afa92b9c06;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1842db4da1bfc287847e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h173607de54353948ffa79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95e256fc31833cc9cad5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10991d9350bef2acbaa7b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ee300eb6e0bb63e93ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a7c3cbd8950284ac25c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92d4c44804913b5bf3dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3afd9e30aaf56e8eacb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53fd0851360bd714a428;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d2d1abfcc8a80ca1f5b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11664c8f1eb89a5b8a975;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a8696d1002a57f1246c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1520771c73fa127c647fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfda25ea9f2014dc300f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha99f91d9620d0b903f5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcdaf1db02166c4287196;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf53c20474a37e34ed24;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b3148b445018c8d4a23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he8702bcc7ccad3b0e086;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc59b30ab0680ccdcbfb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8c80f533547e33811ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1882526bbe4d32bddc268;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h214a6c8a0cb96d4983fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce1ee855dd9dfdfeff75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb82e5f35bc1cf08f857d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd67135b60bcbd31da7ca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb31fc69f5bde6d21b5da;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3a67a818ba5438d65c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39a2ac94d75f6b0f13bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cddc2b1b5d509ebdc9e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12beb0bd24bc8767efeb6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a3d30f9e31a396355e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31f15d4420c4988c7240;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc0a33badcd32ea99ed91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f679488bcec1b43e714;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he243a4cbe50e50ef98b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16072a4c79b146265dbb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87980251adeb34d713ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab9f96abfa10f2398acc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b25448e3d5fe8f3e0cc5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bdad1aace6e919bc6c64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9dfe08f06a3036c2b177;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf67b7244c2ac857f94fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38dd2767cc85305c649f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d9936626911aea3692f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47abbac03f42b72d7123;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h740399506fa8fe629ee5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c028e8b1a2c7a98e937;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h47f90cee841a32edb79b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a35b763da1517b8b867;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfeb7b40cf48c4a468549;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39a75ad78ed665d961e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h698d105223d929037cac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe3fbb496fcf89e38dc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b9b5ee9058fc22acccf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f9972147342630874b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1223d804136662f6728cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2a1d758c8b25e072912c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1448e682f9bbbc4c7eaa0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3dd844b8b5556114a777;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c37e3ef1d98aacfca1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57e1b88f0ffd82ae7a56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h43dcca4e4b343da47d67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10907fc7cfaaf398fe21b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5d13dc3194781a921a1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf73871cdda8ed3d36c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1afc2ee913ca539b2659c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68f6f1a7f1091a043dd5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc2ed0763d29113564113;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f25436bda7d24aa1d775;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12197677698e6a9a60c0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1484a8db246b94ecabfc5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c74758173e1d2cba7837;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a42e55ef3c6f67ff900e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d912f2c530b3e67f43b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e6ca380b8b3d67cc6fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2aa8c8858bd83be22f58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4beb7014d209bedfaa12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b4d2cee5534ed6d25e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f73678fa3f44367cb7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcad2e6103f5d676a4591;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc6cb63b6d7a732febe3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f4b1890681752375c8e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe5e161e046282257c27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d789454622ec6550d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c218ce59fc6bb2df99d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18acf0b8a943dd8531354;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103143983057abeeba8c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4edca3852e381c3cc2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159f22f4f38e4ba26d2e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdfb1a97afc413f5a4364;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h66877ea85e9756c516b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c0183dbab8abd756f7fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h770b4904863d91ee186e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fba144f633614af949a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h125486a3ef72cc2393e40;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14269999763b52977f7ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22ad6ee2f6c216764c51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f40dedc15d5fe464762;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1137949af3348987f01ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9ec5d5e5969f2381706;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113487f452c0c21e17386;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1901d88ac4fb51e13a12d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b890bd82ed4b77e532a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e5f111bb58e32f97cd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5c3a64cd84a6247c66b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19543ad217480eb5dfcb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1567228506ebdae6c618b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c13d17384a8fbd369a45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac1c8ee6f1a25055b1a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c431a006c188cd1d3faf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116d0dfdbbfd011892630;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca456cc96b4e8107ff04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc907e49baa7dfdc7fb85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10325a962cbe2840bac1e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d17dc3eb88402cc2900;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b2ce0e6a2e32786ddfb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12869c00d536bacb578be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb8b1d901b828f62ca93;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h101ed9a2f64b6a8f586d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1116a41e481d8ead8fa38;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4496927f4cfd2653477;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124237bf25feba1493fee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3b7bb3f51fa8d518ec2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11399c34461bf0e6fd549;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e64fa216a8d065562e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a5599615d2d11e0c0c2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e9e6a41dbcff93689e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d1cccd456efd0abdba66;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2fd2d6b5f55c6818812d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1471e6c818f5aacdbb224;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6576ba555db3412bc59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h425fc6de93d12e06065a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a67bd3c2a32f8de6b6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c45ab100c18d11247ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57e3e4826829be34c03e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf03db4edc93bd167c39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcd4d323d4ab4021900b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3387b67a27869b80608;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h534b11f05f206a6acce8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ff98208e06f616a971d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda6d42476f2b32a4a73e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117a547364a5c7b35c2b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc2bd3af4bf09cb94b601;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcdea21839a49e446fcec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d284830544f187e0f70;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ea1c2fb74d096c49f00;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hece94140bd10145bc9a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107424fb4e08e50a8640f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc8afa0386000a7655a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h134ad772eb6cc06d7ebb2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3e01c7c44e257b0a8cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2509bc1ee1eab8e9297;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hacf83a3ed96deb58284d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13dbd47a08c39056d7572;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59e221736daab216e3a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc70512c5631f107cf8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1efe4260cc574d32185c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2452103833f24f0b6696;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1412eff6943fd18ee8bbe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ac075d91c9b8c04c6df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h593ba599daeb3e7bf8ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d9f4e5ce351441cbcac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14869cb12d951042668e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf8e37dccd7d45df6307e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf0ca3a9e82576ad35bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1365b3014a9b55755ad1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac7ba6a597a223847863;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e3ffbbb2810b19a307;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69bd83c0ca9e096ab587;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb162a017c1094498e1f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ca5d37cf0cc0fe4af47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d1d94d027a433018507;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ff876ee3feff2ce25fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbdfbcbccd3a7a9214e97;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154a390fe613a9030e07b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h40e30e20d5b9ae11728d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15aa0e8169e2a0eac87b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1064461070173047176d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15961ffb2c4129e90f1ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18644738f60742ee55a0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h801ee66aa294bde48ff8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c9f18fd30d98c35d6249;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1900302a7b82a04d66519;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18fd7d7f370732b8ef2bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc004790991b80ab3c8f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f34acfa279fa32f944d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17cd5ffce32070e3ae405;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34aa2027faa3ba2d1c02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4941025e1eb7ec9d76f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3b6608f83c20345059c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9434a4aed7c20c8036ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f54931ec4c58b6c10fa4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b8cbd5106c86fe54800d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h180d95f68fa1e101df89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13392148a0528044a0020;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15190ffa900b1224d1c13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha89061be73d1e88cd1e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51651c90b78d0bc18471;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3bb1db0be507926bc86b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4949373967efdeeb6b05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18287c1a5142534e5a3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1191dac72721b91c67056;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h195d0b7f3c209328e0d75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h82dea75d01e882e46230;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1cef7d7c4019387e0f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he02626e4bcd2ba4db9cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6016b5396193834135c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1075ac4869d760dbf9893;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f10f348d095025f1371;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8104b4a4f4eb84d198;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba366cb226a122ba6708;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc9a12bd5e3849a06d6c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h735e47b41500e5e553b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ea7ce23a59032277203;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160d42b0638931ce598a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb13997dcd6ee35f27fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14f1d47663cb6d9e6f277;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1077ee3c0ad0666f9a9c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8df1ab4ad49fdbbc9549;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha244814e9301a87d1018;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1edf802061e7479ab6591;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc907c2c0d81333703574;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heea5308475fea0f33b27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h133d5ed75747b581d867b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127662688b9e38fd3cd7d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f770bd885411c028e714;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ee0f8e8d138733d9bdd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd3b153bbc0ff26612d08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f7a84c5dfb12ead8f6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c621f2cc99d44e9152c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2eac892ffaa3ca8e4226;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h48f0ac38cbbb17cc9c28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d8cb1da3215b6ccd181;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af7f6cd5c475986c6243;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f510a33d2df9026b361;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f8e5efc99448e7941d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dbe365dee66b0a6be845;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18a5ecf11da7eccf60ed8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2112d3acee2d700f2b71;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e3a1dca8c0f088207d1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102dd39d560af640cadcf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heeee68c1a095d53a28ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33f7db5693cdf7763a82;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af6c1e52c23d5a6dc113;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c164a0fb5499281d101;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d1092207d238b1710519;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he55df2937ce1968a3e76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2127fa6b7f82310ff452;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha36a4f7aa992592ec6d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108155403cd924c4524dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6820c41e50b54a309e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158c05eeb6f5140b2dbcd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158e6b1be4cbce864e829;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c59a949adc9f5c29071;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dfa522bb4ea264a09ab5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5023ee13bb020762e5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5a9788630a6428b7b73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d65813d0970b7e931470;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd452751c438fe5deea43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5397b292b3528530b5d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h35ede3d61d14f947d0f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c7185003aa48ce78c60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54776f161e2fb11818a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf61123c20f742f74fb6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18928f0673abb7dc5a27d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164a53c99297f594a59ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ebebfe4602cd2b5ed98c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119533a4e936a7a0395e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115f542f258a64b933930;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ca551b163f3480a6323;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h29ad2b602c3d64ae8dd0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b565c94996caba3a6ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ca003ddcaad62f56611;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd3db22cb3a32683febf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1651eccb46a5fbdf56c24;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6fe440db0abbc8d38ef7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9a486df51647f5633fb9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156094aef6faae82794c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7d3a6012f7da0b85636;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha173b62a8989314c13ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18852c4b950eef30fdde1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c69db2cd933380746d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176e0bdfd9cfe872ea91f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6fc99cb3be13db0cf28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13c3d99b8973e288e33f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ebf27baf8ef56f9de64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8e65343b36379d0a98f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc0d8ebf0dfcb0854467;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a5fc4f5a1f9de40028bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf868f760d7e93803ba85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec1e9fecbc8ea0bd3cd0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h138048374068f364fd19d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0a36fd8f404fe0954d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b826fb17f3041272f808;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b32f4d5732c8bc19829;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1742f61df601ab0911a57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d36e11de613169f547cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16005730f356ee4b69ecf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7cb99e291d3c6695507f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5f0f03fedd53a5e74837;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1205d087d09887084502a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13605caa4b393477dc284;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8c68318b7345259f271;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4224bddb0649e02b1ed2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf592a59e1a8a74ee7a31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c96a4038d21ead0e78c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175b2d41e19072ea228b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196ce4d43cff34ef0ff64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf8ef2590c88de387435;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b03049fc177717ba25e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19bd00ab95971deabaac7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c245cc27acbbb0e7a422;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2dedf8488700a5a0cb5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h111b8f791ed6a99066c32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf22e78f3266f7c056f96;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc8248ff542fa7964c7a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19cfc04959058706ae4c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf0ef2aac3e166ef7f3c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha56f5f3fcc5994824964;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h55163a266bce724c110a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d1f83cfbdeecd438ea5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53c97025253a3b9082f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae1d20761f6ca9c5bd32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7e612cc4cdadeb13b71d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60fadf25191e38e8c648;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d826459a9d1654935343;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199d34465f81cdc862ecf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88d4e23bc5a51b150727;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h682627c243fac3158960;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd69e7fc485b4d2307799;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5eac279145dc92b84cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1551fa546438e59784019;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f906f210f2b13255312;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb86cc7e573b527ccdbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa727be95592cac8e617;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6ecbff321bf22a1d6a02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19fb5b12242202a68997a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba73c511a1b163f75213;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12d5531f27645405b491f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd292c7fa6d13c6f6bd4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2152c3d8a38c7cd2c8f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1183fe89ef766945dd1cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23200c3f586f02f40625;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19012f7e90aa3da5ef8e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hccf8d047e3dc94a04be6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a543290938631a0a40c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5187119c0ffaac7fa44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d054d69ad798a5b8cf1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8dfe980051093e945ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e212f508da7b47e11617;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f3263fa2161d91985267;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e58cafcf13c40af20620;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16aee2d2f9b70ad9bb7b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11eff340177ab0cbf9977;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e55e60ab82ecdfeabe9d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h85c08c8613568c1a7c1d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67da0b7c1167dca83111;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d7478ffda4934d9dc0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1117a186e0ac1ee06a7ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b3009beb992a1970fed2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h275f1044d445750bd879;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36f06277131778921a33;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18510d38952f2a6aaa3c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fb65982ddd837f10c646;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7f887d588ff91bbeb95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h194e36a05cd45a8546848;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b1a41c2e1b65751f259;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5d84dbab20b52e26103;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2e8b045ba54979c192b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ecad4fd1c3d7f5c948a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7367b5dd81ea4a74e9ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbf539044fb952d7341eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72f154ca658390e53874;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5221874941f1855b49d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67c6d3eab0eda4555575;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h110429b5f60cf52c0d2a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9715f0e43224c15fcff3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c482d8caf21600624ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185738968738ccc9cba9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187f935110c604e77ba3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h521083757dfcf48166eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38213202e9daebdd393;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1996c1e6650e188ebab4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151e90c5bf248e8c7807a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7ecdc491ee20aeefb47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha6a2b9a6a2d5753a0f47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178671b79cbca0d42128f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38e8726b225bb0fd3660;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha560e7f81043499524a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he31a8c7510ae80cac4cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1affbca3ff5c13539818d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f18cc0b25bb21977ebba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16fec00bd4109ee4e303a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f3a9003c45380700a463;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92dff641f380f1a11dad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec0fea243f098ac85fcd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa8307a3d395b40ff339;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e201ec79bc3975321db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb05eafdd56ed77c6b15;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2a481df7ea598f53d7d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6045687a025cbfaa6930;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1406f924844648220f0f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16cdfef43ae182da71c08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1961b2df6e2b1797978f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc1e65da8d8049d5ab3e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf32098768893615d4a22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3e316397a54a289fc536;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52b704e14fd77a4e7177;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116d56c249d29d7701b31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d2994099278a386e772;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f5681290c12d23ef13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aff7a8623f57a1881633;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15bab3f64f805745b4256;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13967a59c11efcab9994f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de24d5bd24384bef8267;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc8a1e8fde79ef39f61c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1619229647cd302693376;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1446bdb481a2ddc156914;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a619233599393da9adc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea6f69b1990ab8a62068;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff6897a4ed7069c3eb8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h965481a566b855149f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12df1e69988edda396445;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1df7427acc02ade1650f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1673297306dc757d169;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa1b42eb69212216651e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae11a96539a7108e5354;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a531dc95121afea571f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192f5acbf39ecc8576c50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha61107ecbe94fe55f50f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b39ec44afcc7d9608196;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea7bac0ea741c4d51ce5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heab1f0daf0afcb42e5a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab2297a04b54c4ad6ba7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f67cf7fd62db78787a5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h408e8bd972c1f5525b80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b067d68559a033ef5e93;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h752e56c20d9e46ffe36d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6e85e564153dfbef18f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a4178b2bdd7e14a3e496;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34b3a15f25d3df239273;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1332f30e6dbc3c371be71;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b05d77b0f5d0539bd60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde62c4edddede8dd76bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9055a4e359e8dd17bd12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca5847c56a3130d274ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dbbf3a4cc56537449b91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a52f4deaaac978af37e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5e92d0a678792845e758;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1687cafb30eb02a3eac56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf152cec9571332f0169d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e380c22fd81588f49488;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c439a39ceaf66a90b05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8742b7e9c7c0437e427;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3e33262d2d20861734e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fb61f30447e52d6e35c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d2542066704fbb7bef6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7862e47981588c58c48;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33f8f68a989e37f1d394;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd0f80fc321e943364d8c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a5bc7aee53486af647;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10efc3dae1f80f911719b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h173ba94eef0d00377f88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e242efc6d6932bbc654f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c5684d738c4bbbc07a35;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h169a3e1be07f98cedc732;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h99501f31ad12f6ed3329;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae3bc09fe4193a8f3492;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a73eef15108e4780012;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f95755d23146ffb4763;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf87bf73beb6227517327;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9a64a69517cc3b97cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1576d10398b25748e08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa5b91c909ac5d4ce295;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3b6d78c24c635b56701c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5e23522126003330f462;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4930e68db81daee35913;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6a21e1d61895192b3a1;
        #1
        $finish();
    end
endmodule
