module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [27:0] src29;
    reg [26:0] src30;
    reg [25:0] src31;
    reg [24:0] src32;
    reg [23:0] src33;
    reg [22:0] src34;
    reg [21:0] src35;
    reg [20:0] src36;
    reg [19:0] src37;
    reg [18:0] src38;
    reg [17:0] src39;
    reg [16:0] src40;
    reg [15:0] src41;
    reg [14:0] src42;
    reg [13:0] src43;
    reg [12:0] src44;
    reg [11:0] src45;
    reg [10:0] src46;
    reg [9:0] src47;
    reg [8:0] src48;
    reg [7:0] src49;
    reg [6:0] src50;
    reg [5:0] src51;
    reg [4:0] src52;
    reg [3:0] src53;
    reg [2:0] src54;
    reg [1:0] src55;
    reg [0:0] src56;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [57:0] srcsum;
    wire [57:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3])<<53) + ((src54[0] + src54[1] + src54[2])<<54) + ((src55[0] + src55[1])<<55) + ((src56[0])<<56);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he31739dc8edd62fd506c1b827d44d8a1376c8c6f93449992b1d54fe1321ce7ffc50d751b92bdce378f56a42b909bda4ed73b7ecd7129d9b32a0e198623319bf51637a845219cb5a19ed66d8557d155738ea933a100fdce3f5cfcaa3ecdeb059eeccde6e4a733482675;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hae231ce80b1635d23e0aafb382f1ec238ac30f7930ad14a4417991a8ae78405df31ff80d3604e20d71a5da83346c86cc434aefe9f04818e1c0d89f74adb1fa885366466cb9052d8c49ea5eafc900b3e63504e7ce1841f0f8a4a42e81f493f87be8d6f0c523b9aadeb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168457ffd301276e4009934ebd085beba7445a938648067f1fa2af264c05939f0d1968cb936a0bf1da0980c3dfbbe9cc5782e236e3764bd24e3169168396bda47d9dfdfa9d2c8e5a16e1bf7c3a3c2064b1d0d958c18d07e3fbee3e6f2bfc0b033d21242cb75ad42e349;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d0c4d9235b97894f99759896ef6e345428b2c03dfdaf02d4fb121d8d34fca145fe632cf2963b67326c34b9da6d9434bdbc60751cfe0fefb4d735d56437e06e757573ff2868d74089e7a6e4b4c2e26b669b69b6c0998b504b178fe432852f4e994e17eda7b4d7790f99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8a8dcdd45a5f36b428cf6d938da2b58ef10621932e25a964c1e1cd0470aecdb48d4f56ecacc9bb4bc912c7a88f14a0d38acec499618c5c05ad4cdfc7d00fb85e96065c149c8d9b3a116a109f4a93e4cc79475170d6f9c7f73975cf1dfa7ccc5d6128a201a5f9664baf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h380b417040762ab1d822cf716d04ff41a3da312069f8a2553d14f1054f349ea355bc4395f7eb289070d2efc4d45820d77f838ebe631439f5a5c6d304cdac94f64f1b70687502ef818c861e3a5ab17bcabfbd68d0c10c6f4c8f022159288734ccb8518204a4eac33edc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he678c9f502d0638eff1266477a48110d903a1acabe53aff8ff810e0da92b748d2821e5d0f548f671d3e242bed2323f8934eee313c856d0fae4d1607fd38b162040d62d62e360c4c6847b1b0118843affd812eba8d8a1c7db0d547e907b87a6bfc61f61a5f583504b7b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c58438d01680b2d7187ec0a2b10094f451580ec695fd8d8d29a6f8b2471eb4e3f0f024c96c2dfe0eb4757ab2cbebf111756513e2445b050af6720a82e9d3dafde36e8dcea10f044a539bc583c4c5c07751f114fe57a4956706d2fc5baad275e72dbc4161193287740;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd97a017438d3a91e9d293c197095fe22c9dbae9a0cf121c0fe8e2794c4f3e22e270afcbc05a4a6251c5333f1301c1982cb41bfbc5d0d01f16c964bb32455a9da45734d72f736f76fd7b92ffe0b5bda6ab29daabf276020fc028c6f5b2b23b46291318d3de13350e8c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he769be76b3ee819c67407c41ec2848b62cd5d57f3e261d3665b01abd1da1dd18278d529544e4171e8096b8471db8588615287df1aabd2592b2ab672bb06628f874363f30984241523b2ff72d70adc3e6eba8c9e13a21c1bcb190650048bbbe03d1ac9d208aa309cfc5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99f36beb4136cff9cea7f1bbc311a7dd3661cd296257abad64af450d29aeaf28388a04a660e0a801b07d65e0078ee7a0585395064fdc2b6c368edb52cfde7339624daa4f93b664eb90cc1c574cd39b80269bb50b578f138048660f756c4beda5b9f4481f3908c5b89c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf83b379373fac78891cf4d5b87eb943d8bc138e628ca10895fb929a767324c55ae725f992ab7d96f72bae1fb16ae53691bc4ba6c64b7dd54b4b83a6515064aa86b470de6993eeea4f85fa9d8c46cf97e71fe4707ee19a781e6e7e41a42396b20ca16cc6416e5eabde;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b7acc71c198b722101cbadff2323cc888abe4bc2e6d049efb665925257361200a66713348ede623b8f53323c0cb880b138d577e08413b19c4c3d9f1ab4311b32549a69fb64e04ebafdc231142c893803f22686c5677f62a69380bd37ea4bc3368ba1d87f4f28fe2065;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc5aaf090ff52dd8b83c363c1c01dae702c7ff96248a3a1f14e6a51c910bbc3ec4493d31e7956818aafc84f4420ce4f578a68bf346055e91ab490b608f0ae287705507835ce6130ab7133a9c00baebf14a1cdc62f880f06cedecc68a88874226265d69765a8a6ba01f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4186afccf786c318e4509bb31c90ff638fbe62f2efc3f6ab46039c74d3636e32bd6363e1fb1dfd455286c217c0a6c41b6f8e9a1642322840ea80b5b885f269b45f0e3953430596eb0cfd667094c5c29c9b64baa343eca8bdd79e505a5221a6ac415459fbfd0e505caf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f0182db85669efa86db35f90f5f5a8514192cf8fc4e3efb63d5fd7693022ec6fde2887f0749be72c785c00386eae8226c81ca1bd21e9eb417e4c8e0d335ba791c7e09a6f3e6c5ab3f38a1b889b2fd80e877edab70d182278ba64bae15426032dbf4c67b098c72569a1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf26a2112ebe7a41a968d14d3ecda7445a1742f20dd72e0640cdb8a5b36b696932fd310728ccd7e13575a12e34d7f25c9fb54aabcb8417cb28dd0f5dcafc0e705963f8fe8461ec75ecbc5de63be4719b9497383ca359532cb7ff163eec5b21590507d6f6a3afc69043a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53f563261176f16fa0910217eaf50a5922eab5b48f3adc84b392bc7258c08dfc9b0390528192d8afdd1d3721c37139fea0d6a0364cca5c5bb60dd427b842915cb1c817e9ab7b68261ceecb8357b9f1ea9e779656b285c9047a89e33f9c8ed599492df533ed43b33f10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd722dea9a7099e52a4675a0cce8779198d2edae2ede6b2a547113cb4a5d889d4487c869cb8d50913e43addf83d2cecd0e97ec15e8a984d8590962b8e567212a5eac5dd26440f1960798c044a8a1836304a93633754c1decd1b531598a75cbd415e9b9f9d8cc31d8aba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a8e7b5b12503c5385b9eb4b14aca7716702ae3a4f098eaf87af96dd3b58bf0918c0fd16b2b79c51cd7be1ec633a9b76312edd623f1df6676f1486c20ff2093091f92700e648a7199a0a44dda2bf394f556317ed7835619a8d8eb606237c3dd04dae4ebd3384a9c4e2f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h150bf7bfe99d7f87d8e12d3599f97ffd1612ba22995f1d195a39b61f4ce87dbbee6e4db95f1e5fcee7fa2875c5e7f88d8f498a796fb1828e0495202748d453496ab01b399e07bd2707d62d8b63c796535c55f3262136055cf137c07b116cd6b5807fbfccb0c677f2f3c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15a07e1ba0e790bfa54da9a3c8cdb8e7689676eea8e080112497603b59be37eae001c4907665444f5d250ad7457e667078efc375cd7666ba781d8b55a482310e5f3365c6a237f99eb0684ec98608aeaf9bc636118078fecbe5df88d57fee055786c9b3c70d9086b9f84;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h796890cec836c57edcd05767ea8b783e26f5601a9c8a9f563ecc05a2d20703f65bc9acf4aabcf5d9123a1eee352736ce3be7650b3205bcb20a176dc4d8a1a8b075301326cfd63cf371ab7e28b7c48b4c628004912214a5e6f7ec0c4278050d789ba20c4d1c69665357;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h168423f2fa5be60feb91a81a411679f895f8ac17b415a003567498e6e399bd1c4da63310b263a5e3b770799fdf49e910e0622873fd15bc93584d40e49cb4942d420237813a0696453c9defbb2421b3ef145d27774d789896b1563d919eba4a51d07a7954aab4fbe7682;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h136ff8eda54cd3521ac89d6f708d1d04852c143fb74f79fd9214820073e50851057b54714a19a7b5fd205313f1871611b0c11f66ebd1903e313d282fd8b02f18239553e6850a9f4da6133d4666288541756a4cc7d533ecfc89b57667802b5e42cded92862f1700a7895;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100e8b392df77ed025d1ef1121dbd0d12bde41f9d693400f1ec124de31f42955f7cb2c9d3d42190d67e2354fe96604f959e8176be0d72e0046e0387db4968c9a4ac7ac4a0ef96c6c5560953089c642314ba16d5fc6a41ec17512a819f6a026a9e275161a6dd54ca56e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c46e3dbfe85afa4de3039cbee249544b9ee9667d2ccb805d3a2c4bbc744239bab0f33a638ae8a5a6b77ec5de612e3dca31acde8a8014da884abbd817a54c8671d7ead2ead37faa979628280d04ff72b032acc8ab30bc1e07f394bd9cbbbbfe13d2e63eaf23e20e4a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h186800212a8219d4d6bcba2b96995616e75cfb1f30139a2303cefd4f9a28a19d2ce5d819ac4e49b3595ad7941bb6705cfae9b4f22caa0f17b859418c9f5972b1af848e1a99a61330350ea964bd6761f5c256d01031fc7adc04fc1ff8683b605e40429ad44db9257c76c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b51d0962092fa0221cb4251e7dc136d75158a5b7d94e42f9475fb3ed29b6b0ae0e3c0a006712148d27ebdf54d3613bba3ce6d603f34d628e0fa779db1ebff84ba08a49e945ad2dd94964165c9419e9dd39c9a0ad9f0df0a91142d3d860dca443ae47c97a0a4a54b6fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h71e3739fa514261ecb679223589047b04fa5f3fb3ab738f3ee0375ce5a49e1cd1b5dfaa8a02b455b3c7e4121f7945313b9a8bf3ff4382147e5e267695d1cfb989ef5433b6b68e7a465a3d40a0d721d003de9d6267fad10d5555fb7f394554bfaf6e2a2378534b209d7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc8803468c4c509fbf6db985bc7a0a5c3c2c884bfa04ba2b1939717931e0706d9c25e05d29483ac097541ec3b05a387f9df01de9817b1b651afdc781b3e6d3e377cff6ea5b26d7fb723c9df27f17a8de438f2be5315c62031ed79a9612469f084b6088aeb6f4810e88;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h571aff4a54f27817122d68e12b8938e6e154b4d6ea23bed44c3b6253536a04b8dc4615b1033cc6ecbd693cf2dc66402ef471d2fd19af9cf57873f541b61f459f20e779e0e9a30404201c578c0fc65658f33c030b2057dfe0515bf7cfbc74406a427d03a0b98eac965f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a211eeaf80ece4aac4ca653e364fbb96bc96e2f49bab7eba5a528a04e5baed4d7a5f716c94b759e3173063fbf5a958777e421287f8fcb30d36ec2c919f6c936107fdcd5cc45ee8141563adf4e820aff35467a691f808551803fba9643c062376d1820ca8170e709f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2affd0d130ae1f8858306a3d9cc428c38b97b42292e80fc760a3cc83093b33cf28eb8aee172ed9e96cb611f6c8ee453a6d16088994efa80e60b19262ca8164237e5fafc8ea996f60f6b264f5a8c45e633ff7d87a1e2abeca01e28c44677169f08daed81fb8e3595cef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac5261d0078a4fd4291240d0533bd77d7051794fcba3850444044dce434e490e54cc16342abed32bd472ecf8b5fee835625d9042fa557385a3d12f7937c5b1701f0ed38af8fca2a15452814277188e660408b62a8c2166eaacf787a682fe0a64953f7bae13a0b7da5f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1db9517077d75583a8c161a2dc5006db8df980d005a5551d0baa3978bf338f1121b61d6dc9acf2a5a5428eca814886719aa2a0593267e6f51034270cd6ec6b3a7140e0b7f7ff5c8631a89133f8f9716a79d9d1d53b25a276ce74807cb9c1aa6ff499e5af415eded114f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1530335916191bfc1f6886b333ba819854ff7ba64ebfce7d412780f6f012c2ae15e61690d8ebfdb139dddad6f1a0373b93ae9455b6d60ac00b1176637684c3b1b0c88905ac6ec632ae1446ac1b04256ffae19c47755f80fb12c385b0759ab38600e88376e0937f9419b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d7f146a04dcb19c31de8c895fe312665bb3fd489fc2ecc4bc59eeef251bda6fb223af3eeb52676b89f1d435a81a9b525e477b4d1609698fe95c47819d83a87be8d2d1954ead4ad6e728f7b4e7260bd280aaa71daaf1615c7b4e10132303e6487400a7b5eae1201a56;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h103fd087fcd2e642ec6e6ae83c80c542d108fc85e8501c63f13797dc504b5873b6c2182947f36adbb3e00f90e9dfa2b5caa8413974865bcffb858f8e21035dbdd3d2f0086b4fb78b4ea1f04a43df160c978aab7792bf35196f94c35068185236ef2361b93b7b536ead5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2fc1dd1a8f9dc34100c37ec7e319c60b9d6053271c157850cee9f75956feb9635fdb5673d069486d824407e0b4e6fa59ce68569b46d76f30516ecac6e2fe4ba256fe96e2b8c89f32e6c9417a123ca40c7521e2fbdef94b804cced689f0ed228833e08d36492df7ae7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58e2925826b299732fcb0c96119d8b6915ba1952b5f861770403b7fb5e0de0861a3903f341af69dfef7a01a6a0c2e78e10ca2dc6c279f39085d3044633b906e414e5665e97105d39be3477d89ec6d5b42e1cc060e74ba644882b76fea53e9dd14d76034374ce3404b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af15f01b18fa2cebae3eaf1c651bc4b6a17414d9a034a739fcf870564cb3751201efc9cc4726327f76b1a7d25b0aeeac94d09e6365d4cd2037d4bd3dd89d11a65845a62db0a23305df47bf5bfc60e0ab712575ef1fe070bb91589658553ec5f7722665f3a257a24c50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13826abe2d03c298f3216a6b20721b90afffa3cfcdc9e37b354ec1bcabc522f569050993a4c8c695051c31cece591dccd3f29634c48829ef5741e584dbac1b0156cae717e336e3ff02de89f570b899f1579f11381af660345eed2b570a5cd6956697468b1a4c86c85c3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h487d42c37254e9a9b568b0f32d1e16b21c2fb836cf7d6140e112fcc55d5adaff4e632be6a37b97c56c989320dc58f7ba2c5a189be91ab8b2f084e96f2fe68794079dad63126dbe7c0d5434b1cef8ac5111215f70f94b0854c681bee5b4888884f679e52926ec04b682;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h88433cb6555e35974f8265bfffac06bf842306e1e138977f494ce6e7ffa05ca7ba881469375cc6890e16f9a33029ecf1d5029f867d5225785ec94545e228b2a37a2eab18e343b8f3db7f84666fcd46d4f1b38c4ca0a3cfe77776bbf84528880993d23a38476d951b87;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf032fd4d48be2741d52e23a9c9b125ee825d384328e1f878352b08d8c28362621aff594bd89264da80fafd608eb41a88264541488131ced41be89ad4110d9316db265581b4b244406b634edd0823e55c27574a89f559bd62d763e5a29d2d7520a548f9dd9549ed2674;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h52f5331d300c3f31deea5ebd84f1df33c1087a516ebf5264ae8ef52f2647bce34a93fa547ed9f48030193ff7d9430a7d1c53d58d23d7e612e580bbad15b7da12333744402f9ee1daecac25815e522d01b4fff958f8d5d037f3507d817a0e55984a130f12c01deab7a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0945c8e439601aafcfd302b82123778edd2d05aeb8e71f850698dbba8d2b5b95f6c1428d40d0fec0f83cfbf3c876294ed763d896736daba3345718db9f4400127ca34b7a94b036d70f15034fd0350c24c24fb8b0a05580656c45636a38bbab55e61a1996ee72a3be7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3f57d6aa71a675260bf475aaa8d635596db3e599f5fb51954f34245dab7b5e422537e1d7ef10514a6acd0333a1e9c0a920e2e9ff7115ecea981ab7df334167146314498ce2b707a39daef7ea827d6d5aed9fb0d9e46c3709f7cdd458eabc04c768e6fa55b84cb23b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h154c764ac8750da12563acdef84a9b1382abd79d3acd7c8bf68b4704fcd63894cf290d416a6f14ae0251d6637c4ddbcba22c1e0cb2e40a1c5e25e7f5fa8af03bd22c08f6d0cd511e4f830316f1d0e382544d67641151d82e2b9a464be0e16061ecab87110e748a88fac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2b39c83070205f6ba7045427cb64aecc1c639a617b95c95a250563c5fe6fb2485d1400ae9fd9053f22c11ddff103c604cab0e69bd5f6b3097d2b8a9694c34f59f04948103524654037cd8dd16ef950d7e87b502590a98d376c35bebb3c77e85ca26d03b56666adf318;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0644e3f5b0d9add6ea5749d95dfb9cc16dbe54fb130cc0950b47bcfd154a22d3953f15e9529318cd8982742e842b3c50d92f1d8f09d11e045ddde9a65c42456d0fcf91ec7e3b12080f5471aaf32d6ee6200444379f9f6f754b1629e098fc4f0adbea6125d4294f205;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6484d6fd566f4d3b022cde7869ea7752db41b4f9e62bdace6c8b143905a56e296df84103214c5d72ce2941e82ad7d6209db75708faff1a983e96989e69dacdd323f093e1030bf28cc8fa2810df3bcaf72d9b8ecd4295a6650df3d4c7a8c7d72354485791fe8a900d9f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2a5e4cf1a76b161bcd38a18b2e188b6f981e40938a26a100a218ebaf613e7e35bc4558b671e06d925d0de79f3dce8533a439f60390f74be1b560f3c6ea47c951675cf36630d1064b9a1ed0852b38852aaf3791369d68b7a280f9ff334ef45516e0f962b8fdd06b3ca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb2e4c5567a81c743cbb727984e6dbc1d357b1e4bab9b3ad7f3b727c62c5b42a54bb013a1f1a38d503647433bd29f2ff76b037a8c1ec4760f9548ffbcc8df24a1347f6e8a2b0e69f4aeb924148f24cfed82a3b94f221a39f8441a162d6f2d60922586901cd6821bbb55;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7b053cbf8ad21361bfc10d451d312e67a1d74b72bc5b5547b284f00ff0f0dae26b0c67017f42eff3e225a21f0b8f17a2aef33403c812ae4c72841eb6dead0c027ae9e0258e48d6bed16f5f4d94ffbdb37f63e7856fc3a45a0f7e315d5f6052ed9478302240cbffedf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f88fe443e43f3764b995b738e07f14d6011be07e6fafed03e8092a6886ad6ea113863ed96ecbdaf53725fca93851548289fbd2403f88253be80ce80f4e9cade6eaeb46ae79fe6170d82d6b50926621a960e0ac96ac5c599d335cd5baf1c2af72cb08882f0044a7444;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72240ec4d23dbf2e299f7d1b55b3092d928fed0e982a678a188db8c3765c4ed8f556d1d70c1873b865e6d99d40f5b60f0ce7e32c6e765e1845367df6856bb6091af766643c4edd80a2a766f45127867c4df325da18a36155e8518d9d2ea6b8394cfa2656d5aa0f699f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h141d2a78c14459b3d2f8e1f57a66dd6b126496e4ff3b1d2ac0f2450c8016027a1a5f62e60e3a81a608f3ca57c08cc5bab324a63f911733941d60ffab1a9eff80389b3c7715b2c050234418b55d481d19dfdcbf63507e2ea1081a9df3523a8196aec88c14a75e51777f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h105ea04013a82bd69c24627b7976a86ffe105a587d284a173771b0a09256699628f5bd5438a83adac2246658d7b2d11729fa85d4cc166c1652d7f384be87396a6a11eb6a36f0b2ed08f2651655a161da91ee9ef25174cac9898292956b06f382f24c2f0625ac53a939e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183f40da3e5f577214244f74bf1b4566f58f9786fac7528f865f83529f35469045fb5b4b40b6ad8840d28deca8fd9d7e55cce37caf617406c19e70cf28eff01d427a99be868fb2567e5974e4e1b4abaa22231aed1d83f850e5212e3afd2fc72e35ba173cdf8055d95c8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ac120c387a5da90669a10d5e14eb5a7bedc1c46d41fa2f529b928cc3256aca50fd7a6e43fd593b33fe74bd6874b051c0a0d9373bd60a0e76d9f954de1019a00b0dc58871a5189571359216e1d8ba6fa0a44f84a2f4d90d7b4c52e6788bc825bee96361e7370ae7337;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cd75650871c76c1b5f2060ad3b050283676ba28b929ba10f1f5b809db599a59187fa4b033cb24f892d5c4b0600fe64351380139abbc46817e4b655e0bff181c9e65c9391ce342f59aab6615f0a53ef8dad02b9b0d5909b5288f25ac4b2d9795e1c1bb3d0903029b004;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e7a723ec88364150992f689f10274fbe7d9870d5ecca261b8e63c1e35f512d2414cac2892198c1fd054e58b89e7231adf3ec21240e89ddd4827e4977a9a65bb5bec2d8fa2d7375cc83450606623ed3461ceb0005fba045c6bb4e16d2e2cbc4f9c5d19e871f66d7d4d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1add47e8ab97d05f370415fda2bbb5324a764e5df7892a8e00606339f58362f39bfd63e949144be6599b88b23e6c0d6e179b7c426dece396f89234a30c472f0691fc2dbe62827fd738d644114cf09302cdaaa72769d7b0a7795972eebaa030c484a7f8e2c4966a41210;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2edba752468249d1b7aa4039717eab0fdff6e908823f9787a14cec1877a533621ac40543d2c539c8cf82db0b408119200cae8b4d65161859d4d769433313bb4ec6f4e8b4ca3e3f48fa6a77b9a701846b3f6bdd3c0b90106d3ad75f595da4b47ad39f91b3b6e106b701;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h129728a412acd5ee711c8a9beebec256580bf8bebc1a650c120c8f5e324b298a22c8018f550b2ba92dca44d9860ad8eb01e37eede0cc72a6c3fbbf6b85d65910dada213844c6313bb514bb50cc2b4f24c57a1627ff361fbe7a8dc8120d1ba909a4d02767844c8b161ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f56f02743429fe34fa43ab181ea4a6cb005d4cde3c3cc1361a594cbb6ff3ae291e95325bfdd24eb954aa212bd2b4d8b4c7181aa1927d021f92d34e1e39463b00a5393a058eee7967b578db0ff0eb29da2d34ac69f05b2e97f55b179130fdbc241e0b34f5b232ae5428;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12a484636e4d560fd7c92f1dfa6dede3fa356701013c2911d03ce43bb8c92f43f7735ba7c11cf24e244bbad89044303560e1bcba5dce195612b08f116232171d6af49b3191740003819a9c9c444f222757e3766e97deba818938a5bee3714ebf36ff34601544412e58;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha69d91cb978afde469314346e627ef966ab6386cb08adff6896e238424c25cdb4803b25c76b79410cbe32ad933c6041e1d3348d90b84d5018eb2e54422f3f207b256d277234f840478306fbb4879330fcd697b05b67de3d3b87fdb540aa7a6587756f350c229016cda;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15b218f220c1c300b0ec6726cf74841cc87af4eb8a5c0acfa01fcfd0c114047105878d75f6da54dd9f5d6873db01f13fb95d85d075985610004a04ede47d0b00a05ba2fb6933367a8b067dc50d2cfe536f196a32b4f5e51b7e1b26d80c9f8101dcf123bda8db046db3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5376b4296d43ba0b0abaf683cc7e5f66631d14c00855500fcbb48c7040a1ca05fbaace48697b9a46abd47a7ccd1f8fdf8ecbf240085da0e3958cab06ae1ff0fe2ec5018e6247bc665594c6d1f84005f2ec751c9d990c2c6ef75cf7e81644a9bef2887d76da8acec872;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dba118e66e4bd2a500978e7f4677e027fd1009bda2d063e98b044d867bfebba1df794c405db0750a332866652c29c48864df985bee150c574c6f093ed33da150bd5788be9f58d020743cf7ac88829063aba63b7b8a6b3df2d347f5c813d3c314b2a8ebdce1fef9859b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169c37f5d9cf316ae91cec1025d49e5e1268eef116262b6edf87c2ec1f0ebb6c3938dc95bb16b3dcd51ce4f05c98737f5a33de3b8fb5d7031fe037ddf10cb7b4437a998d53f6bad8861813ddfeb0a082cb262d75cef378cbe63f77c0b310dd20c478cb664fde2bd313c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e95cc27beaa64b6b5e5bc6236a3b11847d9b00cff620ae2436ad264f098296100b9a98033a6389d03106b9bade00546e3fd7b7517f48ff8a26b2f400c20627dca4f9c2651d02e59ca2b9d870f0abe7e6cf712a7ee2267ecb1c37807afbdd45e1125a96fef17bb7a75a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdb1c7ce4d3115c32b4795f1254e8b2a545907df794715d9d9eaf56f19e33c73596273e33171c36c22ec7d53357db6ceb938f10ff1606b02d501c8c40f1cefe50f754c5e3c56dbbc5d96d009d60db7451a8c62a33d73ec60f849ab3366fee44173f0d740518b41e331;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ce3510ddcea36f4b068e43f6225fc1fa02d548cad58737978b4fa9602a3628a1d62758f9cf1f65e53da06bbe93f0504be1cebbc922101b26ce614f3ee4d371bd44ed6d97f779dc3851dfe9d97be1f6fc180b63d159080f42a44fb75a701a0c582c91be4ba4bbf5d7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133511491f67dd452401218a6d63363f1c88a5cd75694aa9895fd3f8ddafec8095790635106c5e8427c217547f0f945b881c2735f5f311c91b452ef7c8a5302d61574e8ab67cd7b3b8dff94b4b45d1e29a6b7264c087ab929294ae2808b05c67af812b4bea3d04c93b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c06d62970770e1fffe67996db19d979733530222335c55ca6b4cd32312ee8c43755561c12233b7cfa1ecb40f4731937869933fd5cab81fd312ce9f19f82d6a77e684878b9ccf11379501d910b27faa7e50660c2c4865eab7a5314ec5f3583e9df21e26bd231081e807;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73aa38e6cba027cde5586cff377a3ec8838aaf39604bfa0f6e2cf8e303134de5f3fe17e91da625c46f9bfa47b9ca531363ba8dc2e7d6730ebbb66385071f5ddc43708f096847a0435257e45945a858709c3ec9c7dfddbca222ef8bd29b2ee2f2f917170b09d7c60c0d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h178585128053f726d0dda4e60ada800cc496379fe4f30dd06de1860a04c0f0e2d804701b321d6b38d3d0ae2f1a02c54ef644da03800e70745dd6ffab8213e4b04787f185550ac08f0ecacd57c95fa343c18ee9da63f9a9065c4304d518c87c7fd575e192828152ed0eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h463006b0e18d87fd844e41722ad743bf7162eab9f39f847f41217e11ac4cc8779db9b4141635db5f0895454487e0c91c999538f35d8223919824fe82900100e44c1d3b945bc40a9dcdec80e98cd14c794e581e2d4659dfa70fd8d9b8f684ac0cc1797d83c48dcbede;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f26ae3373a67c2114dcc3668452543329392ff85e4476ce12e9216350c72f10f2e57c6f1c30b3af01336cfda52b2e3cb682f5077f404d4a4c4658f8d70cec833c9b5548181d32e439353161c40493d20a7fd99e29e8e197383174f472bb84f5b25b8173f2bcf3750ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af728529a97e127faf6d3f780d4802603cd20b49e24834f3301436fb167ea80810e72c39a565ab22b05712cec14f4bc17a920763e75b856e5031243e59e63054af6dbab21644823caf0d6e357268844a8cb944d5edfd3260bba5a3454bc7d7b8c7e1e440aacd9bed69;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2e7ea3b471380738d3f721ba16c9581cf4b8a8cc588dc983e2f6c65a491d8f6e1d51e821d9d73dfb2bbd3eebc2addec49ea1ea7e7f932e8a86739a202eac7a5ae54eb495a80075f06535f927d1efbccae38eed0c8dbf4b10dc2e3226288659dede5293e9eb71833a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40265192f70be94ae0bf805d244c65efe4c443fc82d02afd7035ea3f20dc6a77d0f27874da084011076e53fc6c855b191d678b9c42ecc2cfbada33c21255aa990c047331bc5afb3fdd8ace1ddf632335092c253c1ee252e8d1a09829404a2951305eb53afe54ab7a1f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5970c59d8ccd548493be6ab597ae2d512aac123be1def30e03d52ce9d39fabc2b1350bf457cb4417569469158235734efb502f3cc8b7b569864b01f14bda0a41e418f2d5cfdc06ff4cd9a6a7a7b24c54bcd770f88d6cf79d8b0588e7ca45bd64eda2aaea28c994b615;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf67dcf66f2ace3dbab7b389f6fd5eb158b423ec18cd6e3be9cdfe8c8eac381d366578076f97630f545c2436551dcddb04f0feb7675c2c12173bc2c97b9c4a57a4629b8ca48e253d3b89a45824f843784a20f08bec6f1c56085cec18391a9c65159a7d913a8c369e99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb55697f7a8edfd225ec69584816351603bf0273a3e8e8481614cd946270a40021457d157ec15b09f16b20c894ec8dd4e1262d70b06a6aadf593e94fc3cb8df707bbe50a3fe90bccd106e5132f3fa380e1dc4b195d5a133048606ff8a716d8bd30b4ef49dec47eec528;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1999aa80c83135ac384446298f2da1a79b002f1ed0f62d18c04d4097fd5b21a5024aad8c5ed1992f6a7b7b388bc5989f8c1aec92f43bb2b2c7707457f956f713c99318990d1cf48250d0ab4d836ecce9aba875c66885edf6dd4dce812beb00356019f3de9a2fa751cdd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8314a6b82b7011fb79e01cd0d009438f5e12718a0ed9c3bfc8bf0bc8ff483d43885751197fdec820220a832f08a3f2367f30b407ba0051aee81f29aa99811a4765c43e48b68929ff6f2fe845e111a23af9dd327b1338889b9ef09b4e88d0a48081bf264c6191440aaa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c6157727071b3ecfc0c6bc86b1afe616755dbdacef2430dcb85dfacf39b4a584f9975e7ec63e65294f7eaa9023827323ba0059fc052c99f1efed85ef43f74a4b91805c01f8f090e4ef3ae8129645d6b241a02f1b1afe6e61f2131ab83058ba98a18d6920dbbb974af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43fdab07947da9c3ffda7b1c62ecc42d1defa2acfc481536320d0be325268571557cd6a18ce67e57bb731596a0382f6bdc889447d9be999b0cb5594211d51dbef6f5dd1caac7ca2cd982cd3f5bd009355ddf7edae76733a99699a6852f9dc8f06fea00c85cc12d96fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc8730c414a0a6f5714144aa8e74bcee67602a78b499fd73bb003a51eb3c62834a268e866217abb09327b05063bb23451e606f73dc1213242351582e65e4df5ff82b4689499f1de4f7daa04f394c9db41551f8eaff7f04778fc4d36a72f5bcbc463c0148631ec73313c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fede9ff5dd560322a9dab3f66e06f7489b18da8e0b555bae5728a62f0837e1056b9b75a5ed93b8daac2caef90139b31697e35341e3d34ee8cd0abe5023a5cfd84ac820b3f81b7057c448c2aaf81e185fa63d5e7d022af14c5435e1a35ff15281b214efd30dfe5ad208;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e78aea4b83c705183558dc13b18efe4eb53f7715d19c3afabae42043582c0ee4ad72b6f0cbf284901d9c1ed71c574ba3e1c7e869287b27a213a872bd232b4f4b5abdab10011cf37eeb319bebdef5effb528c969f98de490d51e0663548065bc177075ed69e1ca10c9d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64a7a3e9654ac0437cc5d11524ef99ddc39e1c13f9187b89d642c2608d01559ef449240e8fa3a1c1aeb55c2177255f6678a554c799e35cb50dbd84de53b6c1476b8b4f5c9b0305cfbd1ba3071653445b9f53afdacc30fa301d4407130ff35f9ef943a31727fd04def6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf6960dc8a06531f2d630d2a3b99f17a585cc9f58aa264d98a7ef0ebe84b43161d287a90f07c066d84115e9e17cb3681efef9fb1500573c9ed28a6b9887f596f071d2894bbc9d8b1a259ebe3a881c2b70459ebf291b3aa3542ebce75c880b40aae7b42f0a649b63f391;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18958cb6e982e3197a7f152f72930b751277a9ee35917fe4cb03ad999a7b2cefb0a437df9be0d8b5ca30c584ca2d06c9322372f64e843bd2c6b508b8dd7b029673522e6be6e8b3b588f8a03132fdef7cbd0e37a7feca6d168e68267de8330974b3496ae7a203563ffb8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1545e19c0c850bf832858be4603e394890454445e562de007e36c82536361ffb9efe1ac3e2d980add8107bc41e3590eb1f9aca3cb85432d6098da45555c9d22c0ee5ac96acb973ee14e6ea3d0ada4d97fae1baca86183e6c082b493e9905c4c41a99aa757e743551242;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8216e250fe65455f5a7f184c16dc0ac52e8d9dffb6ab48d453d9f2c6a211ad52c1cb7d567ca871c2517e967a145abb1db8e43676aa9fc5548bd0ce1b61d05bb628558858fb515ddbe4a2ffb97c9d69dbe8d0eabe185c2416c257ef7e781ee606bf6bbcfbebc76be4c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28c514ea5d59be82436b1a2bc2f91f6202e87292ea446e78d4561efee410af71ada156d9b285be05039d7436aa76d7e21acaf934ab738ed96ea876e8840f669477d9304a0528b89e2f2a3278b37ca3a9b59a5161289ff83576d07f9a5417f8cf36e95938214bead42c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h489f75d3c84810ba5a4c4f6b6e4399b854f965e713db2c0016681541809a4d6f2bda5f30f7f6013c498b0cb3755868a12d64ccefe4dafcdf777c9cc5f010aa08c44043348e6c71a62dda061fff75c5c42ccbaa9596af5a847f16b070bb84a971509f28298b0d305514;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12da3ca6de8debe1b36776143499bad41048f940c31edce5fde930b551ac80484865873253ef61201235fed19fbc208cd45d87221962e57361c5ee0664a946842b8dd3ae61ecde5c25386f3bef1d1ee2adb408cb1e4b991d968214e683a83716bbb895e5bbc0738311c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ae73fba63b5b4234eeb889a17efaaddf7643016907c937b7bd13a58282ceeea5e53fd119e033850632610e17fc9f66bf74b9f96c60a015272083272aaa8d21d53fe21494673d2bab3cce24527f8d42f8af47dd3675a0623391c19c8680c41e2e1ce29728d2a08b33dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h843fa875972c4d76132bff2ec36a095c6e9488280b5d283c4cb6780b4bc59a7a8410e422bf1fe6936c45bf29aa4e537d7811aa1ffb04f46d89e79468ffcd2e2d4bcfc2c1c86b2ad2916df5e7a03a731e637e10c88628523067a2eed3c166782b38cce24e17cff41e71;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h74846a9bbb6f5783c3c0ff23408fb8d22db97d7a7987cc7051ea8b37cae21ba2873e05ee948aeda322b3b119b5aa287f10f552f0fc022175fd4dacc23662041d4206120daeae357dc415a0423cbe445e9142a848016bac458e055942afd24696c1db89317c776e604d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130a3c4ae8d5c9e4cda7616427564ade0ad25a05ade08125a74729f0f1996a1ac6d3cb6b3168f2c3033a92bdb4feed6c51e2817c6bb5dfd8032a1cef60f521acde715e4792e5eafc3277c5eccb8b773cf8ac632d9dd3bebdea1f12447857741124d830b0cf173001fbc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h30a11e9e2186bc6f3026e70514a344d0cb677744e03e516eb22c0c503925bdedf206c06b41d357a0b1a6c2b0860cbf8d0ba137371b932408d6327a96a72cf8e531a2c2e7bc9d93b6e8e923a7477a6665bd15acfece7b58b2db70c77732c4be602a3b7dd0dea88b6e68;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1322c993b564d6c3f9d72df22410443f0ccbf38e7a48a560110f6e6952a1713b0601e7286af928ebab89ecc0cee98abf9012c2c049f2305b975a9118174bff7ae209cdf733e3f0450d601511eb0373f59129001089ef8c5c930fe176ca14aee4bba82bef40c6c83f443;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h158a5a890d13d3b4de098eba83557b11d0262a2fa3e3f7f17f542b4a6789164ade7d885ccd8af19e650f9aadcf5cdd1dc33239a2212fc58e07b77765117c77863bd2130c9941bfea52a25e5202d9aba0dbcebc70f36538477916c8183df1054e3508ae6b207be0252bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d25f0317bb21bdd5a6fd16251e5049a3b543e72b765b22078cff810e1e500d5e9cb0cbb920c2493b88f69f992964c8655a887ebfca0e1a8878f6cb835b7742cb7255cccb711a6b23812ed4e838494e13c9f2a7c37bb2cb5803724467f26961b0eec1882297e1f08888;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h167772c11d3515e469dc958fb915c60a36239e906c81d33056c75d0bf47d7fe799de504c8330418efbadacdcf9c5e0f77fcae763988f8eb1bf3c9fc418d0ff2e0914fe3a813cb9191ea97facf1ce0cd579b11da3bf37649b6b958898c0cbca232218daea875ffdee8c8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dbbaeaf4b919dc30ac358c53d21557dbfca54f44e0d7605360d8f581400c7f69ab2128bad94f66b8c8bde970d39bda3e7f15534b46a2cf4cf31f0119024d4100cff63d0fc648654d0ca317d30be1cb546b7ce08591c1825c606711404df37ae843faab69382e895a4a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a421447e39ceac75df683be22de18240c8688a5af921bb36d97b0d166cc2d4db5f0757b708b5fd048babe8b4a3f7555572663221293ecb163c9e5bd5b6a6bc131f038a398c9228bcf8fea80d6b7ec798b85e6b67c29a71cbcacb98a9989399b56843c42db86d327cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b614b46c0a17d54a00c0a7ae138c9f85fd871bdee4b92666bb2228941096857ef6e399a10fc190b065202215a26c2d80798bdb9cc8c0637aebcd1f869c3707f3bffcc4d2dc95e5d1f838e812d400187a9226f70481f31a08321e049d0f1d16d536378aaa4b8b54a6bf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h366a286a135014481138e294e9cab4fa0632d8aee0b276963a1d910838e18aa39df728b0e8a27a512b23027e3ca48ef6450c93a6ecf6b8b2140a0f501d859d6f3b369201d9c1755e9d060567442721041efb9f10e7ecdf7988ba880f8ed07f0d116273fba5cf1f335a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ac05ffc091dc4cce365f54050651a914abf7433f9314675b50690aa456d4c8437ac2484658844e9018dbe6713037ed1d673080b30e42e5661de1078c2f17562c4941eb68b5769e0c61d7b50262207df8daa3c4320c4950877192b385b3a7fad2269ecc4a99760459b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e806aaf639ca3e2638f28674ec68ddcf5104c614cbfbcc7543a35e37d6a6fea58e0e344177a6e584dd025e80a455d01c6c7c7a683fc945f266e8b35502cf33dd079fbf592f78324acb4bab0390bed81b3d4480fc11de671af0ddf9bc9dd1c779dd7f9427994827c718;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21468842e825f72a9c18cf60b075ecbc245c62a0afa94d4253be6d100645356afaffbefc518e58c9994ab009bb2e232f2d97fd497a7f0cf49436a5e2fd137c77193559cc40333fd7e1df9cee636056b924b8edb87b92f3404c4ffa4450015f66af9b7824f1a1cd0513;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2afb07b4c40c28e2665c2d2efe5f93c05a7da15e3fd445f377f26b88adc6806408d861f5a6bfdf8ed8e9b6eab4916683830751e7e99e004b63281303d2df85d9598959a984844d335a5b81b28dfc19a2f92d8b870c193c459d6f2b02f63b6116695ad5e776b73577e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ef4566d65944ff8565c138e29c1e14ebc185afc1e2c51f067172b4232cc98539887af2d26c7f404a6ae1c665a3c4d1df0236385c380f3408bbac508aa50686e12bd37ba5083fa32de56be6b63138081e34cc8ed407aebf0bd64c298f33b14c8fa5a99bd341b69b7a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bbb211108ee12160de0f50e960446924489b2ec55d0cce596173fd22d8ef3dd2a3790702ea2c18002a205ef40cf0e5cc152063c3d74a4f1e075146eb85a64828a8d92425eb4536f2772a9d23b95dfe4414b8426cd44d1c3069df165a08e0212c8661755c69751c2641;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf857fc36ed052b039347eee6ddad721ba7e3095f745299907fe75d1c646576ad99557591171ed84e618b2a9f9578237ca8bf3c17bb73306017b707a85ca203472706f48596ded303bc1844d5f6cc965ad39f5a4d575e93317ee32538e2bf1c5d8c9831bccb99b0e2ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1273db587851b47bff40e13e1c2019b8b0d00df898fe11e344a1535911cfd50db270b14a95d296f38281ac96615928de41ab60ff7d970c28341b0417b279fe469bed41b1127581f8b6fc2c1a90a2ae7692990b4b656131f771c91e38e56222d1bb922e6cb69104b704d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c928631c448414ad759687a793d91fcd2ba0eae919df590f02279aa7949215d380dd42e3ebaf78a54fe5224012ac2e141f1267c6c7a3f39828321e4ee67d73f75baaeb0262de7c81031570593cbbac3b44a3cbf57e1d6f1ef5d34681c9157923db6a65d14f2a174bf8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea4e44c165c8c4b9a0575d04990431f104493bc776935ea8d27def99dc380e3306cc987583b1aab62e9f84e0982392282351a5cd70e62222e1e45c685ac48d9eadf4ea46ce08ca518088f42f64ab191ce92beb26cd2f73fa2bc670349de00db18f6b0d83a64159fdd8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6e80003f9a3621c65ddbcf7c5abab7811605c8dc6dcee6f2e283a210c1e9da196b3fa8116fa6ec5d7294f27ddece379215f4bc155043a55f62d1e3f92071ed9a2a4f17f2e16417558e358dcb00a4d06d371fd7935a86439b05bcb99fdd7e6097a903468386b8e4f65c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9cde418b916518c6a7a9a1d7fe1658022ec67c2c2338843bcdcb3383e4e329fc002794dda0044cf2ed534a367737bc36c263828e5e62f8a8b38f7c79df42aa5f7b98ecd1a52435f78f2c01be73af5004e60b734e08b23ba365c681fd835e3462af022e1051ff9fe4f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha9eb04e504fde8b4e534af75ffbebbb3ec95a4e2cbb9551e25ed70d4cfcc771ee2bc1cf7d6304cb40b9ca840329e21a0b5be2c7d3280984cb0f10344773dd0326ae78976c6d39c02cb344e8636e110b018c6b0bf50c62cb9da54c4ee8d1c6ee8136f200d9c71aca3eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16b95364b95f56e1327aea4ee9d2d862f9373e1975af0d667d62de310b041072d9a1021e84aa650e042f02e6e63eacbbfd1e6f5a4719ab998d97f8e561a70aa8ff0cc7f43c9602360f21e8f54a49e34ae53797692f386a270aa617a0325cb2c8ac0d0a2f00e71460fb8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h436c581320ef88ea7bbcfe1476313610b419883344a97175b4396939ffc13f6c0fc5eff76e00e28f2db85823459dd01fe276a6fe55d272108c810e7d7b6c7f968a23a6922b8161efef400b3092336b4d116f2a6a2818f7cc76ce63e1dec10bb668ea037535a5e4c197;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1347c3ec807a74f9ef4ed89659d62a10ec3dabd50b46f800f4295053c6b1f992d0d8c9948545232619a528259b4851e420450ed983dec9c43f31499b21d4c9672c577d84d53a4d3b4a341853462941383303c3bcabb77518bb869f5ec04545852993dd3183dd8d2db8a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15216407d03ae5d6c7addddb2406cbcf3b4b47e7085886ed399df7cebde7cea3e0144d1f83ac9d488c7f81797c1875d2cbae5bea0879524d2f9520bf4c21ff4a64303be02bfb6980a94e944dda0060a75f19b109f7fc6c9d767ab1c2225b78e5ad18a176510d59f35aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf0b6b394bd2f42f6e478ba08f3e89a96a759064ce313ee64ff2981f08c03907676e9a4dce07a7376770d0872cf4618ff92d89725a6eb61ea02da98940a9a98df3779549eaff63997961289b88f75d869fa9c7eab407fd7873b9d5d7913c2da4b33d8db65fb64677d2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haefe87ac6f48b71382be9243106ac74d7c1c10cdc11b76de644ee1a9cb975817a45957e225ecdf92a64ca14527e22938ce779803850decce73a6c9f212ff44671ab760b74d16e685971b681f2561f741f0c0348ffa02833f452046fc918f3c929d984d69ce3baed3d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3639e0bbfd1849fe8e8cb7c63f0dbf67fe754df35cdb9cd4da129f98cc489bab69963debc061fe4dc2341d736b516cb01ee3b86167f0f4eadc02915c52c08590a153a87e747159635fee2ceedda3495437c74e089e2d202e25e6db582d6d55afc4bd93cf3bed7813f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17452ee975bbcd21e47f5f2383da785b99c71af56aacd1c2d1b1a47aaca80eea1c13b99c408f3691573c93788c590b534e52a3d8b5b00fdd4dc44d893915752ce50ebc7269da89747b2986d78c501be6a37664acc17eeaee1fb3aa45c2f04ba70e7da556c902e39b22f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13dab60c8a2c1b7dbeabe4059d67b1b0e619b31c08789c0dd489444a51bbd681a1cf8a9801319568ba9622b088886d60a0558f5345e81c6c5fb952ad4cba031547a17bbdad88e1703f66960f1fd37479538e756068f0b7b569ac4c958c1989a45130f706302beffde6a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bb74449c6a16354e5f25b8b9fcf1c28a1647a020bcc91ca6c784305b4469ca517cd8a62bcb066c5994b667b1ac7ea5218b168fb481c7a689563f0418f206c9377c5c7f386ef298a368f6a7426b4c98294cb281ac9d415202f552c046d4175e9e8f1daa5dda42542c04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18331060a5d1340d363acc9185d583e2f44b3629c5665edcac756b02b99c5aca4704799fa1ce13da1c17cf53b6b2ddfaa627e0aceb6713fcc0c0382b0979937166ab840d9b746aa5abc629298d75d0a0ed84770545dd21f957a337649c4819114f715c931d346304504;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ccd18c382b0cd748e1e0bf37e9bb550cca7b94469d19ed14cf119c62a75fe08117f1e49bcac561aeaec7bf74f954e5f81e950d8f197e77c1f142ec9eb0fdfc37d8143a0a26729d85bf9f6dd0936ebf8a8ec1713bc3e6359713ee4254ab9759dc25a5a4289a601add90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ddcc22688af2f6159a793e943bf954de740150e66b3851cf4d16d987d6457a2f5aa1f21d93b14348963a460e79ae39627f9b808c360bcaabb3786bc9bb99bde9eab71d5acb1f2f694ffb7f3350e927b02edc5790e61249bb46ae4f12097fc9444c2149fa578507803;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4cc7f2ec7f711f6a436266df795b980f14a8efd5d87a0506a16510074b5825ab53dee1162baa8424ff2c93667f6cb481145d2dbe62660bbf24cdaafa731f1dfa8b3662ede28eef4d058e5a063c8acc947914f71983ec79640b6a115f1f16ecd60bd75423b94b5149b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17fa9f41e1fa5419197373f5af1fbb905761c30437d971a7d5806c9582a862865dec9781bb85052859b49be537db14cc545337afbeef67f197aad992ff380f020cf20d12b4b0ebd3c49a64c6132ea1a34fa0cb6159e63630e3c6bf349fa18b09948121839f18a7e9216;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3f8cc1ecc4e8062d5cea9dfce02232d8640a85a2f123a9ac7bd2ab0bf3dfad344f2b6a4834ebfa759f7c36a5f47826d456393bef939a5a48b46cadb19092392cc7e3471547b1ed700d26093e517184a228485a3c0f912975a604847b439ccea5eddd02f1c4cff234b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h90dc0e022180f8ca18d8d04e9cd9ed08f93b14304eae7488e8ced68674d8d87bdb05883cddba77b4e435663d9c17329592df0e6ed182ea1a8b934219d2fba6818a64541bf6b6265fae54b0edd2ffc81472ded685eea4a3bf4923f5fda670f9bc10f8a1ff656ebf0c47;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1005113387416461ab0e9519f7c00de40399da82cd376dc50aa1a9abeffb487ba5c3d46cae42f7874028300c61831ecef99d8c3767b149136412aea4116356e91dd50a13abb69b0f7cccb384ac63483d19df01b0321f6bc06fb22deb437db8890915ef855083d9e7d78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h188fcef70cc826d2a95f2f4f571e630a78dd084aa412394019100bea56492b746c5a009895d3576ecf44f4005c4b800af9b6f32b61d0ced138df6087fe47fd59a1597079a6f9b9a528ca3f9b28a9fad2ebbe7ee68ff95ed65361535ea4b40225b7e70390e9862ead82f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d41e31e3dc0f3b6163557c7de95d420b92969ad7ad09766816e990e9647fe6a16ec1189a42878e5d22f86c25c45f96920617661aaff65fe3a2097af675fca8184443a6acace9f7f058e148a702cc79cc8b89cb7dc30f73c07d37f344c94a120a5b2486ac70828f8f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4ea574379d28c299958c4ebb76b51d217650021a9d1b8e91828123f80ce52ee91dee44ae3442d2bdeb5d5cea5ae6267c3c98b9721863ef80232900f1732c777644042ed06886c4bc91aeb25478b3b887fc6634256a9e31087ca484b6164dedd3705dc48d114a589f90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5afdc9c1a6d783dd5ba364f9012f339716c79d6e7a6dc37ce85a03c681c99b436184e3f10078a680920ec79a51722682795b03d009594486454e649d0f007435493050018632bd955dd37305743bd038af3981811f3e34a4f89f25907cb4d7d448a0c4c90761f4e9b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1192df7f52c462da404e29e39053a885e2693927ac33a964ca2233e9bc89a2e97aecfe14d8c998bb0277e3bdfcd3aa75472b598aecffc057cb9d7b2a4fcb49c440900d3db0d338e838204a8dda2f0f8378c7460cf15e8e2a995f3ca88f4bc6ce85d1d44fabfebb1427a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h45ac75269045100df67c8e1a572fea51a5c7ce7a7ec71a53ba8038c4676d655352d59f45977e960d65e942a1b983b9a0980bef01462dd715461bf22873a2fdd9611627c1285a9687b2a91b2a81a80bfe532d3f3e988575fb4d0ca2541c2d71bf598ff4ff0616fe8a8b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11acf4189dd98aa27d99e803dd1de55667efb7008f14824b43558b917e721063a345c84f42ebdd2f8f84196e9724222aa4d1ac6df21636bf82a944d5c426fb343f0f1faecd1a082c35dbbd4f667d279a05c6a42d7ad2a5913c755dc9244574bf48446a76f8ee6ae7816;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc9464addb4b711f273f1e2d47bb0c91d69345577152b9293159a2ac29fe3f162cc9e3fe85bedcfbe705cfe3d8298992025be73ccf8c5abf55b3c5a68382d099ad240625c6a6f59a7ed4711795d8f9c5f81b658e87698904886fbde9e315e1579335e7273257e02d5b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2efbae8abf4dcf28ebfccbf4f63fe33b76dbeb5581dd1af29c137f4a39f5fb5333c96ebaaa1f637e7398875746795360b00ce6f0515b1ce549fc07e93c52f135925f54a8b36419f0e7f048a612a51a19fd1d3db521ef277e0b8b99a5e4ea3f595f758c29076e0f8409;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137e621dd584613c3a43d5a0482e75d41221291bf993980124a23cbc59e423fadf88cdec07681671b89f9b2922102cc2254d9abaff77b93485c7dc47d8d511b05d3f00f2c65d10b95b7a0b9e6ff183eea602d013731d3a5c288e582c9326a7fe9dcaf8eb12a35d14cc6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hefaa05d631b74283a86bf62735c9b0a9308c53ed666aabeab73336144b35fb383accdb20fbf60afc5d0de18155f64e77cb77298d01ab825d4336fd572a7591a2c2bf9c82e6313ccc9bb342ce083bc38035b3ddbe67dd7a8f3ea7b6c6b906b86df712c71a6a09dc50c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8bbcecb0c47a595b002799598d0bd1b5825beafa65ec36cff035ec0eb49a5ac76cc75cd810c7336159bc69d0ef0133e88b650ae689b2041e166d890e4528b02f8a1d15453e27e09a0d114b3174a85bea16de47a229b478f9f0bbbcbacbf313d8bf0facdf32e9420765;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h179c63d2ce5dbae807400b012173e94bf5859b8ff5ef56d9a5b545a07b246d6762ef583e2e404658c8ad703d95df27615d19ebd7491290523d8f0b514eda9d4ca64866c770e8fb0b48f02fc30e01416c2ce0049aa42890b7b48a96dca92f21ee692c8eb9e995322c147;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b2eef8f6808d8517726236b819e58b280407d5d4da9314c3a9f673e6243e40c3e61cf9a5af56031c38cdd97c94d99e033cf61e48f34f73d4b1deff107aa65abe17b13d900c293ee2ec238b6b51e9b1cd4e95ca99bec264bb316e6ead7c4eb6412a654ca5b71c661a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb6b51eb517bc5e5dacdb64b91db1c744d531fc2edd524fcfd1b5f894a7b0d21357c0a18bfb08ac066ab2843dcb303d22f10c6311daa38449af051abbcd74c598ee689d5643ef5edf1de1713867bad0c5ae4d8a0d916c2b6863e403c10c7ebd448229d3b8ebd463b35a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e280be6da3d340ed27be819b36e89dcb784714cc4fecac11e1ada72b94739ea40c34ef472e5aeeaafc09319afd367651f74817c5e26c55bada9a0fadbb3a988b5a9c6ff0c153209f9fe252e40ac925085f824fcae7bceb4da5fe2612f194a37a0f2d1fadf713e20136;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h958a734bc43d7cb19d1881e86f5f00b36f9986f95d96332ea2bf304db3f8926794c78ce94acf2985084a76da9625553a34ac507f1f07581383a174244da3d327d093caeb3e97b5800afd62578c071932d0de2ee99b33039a6a420d2ac553ea5cff8a4a7bc091a77b0c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7492bd8a45e8b17adf8be6e09e1c3e814c791330c4611059777377a3b1db09f5bdf32da42f0f504b2b5ec2e21f09543c7004a8ed0f77c4971f168ad2b76ea24dd412f445d4082358574499ce387775b4d139709aefdf4aab78ec6321a728c7a4540a37674d269d8201;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aa72baca6de0bbfa160dbf9f3ce436a908ded1105015e3de3e4eff3714d9059ccbe3bf3118af6e123c9cd7c9adcef323f98c2eab324c1dbb3cfeee4aca94173d5dbcc5d8a38f0b9970a03c384c5d266621de5d0ab66ea08d2fa8273716de3fb4f2e736c189a60387eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d7c28dddf5b5819c679012f8e297cad478e2aa1823fa0ce5aca46231d67e6e0cddb2199d9d23a947b658ab75741416bf2e3a0499926e53af540cd892f69a4d04fa51aa458b44069a7f53633a9b815669157c486c968be623a04e4a2ee12458f1998c8723003725fc5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcab952547c037e36b8ffac472c52476d3f06f797dcb9657093ec748816b847f382314e42a0570ed8d3509f16e61f424d9d18129b1659be3a5a890aee4f71d7d6d016c96f8fe8deb6a82db52ec13b16e1d80650b038e5d45e829c687c959d12dad1fb3a6239e4e4cc69;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb1ff8b7ea25ac01cf4109044d3abfae1619c64721554cfbe1dd238a597e14a541df06b05de0eb6c9f0c8a149aed7a1c51ef1e515d1fb362f36f0ac7616f8e2bdbd78fcee1cb23f33dc34751ece2d36f1b0e6630b2801bf5405b25b3d194fc05f0fedc3bfeef0fb285;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h655a5326687360582f8eb618bc1c4cfbc7b73cc47e6d4f7b5700979c6910a786ad2d40be5510a54d40890ff9da691091875d067d330757a285f5f514547ebeafff2ca869419f1834629f201331ce267d5dd17b5e4827c1bf7032f1fc847780ac732cd0262dc652daca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bd2c6bcce258a86687643ffd25236fc2e7767df62b7d37085d9db813bd7fb95bc05e692a232f06f010269899b02124b3265c3d1dce61317e7aa238ae1a0a47096aaf128a5eaf0e0561fbf7d8b3d88dadfd6753a53c6338160805a5ec3d3b3297f4847a35bd2167b60;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e808ee8eb1894eb72bbe314ae3ecd188336c7c69798064675c85a6be1af92a690125931e19a7b985ec8cf859c32ca6a89ca05e9526177c222a055fc22cde1318a904cb3c163a2e74f118a257f9bd697e175a2fe1806994a442ddc50f0635a802582ee1da7275ee678e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cb8cc2e3ea30d2d39cb1390920f1a0bc94b183a12bf544c3537261b7af0e1d8bf56c01378a55180a895c54d46434618402c6b9f48387d67da8b9a8e8d4588f5b1fdb17509e7351b73b75b637922e2b526682a71c1fc83647534640f8bcd829af3e2a0be52643f1738a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116fc3c7af8e83d1454a99fbf80817859f23ccf305487ff840803532de7b4e83764cc33e8da59418717b5e9757037de59a96ea0d95591533d6e415f0b3d5a0364183c6af823271b134a5228651845d64a4a03b942ca8b9c44ad87f78119f0e63028cb572ef7317f0ff6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6ea7e840d2ff30c97b7c91e5b5fdd242eb84f89f8534d3b88895164b1e9be4d5cfa4cc5a84b4bca9dd284592d5c8f247390d9a5812d85a278374faefc7a3c718da1f1701b17fe060293225b2b5cf8568827118e9bdc40a933ba351d96d3e9091b6e8f05fcd85ffea33;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h558e3c83ab504fb49a0da338b754dc47991e60e08960e5bb476933614e53f67925c3a5fb2574b3c1fcc59afc9dcf6a777a18816b6a8db0605280f78cb902ab49019c8fe13f47595906d4fa583b61239dbec5258f8049aea0c0b7241886b9e057c36db3b445f2d62eec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h714849cf0d546a4bca72b103d2f0fbdb4f5a37d2cbb919b264eda1383ff6b8329c4f603ace330818e0c1514e98f65be6467b262f602807c9f6d46b4708c3fc3bf079b18b43d0a2d8046cc1405abda80c1bd301a023b6662ca9141e818ef1897a988e91a806ec7fa85c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d2a356acfd5a40897da729eacd817c88409701b00a5a510d41fb0049777294cdd18406617dcc6e3a28f15069a7c748e7ea8614f7fa9df2dfd47ec45d7dbe042d552324b362e50b6db54258d406727c71b585bb2b38e88a182790c6d77c8421249b5eccb6a740c8effe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he79b1d7c06041bcc2c760e2a7b9c5c841887667e4acc3205b83996a9ec75d9e2c0dc1e44a460040536520d41f8ff9974eaa84e3b4904795109569041070679273a27751b0c9af0d81da37a92d4d3881c9a0d9247bbbee293f6f7aeb0d82bfe070b94fd08ab3d2267a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d54202f265b52a782d450d7cbca8810b64584e202f596971ba0d09363cca92874e84d0d704c49df9c77cfbe953da73820f720f7ab12f0bf891f7c7dce60261f65659fc38f2d3b890d414e6e32b5174acca556cca13fefd26aad9bcecee80ad3393da3a91f3d9ce7b0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bfc44265c7a7defe35c46f2a5736fe9709e078074f0ad57cb2b3987076f26563a9f55c705bcddcd7f89b141999a0c8cdd4aa7632452fa9c9b110d18f25abcbce9ed649a78d154493210de38938324b32b112f043801ec3cccb822f1fb993c122101254248ddd948639;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ff0206e2515b4a69750c02c37c743c58726350b0e6e0ae9668b5a3b1fbdc825a673eed1318255d4b5a727f2685201d54bb2c1733ab7376491f82ac7a2bb9ae511a39fd8f78d8e060f876d99c1702bfc5719a5a4d17739d560a229f32ac00884cadc498fb7ef94064c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54aac378e4c731d66aadc04e1a176bc11c5e3c4e46b2e5c49a695d71874c16fef3c50e76590f3238cee63f03b0bd8d01887caf970aab20e16f4d21ac6d03cc23fa067a056170906e25f891abb1bb830c2016d086c4fa65aea9ac0b6611509b5e77c96b0dfd0ece1b5c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbd40430f13c0b2a30eb2a2b1aac393216d83244921e5e5b64d12fd9cba0d7199a9f8c9d2007675af4930cacfc51bcf3c20a951c04198cf7819dcef41b55176bbb2075396982fffc800aff167bed868e75c69c3349655d8308394a80fd1ef4be5ffac4566a7ef9c880c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed4cd02df2c18d59c6579fd39b73eb08a6311a650ba333e9fa61d96466472f93fd3c9f01dbea64a2d39259306a48990edb4f85b651d3d9055993d69ede2065298545b3739e9177d71302d656be8acefb8aeb59bc3b930bb89f6d65edc8f29b3488d01ec128d93698f6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he558a5e9c2c36caf0e79e841cafd24386689d1711f5ab8d497f9f1b733c461d376f54b7bde2a65be74e3bb9a94515bf9d478c40eb75c127591f188f72aa983fc172c4f20d3695b49522228ca88edeb5f3ba7cf21455cef86de10c447bc9c6cb93b97ae210d82b06371;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f344c0fb9fab9cd80611a807cbcdd27cc1a8926469e6ac237611ccb1487041fe4df2d3d209c28ffb87ba02b2b581cc3d701edfa5fc058bf6448c894e78c1f93600fb3873c57f1bc11ff80603a87992361e29e9d6eae182a3f4461958391664bcdd6d2b0eb3f52c847;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb77c0d3a0323f9f177f230d253591c4cff4b0d27ca4d06f1ac05dfe1d6420efef8744438b0b6ea0f49a64aebdea2445656c9a38bdf761fae7d8b79ea4861d3e96d49ca5c408fa51876e43d181105f16390e946499da7d06d0bc1a9b443b12b8f47af56e601b0dc6ba1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c32d0300e67bba8eb0f073f896fa44d89f71c92fd6cf157cb180b6fb95ba9422abd9c0a95de50232734348b0f00004b2937a0cb693c9cf292c073b58c46f6558aa3b2a9342f261c588f9a5b906398c4e7fc070e7dac76bcef30e9624746c8ebcbad98fb2ba62606457;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65651902cd555c3f1fe733fbc0f6af9458067f0121a73ed56dc98090255d1243de02d282a25565df159230e84514b34f86ece55bd7782c5a2a3e08d72798ec1aeaf36d9cdce20029287e4968ceef83a47036db5a6fd580e3292d297b0d8a9422065376e29928730b4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125f11efaf296e58dbb65954e282c6190809d3f5025af7aaa104b95625bd720cc8b3d3dcb9ece44a49db926a7c023c72928484b55016538fb012786a7edc3016e40698da3c0d708d402cc65294b3d6fed7fa31b734beec43f8115254cc56e9122657a4a23f1b1cbfda1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28009104a928e39355b6b9c8cb77ba9866d6ea63993741c4a0af86019f582a8a6850ba6ef3c23ad191f268e0faefe9d5e0bba4d5ace3404474a10478c3a58ffed7fde35be6ed62d7869e0530c9d1a15c00a9989aee5c0333b701679eec9c557f7c23956c57c2415d2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb89760e9aa79fc978fc55ae9a5894209d54198f2fbb4f6241d4e52591ab2686edfee245a515e065582f7a4f07201d00996da1bb71a20537f9290dd2bc047982a523d1b5069efec15a0ac26849cf1477b0dc7a83b571bb54df3f9c2cba01f7f350f0eb6baca849242a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18207e6028d534da8c964fad6598688e55e34edb36a4da6838735171724375d98360d1d1e2106a4e8c26791bb3cc646f3d353a17f704315ceaa9f2d8e704b0c1f1be4b7ce1455c21f7d111ee562b075dc2dcedf492383e5da49256cd2482208521bc5686acc8dc169ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19214e784493e94502729e196e9b4cc79cd93ab5f05d367e7d854b4465f648c91b3f2d3adc4c12015a54aa35fdbe5d84a74ff1d455b9d9a312d281f5c5c327646f7c448aa1eea7387b5d793034c801cb13b7bfb42d995e1c47e38f530505a8d616d7e7cadeff9c6f49c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e4473bd7a8d635a542a602444a5525d2f9f3b3747c29be0391f0c831f1406afb3e5b884e261e4141c59d774f68ffe3ba2c92fe96a33c8435cb9e25c5b7cffd93ebfde769b58cf9ed6caded63cfc70ea2e798d4232852273cb70b362d14a18897ea5d1708c2325c0bba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47b73411b18b4e032c291391cd7e491b32f4f68aed04cd3a91d032847fff4e825370645b5748232eeb27ac98ca9d7ef812c88ec8263f67a18195633772baf7eac314cbc285e3a2648d8360f7548a70f27754a9ddf6f3e76d07222b841a7daad3fb6bae44bdf1ee4d28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd0636bb76f6eff3cba796c5ee488cf44860256c354ca00addf920da56150f56115fd7b90229cd5f08d6984faf11ad5948cfe85dec577cb2483a2a970d06f8526ad4388877bf90ccf18f15c462ad0e39d50de38784a827d702d32750759bb7a05667e96c3c1f6bf6a3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f1c9e3690581ffb6dd4756ac96c8e98666ebe09b94892d03537f81b9f222692d21f8ac3b47d4f158a956ffddfa27b63ec0937ec054799bfda6d2f8c89647f99ca04b04e50b5126e05cb12fbe331a05afcffe880b2180a716f18d0b557489c32814c5096a5b90187880;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h783b5e319c3b80a995baad2d2c0c3e47f4e099497381393c7d8ab1ef0b24e92a9035ed7efdd812730d17f4ddf431a25fe1db2a4a00e1fe6c01d729b55abc0d328097bf9c5c119648183b89d966f4edba965e2f0ed792d10a22605f1c8463748a084ad9f34556241d4e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bda54449db6b862c2dd0cedfba1d3e6336bc776f627e62c020459c47bf7ede6b686620e8b7eac5b4327f88aa0f33507d2e2a2a2e33b1f5ea2611b704f0101bd4a6a6bd11519c7dd7e27968b4de37c534090ed164ba9f81161b2b596be44f27dc6fe1d18714f05218bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf41e7c1e55b7a6bb6fd41bac5f40bff6aeea6c662a3a2643609e357dade903985c67dc4c312364ca1a8f0f31f884e1b56a87247849490aa85d2008202af21c0e0e8b096cde32925c3c3a82a2c2661454c0e3aea09a2a622229cd05fa691e7de9ab01a8b93277cc2cd1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18042b7ecbae1a856d60b4cdf3212655c0f91e01c568535917ec374c6b2411f8e4a4446887a6acc8ad84751f6c035eaadbbc78c76d3ddb11e992278168d313bd714fa83695234abd20af1d1778ec1d91138f21a3e85857724c956e87266b6233f2363c76f24b5d0f3b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbbe454a094dd295c7fb44f4813dd3a3e1ead0b43f8f1e7e582e8cc37bf2838963c687247c8fa0c8b97e2788e46dddddd48d720edb91838da48842325490b47bff9c50d0c2325d49a49c3ffdf2690fff4291c16d556fa9500936b042ca2051158c9e7ec45fe9410c162;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81e5edcff9a40d8d09e093d7738629f3ceecdbb63fb9eea5a9651bfbc3115b66a612eb1fc805c7caba408244cb6913dd81d7356fea734773ae19a14d5262b09cc177c8ca946d821f3655db794f45ad02f9ae95ab708ad8df1f9b1089e7bc53c657293f650f955a29ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf95a006a08318e0cefb689d5e9b2dff627e980f77d12f007b4a365a8953cf47e213de10dbb8524469672ee999487bf08d169b5059740b14339c40c293102d645d16390060db853df4ca19d9afb0464bfbbd7f81a69e684b2e4202b6d0000dab4e66606c6fbfb863a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1005410d1b97fa60b21a9b737f4a1ce36cef1df5db6c753f14b8e340f7fa493385203cbd39e0165e55595eb0dc2521df72eb15b93fca30cbed5879d0223719edbdfd6c7f434b212b1f771f3a1f6008625eaf61fd6b833aca8d74c790f2733ffc39b5200a221f626d41b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a697ee253fc98d246c25e368ab0f31237254163ba972199b3da5f4ed93ab516afcba8e63daf99e24ab99b77b0defd934f93cd6284ccde6e14b7f78862997c42a1cfda0dd1783566a6bc6d282de985006bccd29eceec7c18558137fedac69e34e96bbfda816143994a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h727235d8adad27859f0b8eda8784ab9fdb85b8af7888fb9af5c46fd96eaa212306781dbb3317fabe17de972ac20fbf9ded58c4239ec78c2fe392e8ece6ab7aeee29a9b8b426f2994b5022f3d2529ee91db9be3707b805f440ad13d569071a79b4427d2a0170cc6452d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31794f2140f6700ce8f163b7ce90de55622c79e24b4935e2f6e198b68eedb5d08880fcb2ac31c369f982a374b32ff4916fcbcebe4407697475879a2292dea979c6e36a746c43f2f77d34783efc4d689ed3269d40b63c737a7235a3a29ff0d34f8e614f3a2b9a1e259a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eee4aed4f81cc9136a4f70547402d1b9f6e9ddd8abe892dbfec34f98630b846f79e9ee4cf386a6d821d888c26c19d41d91df51c53f4c6c533292a8b4d91242d3394d22c83b5891a8834fda531bf8362d465044f6f6aa5cc65c2106407db624f8175c80ffdd17b98841;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3d11220574f169f1fdbbe3d20457ac82d1ccd4d05cecc2375fe00ac92192769ccd30478d398ae77452a8c92a7de27ba50b2f3b0fb0b24d0511f2ba513bae3c3ffacc10c7ee9bd95b7825d978bd46dcd359d31f3111f743addfa81f278a6f162bae42e7f7f7e1138246;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d984a8d94be40c10a9572a6a3e5c827bbfd0731580d965467ddc378197307e6eee52ba15c75270fb70eee79ba03a3b5da2bd908d553c0a80a0ae7e55a7e38509b244e5014badbf66392f805ed4c57e923642e5ab1d27906b65b95e91b33e2da24fa0a545ebd7b5cde;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7cca9a015f7130947c5b59a9147a22f949fea5dbf5e45a4bf93e7b5d0dc61dd07c7262862ce76f7236bd6146c4caa0fdcd8ba14a769063db58043cb08f54ee418e34f1ff6d4ae186685f3e8da3147bd5ebb2cc514ee357bc4cd7cb2ddf500ba1f32651178f1d30ac60;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ac7b67ed51e868598d18a31df81240aabe3801ba464c8e9c8b2baf354eabaaa45ca78edd2dd0a1757dbba3bcbe91a7a3127b28f93741097de0d23581655bd4f8ecb310b51cf2ce589a991e448be4853f81ed218cff3bd55c72a09fa002c1b81fb2839739c50d8daf4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1964d5aed013d680ba298955e4995badd184d1331a4ee0d7ee6e4ff899c947a6f77d580c7ee030cac06438f24051ec4631a580a09ff85c25468edc6885ab61f979d8adf3216e38e390fd6c443a6af534d2df193393bf850801558ec269d58812f73f8a7e21a011e4f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf9905d9e69bba3fad350bee2a61273fd11ff1a3023a9a313faf10694bb90f69187018a05af0ba611381e753df4e50e3611cec5582ff1a847651c291624ca711ab016c3609d08b91cdc84b7ad18b44f20b1aa24f99aeabd84ee619c49df2d0d1fd8d520df49e99ee99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2ffcbe8b6e86da4be629be0ed2194ba0b87b2c680e68a90ce24df8c4dc83835556c854a6e66e5591c3e38ccfa973ef46f347b62daa77865d999f4c55ad2fad2be5a6c1c193022b1006666f21f35ceefa9124ca381da2cabf2aa441596807881a0717a73ff61f728c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4db15d49dbefa7d1854cbff80761e5e0f5cce74530cee78652e2a1a7b7ec25c0bf3518d9c98c585f4932c965fb6397aa67b361925f850e72f08ed0d55d08362c34a104cdc3258e524204463804d31f348de2b50ffba678a3e68d7f613dd119b548e39dab4272ada7b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h78589783efda1991e4f370ac9cb8b74e4aea23f032046853078db6fb676389af85634172868a21bffdd2a2e969056ab50508b7211941c716e4fb5628b9f3662f6534ee77e27eb3a886006f83282e9f49aef4feda8285aef8e7c2e1de01e02d37ec2ad9ab61a2f4e61a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h142a872dfc1507927692c066c681daf6c46387186960cca090b2dc4da20b3681783d0e4e741e85e08e5d571cdfd69451386ec776b1fe20fea5aff6fd1e2e04932509dce34abf7ee889430ef52a9275348e9e07a60b73b52eb4bbbd8d00ebc0f3206987fb213196bfc34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14f64601440236d8906106621fa03e5975d4f1f34b1b1db5bb391e430437b8b292ebd0b1b797884a443f22d4cfd0c7a1f2cab4c9e46c7b8a6668656d2c27687d04acce7bd7f96c2b5f8935fd990f1b4aa1d35db279565b8335e210b10688975f14f34d17745bc3915e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hecd2769028bcd396aec1446a16dcfd2b68784cf532b891838e359a0b9a675a463f1822b7a5b00f90dffe202a4fc4bc52453b642914c30941542b72267ca58ec139ab9a567188ad55f97ff390d4272ac7f1dd0fb689cacb93b8a551f8bf23280da91b455a378684783e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7f53bb70cb58a43211313d60b9488e77972b55407f05dfbc1403ddfc3793857bec074b14677c5114881960ef87dcb40983d21cd6898eb560ba136b99132c3b9a6fac9f3397ad3f24b826d64b0460ba6f6dd5bbd33e649284db8613ac1759e2774b6cf290fba5441890;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h146b303e2b7d13634d9a8a0cb93641dfa9544307a70b5b4fb893a8a0c9bce6b4c1f709f5aa96a85e3eeca117ac7a96a6b4325bceb016b8c4967bca82ce5b944552734221c47ac405981b6ab81c8090bfa51cccd1b4bf8a9ff45aabe3ed4e5c08147c338a338e25ad685;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8a143238402a4182f9d3235f1c114ca61fa51e7cbcf7ff6c54872a11b74a8565af2cf85211e8855a5b5333d5b46890dc914f254b570ec9b79a82323fd776b530b5c948b6a29af5eeecb61d0ccb59af2c72746aebb91058b27b423c223a6e8f9d51e5b9fe68aabe44e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc761cffa774cb3f251317cb6b4506118147d09033c91e4931495e704988d688ad0cd41b27057ac78d4b0a7f9686fcbabf2595cdedc48aedd01ffff034540e190e241fe08860591c85fe60b349493399432dbf248c84414d3b80093911f16c280dc3cd87c3db4cbb727;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1adbcd6f363392bbc4e031595291f33c858ff6be1de1422c178dbd07a761f581e019491886e70f9f93f7c09fd8c3df6e61fda4373c39ec17184c4b7fd223d23eb86910bd63d864bfedbedd80a8290ea598a8e33780da43b1dcf77fe044644c51e3518c81fe03527accb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf737c7880dedd1876067785a2b5be99381d6dedcb8ebc3518a261e9c2f00ed4ee444e9806a33a22612ca52f5f29462eb1d2d007c880859f3c38b30c187f901db50b3c2d711f58a8f88e3b4954d4bc374bdf45414ac460c332e5e909a476917988d0c08547acd652690;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79359f46bbfa203aac7f1e6232470b02d719039294e062cbd2ac0243fa583284ba61f3c98ce12aa1063d8665961fed660df1327dc17eb7bc75677f5ebb541d0bd312186a4c98fd97c781bc45087213cbeafc62bf03f858bfa515890493f6eedb4bcc5ff8a872b21601;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a3491dcccf55c8945b272f2eeb118dad3b7071728b7947f54058a4149b35a5c4253a8e6e97b58c3fd88f899dec16f689b56ea885bba34daaabc0d269ef595bff05d1413452d43bb07d4f4247c2c85ccd567602a9f278bd986820ac99dccd76fb7aa7160b704810e76;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a3f5df13ca6a000eddee5bc530d593f5cb3f2793fb10cba06eb948079c17d82d19a49b6dca4537be524b60adad3f0863d5584c9d6a53b6f2471098e3dfa3103f91f6598bbb232005fd47a689867d3f700318c8cbf61062f8b14ef5e104703f1704fa375f7f35bdfe07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16175e529bb2daca13575974ceba9516b3a861dd8930b2210d6c63910bb3fc9c06870abc6ccc3241f2ddc58023b9ed7b8fd55c5a75befde79e7128e1f68ad149077883e5065e319986e5ab17f8bb435b67e38bed5bc01a7856c81dfa68399e333bcc30770c04c9f84ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c02d882baa10fd2fce745283b926a57bf302c40f48181c83ccb7d3e32b2640d30a159b23f5dc3d05bbe33f9be1c280211b6459fd0b616eb46d918a6b22f72d247127c56e5fc2a622439de1762bec23bbc543f5ffc6aa8e04f2604be66674583fc2e13361959875f4ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb8ce9b76581c75fa467406b44805ba911d127afaa74d0b26652815aa3cc534a96ab1246b2b87753eb371734e769010b8e58c283f664e3a214f0b94b7747db8cf25449e352083210ce47d7c6d9b292203aaf53bb40ad017ac2cc06268b9944da12d53f6ce1aead855e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h970c312c052ccbc433d2e32d3e884e44222a3bcaec656553c19d0830cb00d075173615ca26644b73d11af68f5d0d8d168ce0e32e672648b46e032e9a0b5a79000565c45818c59bb6a6dc8f6faf88a04e7b88ca68baf4e2ced9d986273638c0f8dca8c59a5adf0b905a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5d7e971de79310276a9bb6d831a4c0fa28da1c7d5845478c83898ed6d5b650542e24b468744eac7f0534a314065d89175e77efae7726ec4bb5361d2e30a9dfc3806684e7d2265fe47a50b7e1275e28bcebc62932632c09290bae89642357746b4dfc6e25bbe39b057c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1706f1f6540d65f854517d18a81f64eea65a701f5b4e4c20ee43943dc983e95970b80535fdc084f56a1c98140af23cdac54b70c4ad9a3634a7b6a2cfededc3289ce1870ad2e89b2b0e118262b3db174eb355bb2fb2287b7fc8ce6bc3b2d7dd42166da31d12e9008d7fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126926bdd2e24d63bd7e3655290a3b8d7447976098f375c74747abcda469394f81f8e03880908ebab463fe3d390c54b290ae7deb0f11c2173140815518eca99200f8ebc6806b2f91d0430492027282ca64aed79ac8bc6c16f07ebe085cb74d8c835369a5cb8f1eb05bb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18329c867ca94fdbd32bfb689c0b392b976a67af7c3fcc94db63b159202146ccb2d4029dd2c2280dcb84781b31063c0a34f5b30c3e42b590fa5248615f99227c6bda6f37997444af182a9e3cce5606fd1db331844dfae5eae4d9a3becd7e843028f451180dfecf98dff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h821e8561221ff936b81ce2ab3424b054a36bc2208f424fb7cb76e2a339c2e3577251faba913a202150efe4cf99996b1a88a4cc9064dda13b6640643c35d4e9144ce13e68d2fd4439ac9997bb40640da38babaf751020b60d64b12b633e5c822d59366b4849e5690726;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc3ecc5f7198674a7aff319bf77efedfb2840f2de407c53a5ae6b946bb661ac0e7d8d03eb6bd2e672b5590594e321f44c9ab223e5879832be14cde1a41f44c58abd355f31c5b778ac1688ba846e9befedf534818d8713c3bd0f729e9fad805d56404c2624c598303109;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17174d5921d1447adfdac70dbb9952036b48520f5ee37cf38393149dcbd48ddd549ba0c217416d222ec462f6f9adbe844651ddf42c626de3756d4b55de6adda721adb7d0a15eb62849e1f3e0d806e23f72441bff095f0e77efed6ccfbd8096dc3da71d454661b4df0cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5133a1f0ccac652207bc37d3c6f4a5a3e8ed98131813b6650d78a4a67b92db031403c4bfd2fba8ff06b46a8d3f2640d36df80cd5f7190e6d915fecee8acaed140813f2b3fa5ccaa4e9e216a56e6ed9859e4f8c51f7f0fcd52df23fc30567b2c84ec575b8d85983069;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h852460ce6b63cf6d39097f8d2a7a1aa6376ab7f8c1a9652465abb5aeb8002549cad2222758c0810e44514bb576e70f93bd7fc40943a01e051b0f78cc885b0e2df66c17513b15f41403cb01d2d28f9815064d8583a2df42f68f9f5718bbcf938d055a0ae172ad111fd1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h23be454f92c29d5818e33626c0bf229eb5a2649a00d3b66dac50baeed7724b6ce5dc1988d45b14151be54342d001238a62fc9b57f991059e21cf31c243559b9e15b51a43a7f0927113f34bd035cd018a9b9a4938fde49384aac3cafac0d6d13157ddb03ec6c543eba5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a1b827a34783928b7095e5298dd602806dd5adbcb85173651ee0a8fb8f7c7454f57998eefbc025d1b49ad58f62ef2055647e4afcbc4adcaebdcc656b896275801a5fa07a2d69eeadc0f580e533bde430c825d5028f93da43de4ee560955337c23dbe01ba720d1440e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1aeec66511a37dd9a26ddbcb49220b8d4b3a774c0dbb84a36927ee56f9c260d33333be62a134249f8d12b52c814c3a3f4286d685d516e3fd24a01b882ad690c9c8de65e3c2d08d38581764ac7247c371c8e64b2e8c1c1be8325d7cb392557916bc8ba80d12d39d4df18;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e41d27cfeb19c40950bb641a180cc76ce8a7148c8c056156566257b04748c2943b14675db979f6bf50285992e10906830771dd209fcfbd9209e57bf69d34f827b6f455f9030c833e716a821f77ca2fbc90f0d321bfafee8e170742115160cdfd881c8b6f7664667a57;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b86039130c4b614c44bc585339a72df99f10ede53f9dd6650af1794932026d30a7d1dc61830e023b1295a08e6deecf4d0bd875d67ec17a12a5773707db5e8218a4895d01dce8f45f89a3e33e6d7ed5b18ab57492596cdf67d3659ef452337d82bf75cfb869503afaa8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1265846830b62aac998b953059e287f4b4367866644ff38cc9042fd47b782a4ea99bf04dff04ddfece4bc3d403d30eab3ced24ded8fac41ddd1ddfb4fcf05f352fd0181f2677024c44d004457b92219812883e338ed993cdfdb13cdfed11a9e5a26cb54e111a23c7a7c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha3687bef09fbb2582540c91ed7527516bfaa103145a2474a92a6b09700b5c4b329e585f63588404c3c76bc4a643cb47e5df7b8d1b883777369309d7cd5abfa26cb3820602a0098c4cf1f73e3d7506b4be42b9702d51d1d4da8a5a86b73315fad3784ef16e01094599;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a556809a001870d9d86853c4cbda7f6904fe5b0323fe38352a452123ecb3d8991542c9ab082635eca4f09a41fd196459c3a3f68ba5b1ca0c63e96853c5d732b34e249e9b48bdb50120aa10a9d5a85bbd206ea2474320f9304cf5a8c4aaf4634de125e1f68a63ac899;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8a9a79f47dd74f7407793caa2ecc28c37927e022027dd15789b10ac684a199ac16834415a63962589aef1b7cf3f05bd613a6cad63e09b9d2c28269b5905b42198bdd63cb1d205ed860e3e0158d97da2fc57f873014c85810d1a26455cb3586a0ac9515c4e974fc45ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h591f7114c74489d9d841c4829f3df0e5b883a0dd2b74881831b74a3a3e18911a3fdca38f2e8078ab4e3225003e468a9254e286411f61e9ad46b9828d425a3b350a95df722590b17b4e8581a3c7986b0a57cd6112d7e0724df1849d224329a956185f8b4e59874296d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19dff3132d4f6bca685d76ba313f8296218dfbc0082a0dcc9cd20bd86dc1a50f6f2c2108e3ec22a91ec8f63b3274df74039585c24745c74c039b2a25e826154fe694d816cc9c275185aed7891263d495da9c2d529f68b431b781ee495a6b881bc19a29d77f7a8f63e9d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1190754397105673ecd2fddb6fad6b44cbc3ecf9953657512d74b331e236a2b4bb1df9dd2c348466f642d4fec248d4d01b599d6e248f956a1f29c421f1de2d4cdd16fa470e80b964af774d4d66c60de83329045b249ed4e86fee5af8744485968bcb379ff5022ab9918;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147f5d02b6b6115a243fc06a67573458d7d10af55669fbefd2cd783dc4e2c7271c49379f67c6a0513bfbd3befe9c8a22c0b09ed0c78cb422cbce24ad022cf1a45c0e7e3cf4a407d7a76a474d604e98d2b20476f2f603a77cc987326c2e190fa472db94896f780166bdd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13b4ac77def6c065960a7f3fd5487bdc227e5f66ab4461af5c8cccf4a3abd45d093afa412b810a702cda1fb612945d98384e51f0c074a3456bf42aa8c9729918db4583e2e84a650a3606366ffb4620a444952ea798c9d24d3f2829eee79dfc5ab31a04e462a639855a4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1121c537d4f46fa98380c47dcec60570f0d7d0e3e8aa5beb9850cb220a86fd18b03f76d0b1be027b64849d2a2242fd75f361a5e9e8b6db67de7a53cedc5c2efbef6730a687e2d7233472428e4c2a76f9a98113f36ff89bc8d0adc302c4025dd80f9bd2ee17c4b03032c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h178b45f94cd01bf36aa1e3cb9d0706db0c6f77d7103e1683c152326976530c0c86cee39227b6ac9e188dc5251e29ee8aa08c27376f1df9019d9ef953d393ac96573523576fb5973eabaa7f9e68d3a4db5596fdab3d85a63c7a6d89f1ba5f83ebcdfcad280448fcc7fc7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10267fee91dcba17500eb379b3d8cc929fdbe383e9c9476726d4ff1ad081473c9fde734808d9bf4f9309ccbf9304260a0bd7ae71a9f0afbe09176be9ab6cb89398db3ab73b7629d709d5bdd31f751cedaedfbb5bd9c55daec8d79c5bc2c9a4f988fcc13937187894d4d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4345b7968fd71542b435218c1ff5a5c2c70b1c985ae89e24b8f58f3845abe704f9e1cbbb4dd83342e24f5a2be4ed09efd8bc9729fe18dfac0fea33423ef687b50b875dff140d9f922a83df99fb3b09531b240e9667cfb05d151e8ec061eb99cfee92803a56cc3fec35;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2237271c10b24b6ea84bb37b4dcc39b0368c348111db5418204ec07137ff199bf8916963211b9a66523bd4868303823ae5c9637f0612f6abedb9f26b779519494337254fb422012281ef851c45057da1357545454d7bddf9ab04df6245c9640f00b135c84ac0d564d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ecd190f0a37c9436ac95b85bab0a08905555c6bf261a35d51f84b95dcecc338e59a95089915c2a60d371a355f4ed6ce7f55b7c4a35cd9b3ae29ab6ad942b3ca2caa3c78f9d0ce524357223c3d88e47a42893a09531b412298b6941bbc818aac97f6c0445258a4e59a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d739a5f25454ea5fa2ca960eab0851de1d2b1a0aa5f694ad0264ae25fdcf38279ef703c20a8744db12c698cf1ec7b77aee931156ec7d73b99d564e939c904d4e072b2157b669e8e7c65e4fdec76adf706a02ec7a7efd358c7bf0c9bba6c7511926a9e8900f90c75a74;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b475116c8b200b91607ea5fe1d4610b3f90c76bbd2d438a3594622a5959842a80aa59ff9b72ac9ed1c4ab035e4087a6635084f571e5f33f2d900c5287a925f00ccd4a7d852a12ecf1d28eeaacc47a8f9fbc8e5e02ae05e8beb707b597e474e50ae867240d6b34b04a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18d01baa403c9fba58ec4c26060cabcf91d8293daf84f4b67dc96b2bc2bbac586154ce3103307097794111c3be1a9c8af6759b0fa75ffbb04931393f1be0b06b3a0b77715aceb980f219e718222f3d680c55177ddfde76b095aba55a53593ac2740d0930879f60fc6b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17fa6788fbba8243841c83757f9d4cca7aff223bd437deb66751a7e8ec0094104d5e35fc4b7f078c4e3a579ad81a39de23d974eba7dd1e1d8763cdb10e91cf15e67d1ab2668c900061b0ad691c74d8dd8ed2c0f74759b900ee4fe970b5ca4a25faf459f62a866df8014;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18e1e94b0e086e3a8becc2e64e380fc7080c75ea1a9147a467c0239dd6c6f11a48239aed86b4eed9055d7075ed76efc2bb56faf7f119c04a818d77c93ac412a07b18d668c23379e7093161b5531ba30f340f5092e5c5d44bbaf2ffa86b1f0a64b0def88336ac9baf823;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a93e7d39e1cfe1d0b47a5aec185ec3a1b597fb24b7f62dc165cc249f2d06774bcac651ec9c07a4e0a7c774b8f0c08886b3f3d0a2cf591ce698046e7ed1c6030320121416e3267ca86443c0edc31a3f43cd0446ae5d7226671247c12bca9dcd66ab7a269e30a0cc6b55;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bd260d0a5d68013b0a58fb28495ff04ce3c3f93a2725e220a96fcd665526b5efac6c93da7540dab7532ddcd9d73e714e524fcb45fd76eb25f8e5f9d44cf55dcbffdc63bf412efcf3aaabcedd02f6c0f55e2034315fdb3ed1fe5405d12b1ed745af94f99d1f4f0e6807;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc3d3a32cd643bf0c22fce5c65488fc1b5002ace602aaa1a9cf7298a92524cdeb7a589a646ee4182375a0421614c849782648e82e5f3fb7c9776926c20d99268a665fdd4013c6be6ee4a36f1b7b055ef635838394683338aeabb70c5b5f48bfb7998aea134717606ea;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h484ce9cf448ae97faf011ab6be2b8346cda60b3df4bfd69ff496d880be9ada6a98e4f3728592f374e01896e7c8a01e28638aad0054d0705105d883d9fd64641cb99c99de53c000c12a272803b5f4af1dc2d1eb52450f66e09a61cca0e9ace0b764a04209d67a95c1ef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99e52e27cd773d8131b817042c9f9bee560ff4be3b67e859e553182f0a2cfb5761277d010879d7f9c2c99311137aeff32b48a82f9b6ff1fc0b4a417e4fdb62bd8fb955a31496c6eaab991e9e622090bbc827a3e10df5e136783a284c3605bb8ab7403978f640c28c5a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h116541a2e2002f15fce9ec1cc58ebc94f707bfc648995e0418a0959744fb94c625a7ace47291ecf9e0b2b5763fb6a4ef53dc4e9db9ac10b9e79f7d4c6286c836e5d1510650081db523b9fa0e025d8a70e4f804e08e62f09552a273fd3ad4e5e877bc3b89424897e4754;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa2bb158fe69341e57edb6c1da8321a7ee17374b69f380970a91f229e765c074a072876bedb2d1dab9f3bdbb63d190565ae9d18bc78c0077f8f46d5c78e4d0d965df181c6df2af5fb516029615f6fede72352a3a3547c4365fa31e09b5ef1f1d505b03bac3e55ca56d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163e73dfbb6f257ef90da396157444c09cb2850e1cc2e7206cce791e44d8982c2e678002d478b57d82b07ef495cc4cbe6a2ed0dad4c3231ee5aa26c3bfedd6e95f3998276215882d5dee74f96634663813e260fb8a7ef2ae557f7ac8c2dfbb5e3785033de4ced387f9f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9a69a76853ff906b4ac69fe8afd4a69c6bdbda8c637afbba87685f20bcf1960e1f07cef26b930c5779be8e7e362b8b70d33fe32878b596ebb9357b6705c1e803922848f8120819890af15061705ccf6f0ae8292a230763361ed05b1d3de876e2ce89e35f573074706;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d3f84fd9325c9e1228df0a30460df43b96af7255fdaaf02c8c80f6a7720364c272dae9dcef7a999cb017d3f9ce18a9f075c1f2f854f80c340d36f0824e13d896759bb1e2cc345021f6bffbdbf0fb957010b4763c3f3c4fce82268715ea0bc507959502c39d81f365e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ad249e77c04edf5eb12e0d2bd7cb5fe7a5c0c1b655268a7d083be94146753cf705fd14672bfea1940a8c82eac9294f98e9ba54c0208bdea5d065d86880d3006ff1d86c3102f401c48ebd4984f1815dbfe8e6930efd65f360a0bc09d5edf261a3f3bb32c8858a71c53f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c8a85fd313dc3c15ad004bbe88b8644b8975a61f32b9ef9a8dd381efcddf3676b290eb953aa5e021afa30116441a28cd64b913edf5d5aaa6b7c7144b39d03704a28580e357f93367a45f8783295a0c4f16ff0991b5431c77de4f77ed5388994116a6d5f5fc34b0d4c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf07e641ad89557bc1291c234fcc2ec5d250dfd0e2bb8ac7c75c48878485c3b2e39344e06094c9441e22f373ce92e0ee84624e7836e773c8c2f154aac9fe2123cd1b0c1ded62f2d72b13a081673e41943b47d4bd3e70c01a76e676be97de29302e8cb9498d6735cee6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h440046df6460c696e85a57f07a1259f6ba96038eedb701fe59b3b8aa6e71d54bef34cad49938f0ef898340f882d196b8076d97588e5a6c19469e2daaa6cb09fd3a7846b11428587aa4f4796cce1c6630ee61b3a9863b29942d019907f890d0ff6aad92337d24d86945;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c9d52b20073c62547b9a2cf24c3dbf0e98a39b487df1794ab07289d01698028bbb0169aeb0995aa613eabac2dd5996fb6306ce79d2afeaa2b661c3276a67da9297d36aec1a9f745242610296e24c8722fc090e92a5f95fd79c0af52e2f03f4af5bd9a1a09b4eca64e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c3ff4c077affcc6f591202e94520c08c41a2e1a03fd87aae8884b99fe5a6a18db44c45d6dde53cd43623d1c6c014a98b64f36561528122bb5945e267fbd45125831e07292e8a7eb68f5f9971a34d90d13e36c149601aaef97047f7d9171a084cd1e2034aba51d81de0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h639233056623daac15066c468c0ac85cd2c4b40ac14a755818644aa1277e511d8a2b23d263549ed04133dc5957d9c50aeb8bde1b6b42bcb04999447866c7cf9daf26aa021f1519bdff04d0191b80ad30d92467566b664e29dc1ddbc0b609bfbe90ad5fc637d0aa6c37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h339cb2f67359c083e100edcfd3b20ff005f9d93b9e1bbef976970fc0d6eda42cecf923b6bf38e3eef147c4d64e0ba7ea6244da0ce10a93dcdf90b97b1a76347c82ae19d66574536a4073e366856ed4505e6a0b8c541dd0144f2d723e157085427e14b2decf57161a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125d9b36eb3a467c745357726e8475465ae746531c693c7308c75c64297ad0e9842a8556accfdb212e0228f4807985142b552d8180756d0f1260ecd35ca7e23cd9f19d731c843a643ebac2f835815dc17034a4caef2d273f0f6f7e8383c0f9040843a0a1aad1125cab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11e05f1ce81df5e87047fbf1430e91be40d656c13382822b743921b45e1ce452b2ff639a21188435cc6f320913aef80b1ad7b50dc8efffdbad5acf9362af3df612f579ccdab9348d493f9b6d4243af950ea41d551e34a713ab3a91e8627aa398897bb65128ede6797e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8488cc2babe1e8195b80a223ffba85ed66f01962f3f2c585ff378d9893e098b6ee4bd9f9eaa7a340f6af11ccbce5ac66a515de667c9bd721a1c5a13ee46a60684fe2b79de730f6a09906acacb160fc60b8fbbec81ea217467df49a54b936301a7327ea85ef2e819cb0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130f896b5a231a6f78e7e082fa8848af7974b936a0ee9272d722213f6e5e328c290b7fa2de03deba0a23b26d6d44fa5e3f3bc4e756bf7a333c84540e8e1c3a441cfe7c7a3be9345124b692c725acc6087b0d4940d383c41ac9fab72101b6bf48e886a244339d60268e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133f17ecee3609642271255b4c298cff0d8cc4be211ee65b8f7fdda3442bcb25e929bc96f59b5a827b6e13d3a730a7c1c4bb8f881cef09f183ad8a55e65c8a3914bafe20a8445eabf390e0a271cf77fb291c68a609be761394575e6c662f366d0eca8c68d3bd22ddf3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h194ee53c682ff054e32d62959eac7f45b5bc33050b6138a30d948fa2277515d589beac4f035ea8c80fc77f5945665108befbc480a3734df6135c1a5bb53ca4c8c657f162d8499a21b3c1313f7558dde2d7287838aa7aa46c56e9190f33dd493c02915678c30dc588e73;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h510c0cb1b64dab071f91492a8a59ae8818abbb1e23dbfb7f1c0a4d750caf65d66f96f35f426848006f9cfb80c486c1ab214c355f7bf4694b4fd1ecd270e9d78a18fbf0fc1c657cb945fc7d3883329d771bca39a5392a52cc22c8fb2cd009098dc1c9e32077c298e576;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1078da62a72ec96eb853e002c5f28f8c8de549c82f5385daf37128f6d7e7c1d707df4658b885a2a36890c19fd6b1fe41dc7aaf430c4f02d266cef1a0992fed68345987054f8d5c13b43a1a5be46d056727d9e324699a624ddbb897bb535cfab3cc7ad7f0b5ebf1d79;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e663b3919a5cc2f4e27b1535bde39e050eefe11f66fe02d290c08db4083bba6a395ca1414aa39736f47da5a109bf9b9dd27323a7a2b18a08df6593afc97583c931c2172e140d40de3d6b1c3fe8303d6b47627087db520faa86fa1bbc3576f74e3997a2415da70a08f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99716f8049bb8055b248a20fc6f4cbf40aae1642dba50d57e849eb78502fae8da470901964d50a425c4d5faef056f67c765ee22c0b52a3fdd0450f5d97128500d2c4e0e8ac4eb56d959cfefbaa953817a20e77a1ddaa9a442ff34b25ec7920a2253b0ecccbaa4acb58;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152e8a60ad464c2755c8c0dd4bb03ccfd07996d8a3af31f233494e8bf325390f7a4b8fe6995ca319900869583224714e34b55caebd2d092a53354bb0a49c1a8a22abc02a6773c6a2356b9c96dc26cabe62f6dcaa9c1186d8e6fe719adec3770e2d9172beec0bb2a7fad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h95e68df9aacb8a2401a3ed968dc067cf326ac34b751e9f475b5f42aa81378ccf7b0c48eb1b9f1b8fe1605b1e816e15b0f9d311d8e36c82245702bdb92e0fad0cd203baa074ecebd3f9c08f0ae22213a15a04581ee217326b865f7fa5d0769d20025a534fd86ae5dd42;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9354e4e9da8741dd7335044b74f229aa39b92904327455f4ab040ca5051201443625086c4cb578019067a20a9ab57f936c0e3f2cbd7a34499b8d4c3b6553390b1980153d61682c0db1b339b8bd97dea5927d670ea3f52b47f18fe2c1b025783f5231673a173e46d29;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1728415ee41e39a9bc70f1b609c88f0e41aec0973a0377fb267dae93177cefbff36136ee6556eab79c69fd7d0ee9a42c05d4f4726bf34bc79bb1243ca413d986cc91d93ca315b98a22f48e8e256053c12f2e186b06044c3e79639b5d99e401b45cf80abeeb994046c05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1185b0e84fe05849c64d72b4b184c45c750f24d87aac3b5b153ebccf9d87b1abe2f7e65c3aaeddd4b9cbbc6719b364a5c875fab8de785c78f7918c62e1d64c8ec8fb992c0bced5f6c86b0cc4d865f69a7bb3eec981cbef22db427bd7769ba03d65551bd71c6efedf65b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b254a1ea7fa70275c4a32670cd4cbc2789794f87d2a9e4fd87e5306101d31e2a4040a7164b5be5576ab31d13c8938e950f2076d37ec58191cebf5e6a09d078597a3e9a891fa74b8b6462c211cd2ec1e9dd693d13a63a7f9ff2d1c4aec71d996f3097c61e311c08ed36;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbdaec6fa8616fbd1af9141b7958c74eaa7db7f60eba00bd1b44d914deb28b360dbe6713a88f2acfeed9633bba5235d3ec3af75d7437816b8d597d2e4dae028a4b65a84a64df56b083d511427a35ee9d51d3987fa34db5d62b4b120f742743f4aa755b8a8da40d40d97;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b72d46fa1729f01c2586f05fa01be7ebb34e38a2b84a37f9dcd818e802b65b53a521dfd71becd9d9c80fc93beb911b26d59f756c56dbbe37ae2333b64a336432856c35ac49a07196b4ca3e81eb1089e050d823fd2f55234d95d9f9e07f4fded1ee93e2e17f2714ae24;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19cb6d307d89cad74bc31038ef52640c228912df9927488b1d576a9db7082fd29e583d11c801924d07b9ccf5ee97708d5c54528b5cb4e53c18f29613bd18c6299bc0b44d3f45866014424e2ac9b13184c481eadd5473555eed832ef4478d42f4687564412a2f529a83c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h149ce563f418e071aaa2a4b4f3ec5f25c92d879126eb75a6691f5414a54f36d39b69738b7fcdb74f4d90ef951f767f289c722bd79a9a89bb0b104909709cdb9330a310374b34769097520a8c044e4c7aaa58577a7e791850be454dfe417e816eb094bd737649b4c713c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16de7239c17b6b77c4c5c7f4ffba278002d16b6280ae1888932a1412bdb85c749c540cb389a11d1276c306e43aed988766d32fc540eedc4f1db9f93074546361e8b3e4f31336605b8957dac91ecb014f6364abde6cec218c53b4a6b412e9abedac0f8bbdae16a2bd8bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h418dff01cd86564d8d15b63e9cc87cb169afae378163fe0f11acdf16bacc441993f0ac0854810123849c2da72f08f96f97f42c48fe7e3c2ca3e70069499fb7f6102586306b97efcf0d858d4d0cd73af887ada42d973215ac897e30f536e483f7f9563afa74df2bdd30;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1674db1668803a6e3fe85f5945a0058dc4cdb4bb51b8f84330b7431f1045f6edab09ce55458c6aa9ea855bc1cab7a81b554e1f6690e2d6ba56d4af469df2f903c0951aabd84b40a7ee8f40e75b719336fb5d5bd6e44ced3be15e0728d2bfe0181efce2ba8b845068e93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161e3c792d8df1ed63c8042e12a5fcd1e1614db43a42553c04978f11aa2fc49799c978647dfd8ac27c6bb701659d9c7ce179d8504de3bfc74d882a937a1e14f14be038e3c7da60ea018c646cf5d8dfe170f7ad46d16023b285457e0abb0af90d1ed34885344c68819d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h145cf4b7db74c873221ce072bc4fc9039847956eaa2ea7b6dd44510b4764cd831a7a05a1d116aa35aa00c8011bf7b7aa4f48683bd45b78aecd1e16541d1c6467a4fe994a623c0452f27c6f2475d795e2cce4457d15f78c4379040f7fd34db69d09c6d17436fd1f24e95;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108a556e60f1704173e137ce7b4ac10040b0d2118b47bae49bd9ec491d11eb7b682f9c3d8c5820ce36a4a0ac27510b388a6790895dfdca1601384e02bbce000cae33d5e00d3e97b356674d08267acbe06c53ec1945472c9f8e0405d048839d76fd7a26c19d8f098338;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79ef2b96b081cd1a6a4e7edae3347cd1892ee44187901fa3c968f564d8673ecfdd3d0062c71d024064c23f7a732dd0954fa8eac00a69a997af8475c8aa409bb8735b0132e1752384e8e27c741d73cb2eed628bce5e8278d2f5d4bfca23fe8b89a0e7667e6251d91b6d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h653131f76a3d5ee74065cff1595c492931ab3fe017fc59ef4b8bb9bcde40ee837515b939ce84490fc890832c6fab1384208280442a48da475db7239bf7dd221db546cd567e74947c16620b62ab380252507df000f9cd8620ac214d160a8472f556868148d4c830ecb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1104a5a47fe1c103fa9c79f44a4b53e73d62cbb48eec45360b2ccd8b6e58b313c8f32829f96c1143cd55116bcd961afed7230293fffe4b9b4269360b8b0d2d93ca31f31830f44c81f69f4165f56cb8c6cb39779567ad36f63ee6200c31ab4497cd63eb48e2245bc1ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf90a2c532f4b846bd9fbe3be6c400b929112dadd58f6743e2aff560f8ba5a1a61b0d1fb613a3642e3bdad9ed4b2b2d04024ab3f1c50b9c7f26af31cff5801f36a001b1fad600d0811400a6333378a7684510fa844e9fbab701031eec10c4415d1eb2150e44e96a1fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18fd299e8923c8ba15d922c670ae237dd37261254dd798d074793368822ef389f3dd56a1b68497137e4e378e2752fcb0babda9a0e7b60add3efaf0bc49f21d35e53b8e5ca32e286e944e758203dc0b72116cf9a6b800100dcb3ed3447ea5cabcf46fef990fe5ec798e0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d81bb20e9b6618cc54a9336d910421969b82525b2385be11619b13a3795e4d362ac023193b95427abf41c28c887d8dbd30cbda7a187139dfcce48357f53dc9dbfdfcae1da614fa29c3ba4e0c59215705c599ba358d165fa43ca12e5dd30a6d1d74627f35251d5ec75c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1023b4c512f64f713b55bef2b362e92421c5f6f7413a45570b32e4c2b2d464ea9538f1af7f2705de11b30d88c3859395de20c066cba068cb8f65458ea426e43f67bff2f499e7a9bb9cf2c1ada145041bfefa656905ec429914e344fe66f130bf5e0be2b9894f8a02dda;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h172a140d1a46b0fc84bb75e9d9e00911e5b8199155e14ccba9bded528d81cf60107293021aed46aecea60336eb86ed0cc58a97c2ff7fca61826ae0963be9f613778b76425b93256acf79931d55897a0ca7f071fc561281d924d34a786b920c6087a3d2721a4d4df29c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5e9687022dc1230c10babc8e7a4e0e0ff9cd6f7ce80fdebae8242820da0146ed3bab6cc28e7a5107796a77fc5083bd9479324516509475120aa8f928980aa5498041d4d7b6b4be43b5624bb14eecb009875a58fbd5c96f53438c2141d23cba34b85b85d5b212f312;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9974243ab7263cb8fb968e11d5472a2fce9a3c9b622387e170a5dcc2f3f17982114b014b409839931d22e693ef580839d03bc7b04026c6ed68ace94549ff715babd133a585361a326a85dd7ef4e57529937d45b8afc8ca9c73482a35a5d1f8011550c1f3752a7a156b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6fee353700895957208a304adacf36c9befea243ee52a9795c215b28765f57e657d25778297ebb805dd0216b6546b04aa83cc0e85a0bc27d6ebce2ac6af64ebaa1a9b3fdca1d836c6d701553d5424fd6ed6940dec522533eb123e9dba75872302b240408fa87355458;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c9f09606a3183c746314e91fdcce239d0c4f18f63ddea11fb473ec69698943635f560b909c9a9860013455b7e8499fd45c70efdab61ff504b5f7eb1a0be571d38711919b596c1e2ad4d61e57a262c41b1c8e20d125b595d8320ec26e14699d69c3ec5a9b432c3d1a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h22a89e10a35f80bb9ee04d1d619cb8b4a71689186e8863bb0728f87aaafd998e6aa5a18a83673169352326e28bfdb478d27b50ba0df424be211727a2993fdd635343365eca890f12beb5b74bb63cc3382179d66f491390aba50b188fbdbe7a3b8fc06305bc6cdda11d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15250f85619441bc0ff0a19f7616630d538705ac81f67d173f3d99695ccff2bd402a5272236eefb00519f60139c0d23d61c6435d4a1ff4fe702541af61a4c9c6f60b066697b1530d6cc20b9ba38b3492ca6a87d35a622108f38c78ec3ce35a104c50a1435003b5dec50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16958d0a314e9f19f15b5868d8d426cb9956cffbc7afabedf2cf2dbd6bb2ddc8e6333ca5f5b50c2633f8a044da98d31bdbe16d11ea2d128cc3520f3ffc13f86f0b499fb4d69c6465cca67ae17b1db57f6a5d5b75d4786e2e5c2455f3cbf4fb901a080251bfc719858d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be2b4e6fc99fec7b5711bb1af9da891f7c1917bb242a1ce7a87311c434e0cfc4163ec73d571c4cb4f3fa48ac524b421677b40d2d914d623e7bea9f4a45d156059dcbdecbab2041475327ff6d986a0f269c1affd111ed0f6b346200fdfe82ae35f6da1581d07df08d30;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d93d8b0bd4bcc3e50ae4864485c7f4c24039af0c3f487964baae06024d12b7fbedf450ff68b0b9eb203f772e5cf502a923fc6c9cc64888d6e7b9e79be9b8cf06595833900201984b5a1c9c3ccf7f4385b5be4c939740d0b9ce5f573c3e61dfce4ac9a72ac614e46949;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h769eec86bfdba7d60b67e0086e2a8917a2c601b9da32f01de111756ec982af7af80c808b4ebda3890b18c82deaec1e4138d9bf22831376d774d7b3e981429cda507819095ea45715622071fdaa4a39f5349b1478586f049e82623686e97efab6b6697bc035f85f6022;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4c282db1d333b8e783bdc205c7504fa5952dcae47e9d9e53f1b8f52d23a0538f2d36bf087c7885ca5fd4f05a625189bb659f9d01559549d20d9f57cc35d2e5c40e1cfddb423417a9a7c3c1b95219a07b440b344106beff1a8e90cdbdfb887b3857094f19b210797e62;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f7f8a6b49da2708f0fda73903fa98a08888737faf8f2665762d2f724ae8d273643d19bf49c5f5222e92f6013e1247f4c32db0e1bc1a2b18c6f90884de73ded634aa4c70b2113a18c0ab71244fcb2429eef10bc11021128bb2fa92564b114ed3fd1d643bcffadcc612;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e11b25ea35dfdf4cdb329c688a77af66fae50b03b835e735a6c29ae092423021c135984afe2a8b3fa7b8cea223d4a733ab10dfb8bdcf4115ce6ee45ac9dd3eee03ac9bb25714e4b16cf38f936afe0404b35aeab93c182e390d4219a1d5501f0239b172d1b71029817;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14ac3fef9420f9838a9f2b803da425e5d397c03f95d5eb79245ed918136a902dc6db5982b57de10aa7662647433a6edfd9a64ff877fd7149bf9988bba1dde34e4a0406bfd6be570aea359562860a8499e6f9cd33397c8290f27f09400b0718dbde827b3962d38b11c37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf425288d1e4c9b04976f829728815a31a4ef273b731500ca7dbd025284f329e32bbb320a95d39240779c6f1baefadaffefebb3a839d7b57fa2da62270820a680c23b1fec9d0e9ae336110a7fdb82010622a1177027ef9be36dc4e392c4e5607f41e607282a5e1291b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eeb5421009b5b1a12912fb149c3ae091b5e3e1a95a1e8096e5280845fdb07b0ffcdd392a18b7f69efb98d2bfc1545dcf711d63c6512bce7e9953bc23ea06d4d68ebb3ef1b55a7b80a7177adf62dca8980f7ea51da5434ee0208c57ed8ef3fb5d259abfa369cfeb2f77;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15506a4903cdc1fdff19d9ce8f01952dccf549074015bbd51bd09be6ec2475420ae571a2679212b1befa55a0d9e6a5097bf53149fa205256aad69191e1b1c217c48ebba472e57824687b535857d4bd2d8cad96559b22c0b6f0d326ac1f3e70ff47e8c838a0ccc1627d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h815803e01b731eea45cbfa9a24e092dc85ec36c1537731da3a1bd2505de20ff42470ce096e26357694610f2bbc0006622f41f4a32dcb386ca44c72e373f954502290c70bb964ce87cc0846d5a0b77ca708ea1bc14c36f3871ccd0331011a595317c2e6b602a8bee0cc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41b8394536a486dd073995e9ac77cca4568cf4c7c94c8d6bf593e005f7536540c1eb0eb622621354f51b2639df733d478b0477cfb7fa8c8213a5eb5b95d42fe2d7e8ae01177efbb1d40b842199a3ce3349a5e54e8722fa0863f57e09be4c84bce8667d5b4afd8cb44f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5238e6800ff2ef196d8f1d29e891d7647cd560c86bad000c58c8ba4ea5aeb86222b66e32090da86d87de7bbae8a44c3ac6b00782388f3ad35dad794017f9dea3a691607869d52faa9718a1668342c67ba741c8cd25c8b9fa6c331024495add4afbb317c4aeeba1f3aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heaf205ba7478804638780ad9f528815e149558dfd018921f7d52308f04b3ad2354d67720b7a7f33fb68574315229992f6f9c0e4618b4ecaf86bfbff7cc09c9b6f2299101c695f6f0b0325f06bf31d4abb624bebc2e3925263cd6a01dc62fcb17f959adc6c1ea9a8688;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf6506098f5eb645b68e594c539841eb543b89b149d13ef51e475bab485fcf323f81032b6723050811318ef70706bd5c3dc27038aecc7a439915764419641f1ec10f5ccc6ce2b39affa196d7fa50efa37475e6bbd85701d15e520a25224caca3ecb32eacf03fcd0ace0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14943576b4db50493de0c08f45e0bd2457846b8c473994aeff580816054a5ba4c767aaf34c3ae8bade088509eadb080c16b912f55fd75538cba361048e6019b9cc24b70caedd133f298e94646350e88d1862a8c29a3579107a13b260c51987df014afe11ed0b8cd7cd0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6fb3795e053b768e11a1be3ef885aa6b1bef71eaba6ce76a72d8744aa71d7aaf71f9509c5eac5839af1989fff0fcfd64731eaca5689408791d436a6e73d0cae60c26adeadac2184e87903686372a07a82f42d2b449d5017b268f30ea8c3ad82bb139f7488d3128c33b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h60350fa9200023f55bb7b6d67204314596e66c7ad7fb40727bb11b08e0928268ca16d27720c63518526a326f9e2dc5bc03d458c333a0a63f0e4cca2e9f491366ab74dd5309c6f8dd16491c59824f798d95cba20a5f589e0dcb45a8a6ac7ca5c4994eb0a4d91efd0158;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a7782a1cabea28e4deb1c45ba4b74fc28ef5fe73f3857b0ffa67183712b4f6574c6f5d3a3e78760ecf2fc35315cb09db2374b711675ff4d2a87fbb66dad8f686dc001bec9209a36dcb9d7ff7da035a47745f52411d6d59463828ee6c4c1224ba3b52c653f77c66c4c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9b809356da9497c74d469c6250757676a0eb8e7a8790878cb8fc59d54cb2e8adb7508c414f9cc43dd1424743bc802769fe7aeeb0fe88d462bc9176a6a7a1fb330106be0ecbeaa53f4b5078972212dd79c1f9b6fc28ad897c2a8de064119b8e4f351c81dc27514fa0f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14dd3853e1d82386f889ce37132c9a6a844dcf5954d2aec10a4c801a4571ec6d49bd09c0997b92215caef54a4bb0326ce615c71f688e13602dd45d045b18748cac9aacd08575f8ad064fadc73de7b0099fd079766f2bb35b85232f5bca6a959edec870690021eb6b37a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdad958db2e672adcfb34c0b7b7a0b9c84522bb12403d275b49fad5c921cfb5d801bf27a11bd0c8838c1f3c072962f8409982fa9babc8eee5395f9a9f2a496c107f274bee3e22c38bb3d524ab473cf3767e3a0c0f48523bb0f727dc283c363f6a7b1056def59b8d3a51;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f71245d9c33c4f3ef728f85dc09923143c407983160b5e0f2330310ae50ade1d1eb0a9864b22aa1c4f254b18c3b50621c8fcad4d52a9896c08ba2a844e76a271496dcc27b7819a018dae5a0284f46e850ba8c1c48da7176b314651f893a2c29a202fd256ee8558087;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h627f3f5081d52fc8b3c14cbefde425049712017cc37e3f44b37ca18794e7f17424a9706a31d71b74d196f47cc37df17f2c2943e7cbc7792338dea252e8bc9f5fdab934c3d9559c7f99aeb0564e4eb28e795defe2d372ad2990b40af309287f11a97ddd2d06c092fc1c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8414b559684a6664c38687591212f936b8ba3068308b58f4988b513299b36327910730825145807f3ec610b40be9bfbee431f4f33894b4bdd9a720d095a3aa4c14f82f68b913daa10ea6795f64e64d4510b6ea0adf38cb7d50aa3b94fcf090d8b6fde612a67211aade;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a5f37e94f4e23d88840ff2798f1ca5a6e311953dfff8cbcca2bcaca39fec3990f266f848d419083a2b45f800893a69b86ba76249010ab2b8d08dac67af1f43136c2047345fdd16513e51c9bbf1c573685d0ba9cf90f7945a45d2aa7a850dd0642c753f065be544f737;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dac9caa04468abe1b92eb8a3338245ec072fa0650aad48d4f21c4b2586855c5691ffdb54ecdb9ae6717e85fd86cb28ffdff85f8f7b4558c84bc05a0effc985de40547638d431c98f634ee375ac99cc7e6b3d0ed85d831c5fce33fc822620d9efec2e418b29ae003224;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heddc869d0441b4adee18f5a167da5ee2d93fffd63b936e04e59198d9e33fd4aaae2c6b25855ec036b0a72e5abbfd433055d5c8abd16eb0d1212a1029cf040291b6cf075bbd8052bdfe7b0ac1ec3f635f6da3b1a0aaf261ac61a8ceb5525e783ebed11d173ff5202369;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13d699d04547a81e7c5ba77cef2e216073ea48c2128ab0464743c838dafe6ab1c8bf17c0e5de804d4b643ebdb9835c3679fd0af288674a44260c30c05dddb7f3ba5cdf8a6d05f479890b8f44f651a2256cffa9d3b6f5f2ef39ddd20fce8c5692bc6815252967a31250;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h60b8a4c216a790e84e731d505ac14c27389a883f7f8b786bb833b01b907465ce14c747801d59a0251db0b44d85b06162696d72a78b531848380a05adb00a7cf00a8edaa5aa79d15795d192fb3ac50ab853f97e47a00f5f1d6a5571f884b2f6225da3610b4ad8e3cc49;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1effb7055e2daccc0ae82eed304474a37dc7e586e8da14a61e8920dcadf87cd1ee4fac1aed375cab946633a3b1c460b7baeda17625807a807a420639dc21050db83811d27a70fdc567526a8dab31e4c563861e7ea0c1f41c104e3439ad29a4a5a283a3568fbdb059be4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62dae4dec5989cdfe7ff9a5a33cae4f2ce24ff6925a24c5bafd8977d6f011de6ee295d430e770312c40a0d130c644e7696d7f1de5da345bebdb34de67a8cd1fe77727d3d0767965ff1de6493c157810f21faf11bb5348ea240a5dbdcd2654af3a29522d57563fb6a48;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e12774eb046a9c1dcececd238453b781f5dd84d6b5c0e06af80b1ab310abe72e5f9d2e3ca33093004f5af02ad66c2df427908da8d6735fbba418f912db7d965972131f35af90614d1965878a332d9dd091be694c3581dff7bc18f90db2c4a3fcfd16b218c2f72325d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ce1970c84cba78f3aae095166cf0033e1f52c060b49d4c60503765398ea17b75bfeb049e18d69e071bb8326d01085b549f048b01e54e05e6f5c22d9c7f9979e5a2d18872559b21aafdc9631b9b75fec2b26589817d3bd95ddf47441d8a5356699d8f14f1fe54124553;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17803ad7bc1fab41a2ec5d757e4c15125975de1b73235f170d15f59c815e8f6c1530557db0a799ea925f2c53864c3c96f8571b12b3c0e99c1b2f6c221b1a36c4c4b60358fcb5540706d394ef95ecc7fd9eda5da1bac0693be23d01562706da11844dd6ecd27a22cffa3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10060d9e738fffd2632672a08e5059792b2e5a18903fc57ea3d6e1afffd5cf31a0c718162f44a6bb8486653157a71c9735061b47adb26b0c1902184f0f61a53a3dda6537e377ffb52d2062225e17c902c61c101848db2b54ac2658d9d179ecc8e6843fa773cba5e20b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f4ca37774cebd53f3839b1fb4edb7e9aea796e0b6a1edf23930e22da04cb9dc60f90f694b653448a910d291bddd8a2079b985e3eba9ca43912a67303b8a67c03eccedfaba5346cd739d6530abf78ae43b6ded15b3380c62cf5a1bda7827434422b403505b5602a364;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h684b6036d4d1cbae37ff0b694c6640a828e24b6ddbbc4e500047b4587a7fe671dbdd2c9ee2a7694e1ae75398fce605b4190dfffca5b0b46645bacc83f080239ef4ef2c8e161ebba4b0b3d462d66645acc99a294d06240989ca3a27374afdf0b6313242212cb3459c45;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2000a4e3e1b377a933d2a22ee36d66900e85c1b596b9d5d82d6b5314c0874a747bbc94ca242d08db462566868311a8591524717aa4bd4f7db9a2b7ec9ea3a77b5b91278269a2c17f3ed5d28e0d4d8503f402cf08e5a268e0f334b4a63b5fd978da20a2897a143f86f4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc00ddb66484e66277202db4d72b526a35ccb0631d19c29a72cc0b711ed3272aea22c165451baa36906a433395f994f15f84b90fdf91287d6f1cf74f432e56a3790d63c5cf54431de2dad43f5fddd75704d19e02090d9def677e2db6ecac5ac0dbf224016a744370f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha4e9f687599dcbd51366d7cc5ba4ad45701123ee33c1a5709a47d799a44c1c675d2c077da1a5917e0ad666a8cc13bf78c11ce069faeec12131d155d5f2e1364d1ffbba83dc51fd3f9930ca08e2ba0f4e2116d49e0a5801e3a05d3b2960a133571b604c9367c4fc0a3f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16972aaba4a05881d05ba992988d4fb4057c1de4d47ac7daadc3232c26aa4fbbaf789a963d6e8af9deb984f2437f2c5518ad2a23d5b44030b09d447ef663e6443021262759b94e91e6af35793d0eb8dbd7a94abc7d2a62b7b7fb65f63fad106bdb21bc8862f9852531e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd7e992d636440ed2ada20debe2f8ecb9cd7dcdbd9b09ffe40b0515c882e67987413510128e59fe5f24704e8abe8ab29ddc7f5b563ad344eec6e6cc130a35a9a7e9a6761ec2c8ed0be5d6ef3c8e9defaddafd1e1380b1d133eb937c06984fd635673f15645d08bbd7a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53bd69904b88a7a5a75da5e3103903b7dc44f67579d27dc221b45997e70748cb1c7c6f7e82a707c54561ed75c1c4eea6d2d6ab5dffe229003c85b980d9d2dca636ec7d7450d5a1abcf3a2e582dd98dd736155e5c6d21607915bcfd141ad886643f18520938ac75e6ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7e510b607e48682f03af62ffb0fdf052a2895d7c6d2828970adc345fe3247df38ce0b9be8140f3a448273137a1d3f11de94badb864907bd9994439a6780c14dfaf3426007892a12e1fcf51f75b4f405d03cda8bf6d41bf9bd8eebca7e12cf0320e1c1d3e647406aa4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hecb1f8a0131459cb2b946b635e889b65455cc26ccc11445a5031f1c7dde9881f34107333a595a2aecf879dcc3c3ac2527aa8e31da622b7a27bdf736c6f5f8f9eb2b31949679e0260bd158114f43500b77182f5ce0eeaf1bddb8b98040c8fa5e861e4f522335889450b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d28397476ec48b2168530265c00ed9e1d93ce2ebeb7f93204f85cd1df1a18a05057c3713252bb679086044db90b1c393241f8a7cb136426781fcbbf3871a957b30fb015a5ff0582912367f28c6384361363574367d339b863314548901478d3535e1d123253d1145a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2021b89910e7a1e6d2d4c7778aa20a085c6a17bc645f17d0b2828c75fe5a185764131edbc298e4fad6b48e686175902cfc233ce1ba201e63e4c712aade135790730967a78e86c1ba8eccb4eab9bf16dd13cd6e142c47a42fc19b59fc196466f0433e30db70288985ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e1ada88c38b902645d86e781948075b4cdc73da861f3c53c8187ec98ccba257f1e9017e68475d1d9d8a13faba6e06982a3b72dbe695233952112b78c190984825d7be3d7d2262150948f98de9433e3ba0074552aa6baa58c9aecbc4c1f0e82d3bfaef8f595905b827;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a9349bc74272f585c73670361825e21924b383fe544ddc738a1e06a123e90f50ddfad0ee4261417bf73faba96bdf4256a8875df48a8510c62797bf4c47173ad0fead605ddc202210de8be91af43b44322c9aadbf2b2428a225617466b1a0040a1ef6b0b9b58e89cdf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101fe8ce22a8ccb6e413a6b47dda1818c6285212f9a44021b14e2fea56c9f6511d31cd810f32dae4745786f5dcd2046ae9ddc68c3207aea615a3cd3df4599b4ee0810c752c4adc8beaab75cbf553b106c8a89a440fd6d10a5eafaf85b88b937f65178b36f84206e2492;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbae3ef48ee682c00627453e139e24696783442987a327097020605ba585fad1f94295d15d46e723c54cf9a51eb2b1e169fe79d518e60a0cfb9377590c522f15b3c549b18d2b7e02ef7f29905d7ce384ed6944fd6f26c844663720ae55d92732ff84634fedecc76948e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1588d10bbb02e1ea75f0af29e3a46100c4b66065d47fba78fc27f44c4e69d75b3152e7066bb6433ca33e8a18743923a9850c7f3f521139bf06c9dfb3573718ee8142cf8a324a49b827fdc9ac872f2128848c3e2a9114967ee8faa5fd36b7726a953b52d6c177ad7597e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d0a0559ef876599bc8a7c11a80e6e5002129d2391741f0d8d2a2b098e87c40e7537eb47ef8dc06c38515dbbef9b03abe49a1c9782077975c5871155a6477e177be2ccef01e62edcea0042106851dfeb240a3034ed42a0711fe5b96d4e8a3fe7d1abd11b3c3ea4c333b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1335542ea8b67fc6fe47bb498aac0850924e3bfc2c52d321250e7d5d0ac70c78818cfec99b49a7bfe43b8e00f172cbcc05cfd0935ed793883efa3b016ec252283bf459851f5b978b4d77280782680be7e8e306d51ce08a52da2d9444ea398320a6d77a33d77bf78b190;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc6478a5965c4a3cea57ab6463ac45c3f050cf73a57621d631be6aa4dea00d0211f5e340c8ef2bfd0da21889a0619086751ff990bc90b5197c00eb452819b45f36a9b77d4d6ae03af53790a6c8bf25321623f2d6da436db846c8204e557509070c373c10b7849a20cc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ea9a5aa3eed29fb31b7367f29368f486f0306179071535496b589eb161b6d41fab8978a360d71679a576f63bb43797ef21ba039ab35e26ed94ba394962931aa00a653ff76bc13ced4235eede592ec6a98ac190e2939b3410156d4cacdd8846dec0fd0d7a7ef59f9c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c56a7cac9f9dfab582d6206925270599d94efc86ea09ec3e7db037da645838f2b3c7d572d8dd8cd697fb576f4cb3953335262f8da48cf008a11383060813f8e2f753ed2842a9fe7165eaa9a1f35dec24b58a27fdead03d7b914aa796388e01754145275e77603a4b7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a5e9ba5b028bf09e6d2555f9db54616e5f64346796b960fe256858be8ffc36c6e0ca6636d012b09d880445710c843c3f0a3a530df41925fd412b0a2eef6332d50e763057db23b91a5ec2be29f4a3f24cae6605f7728d3e9e1b30d935efd9224bfec3c9eb5ea706524;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96ff8398d0fd35897110d613d4ea415b0ff13bcf943080dbdd9845670f59d570b5bcbbde26d8b83804718f19ea2ee56b09200523f6417f54f657729966723647254c7555a5b5bbdd2647167f92ab222ce537cd5e1ddcefed329eeb1072e877118006f37cae1863b7e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb10b6c6ee8ed094b35e8bc9ef28c5b586e61a2e4c186d24ea94cd73de4f1d7baa3d437be21888fc8699f77e4c4c298c056b218fdc7a88037b33eab3640bb27fd1d556c4a9fb8ff9649a871ceaabc1ae0bcddbe6d77905d353e75e09fdf3a8150aaefa5a2c62c5cc492;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3024d9ce2caa5cfca291cd4006dffb2783586d181620a6acc57fa15e0e90bcb3564c036c7a5ff55d6a889fa1f0abe2cee9083ae3dab33adc2e7adb8bc3023f96d9512560d5d4cdc4a3b054bcb7b6e914423218a2df60152372b6b92668781c133ece02e966ef972508;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b48a4adae89ccc7bb69352f10834b021ea2e0da8f273c222b42118449b7150a73716cd3b2aef3665b068d99285c090930b0707a8ed6e3bda674e2ee2d08373988cafd038d411453f2e687a0ddf530f4851642479ab2ee5aeeb57271ce2b5956d005645e0c6cf14b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a7952cc07d27a91ff23e1dcfc3b5ead9d72709191ea83495779580a469f5976ebd4b0b3a63b8621f2b6b9d5fea0f48fc9cfbf2b624ce1256371bdb34ad617037184bcd2b1783bc447caf3e735c64739e1e57a9beab046144dc71bec3c5d289be9a74b7a88a834a0295;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d46abb8abc96178169be85bad9c3f5374661eaa44c3cd20ec6de035c6192c29ebf1c3745255e324f39abd45026b5c478dfd021bda5b4b95cd57c255093a994e63e96bebe878ff41260fc8d9ce6388cbee1f83afc7efd5fce5860558f41b49f6cc7cdac66baf93527d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h326efa3ce31379c84ab96c5c3a4f7702806415ea7a9ae06bd7de7a83b241039857cae5051ecff4b6ee49b302432e7cc429557ae3b122ff2fb3b18d9046d94853736e08ca582692a9686dd13b870aa8034ebccfa3c0bfe23cc713ae88538b52ae649ddf9713bea75237;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea57f00b9ee45bfd744e3572db9e08fa2d133d228eb9306b94cf57ea03bfce70f4471d772551e3849273f5d56dbe44a461d846fd4fc87d326eeda30681245eab151cc012b447e8421b04186663f13211420dfbcf1f0316869a13db81155a5ef6531c22b2e1cd2cfba5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcfdaf7db723027da96acc0690b8feb625e81647e4c8a56cdba503f4e09d244ead724ebfe7defddd65790b3dd243362b005820c41f94bc3f3d49382d98eab7ebbbb4d913a6647d8007982ead29c5eb79b264e09e71572faf6459eaf567fdbc5f5033911f3dee79ef739;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h152ab88d4940bafb5f80b0cd77fe10f7d5a165c6c28c5501f03269ff627ffdc624da75c2a17192a43d3071ea0769c590e365894f5ac8678e2ba44418ae56cb51ae17369273f9af11a3a37a384d75f6ad40239de10cf23d22171b7c25d096169fad945d024a2dd5a26c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h130ddaa71d24ae2387f4ee9b401b494572e4a0d969578e41b24b8d3ef2f83fc3be4ccac90c1b865d15bb77cce3b45fc4de9b1943e1ca9cf0679473af93791e66f3441acdac82e487d14b78fd5f41f70252ab84f3c7bd8a5eb04397229d28c8e0b6384927b42bdfc6a50;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10de6f6c211dc332a6673972bea67f18321fdc8ba3c5a0b0e542a8a4e09b607d0d70dc8db52793568796a679ac072d597d0caf26661c26f4f8b758807fcc97fdd88fce55d983a42b5d910e39a904263bcd40b2b6b4c8580e8dcbd8a1da04247d903c2658bed2ba16be7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h131a459f62dd76f77ca41c46fc39f957a27f83955dca93203b2cc7b54589d27212b55ea8f4c20fdc1945a7790e520ddd78683d2ba13e841636d53d6bb10fa66f87616a357ea17883bc2f839abf731213d8c2fd71cc0138bce2dc289ef543997bb5538c76da57cb06d14;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9d220e7ffa8d287e0b9f783fbda1912b96f6decd223f6fde9bfb4569d16238deff790a2b21f39eb7a374cf16d4e5d7aca9f15ca5948d4067499719f0c65298942542e063b767c97280f7db9fc10057a8c2a76ad03c7ca9ec281f57a3d092ae18af07e2a6d1bbf7dd78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca4f332791180eb33867d2ce289bd250c562cab32843786a9de8104f1f1e73663b8771c8cab5a5b8c7d42eaff3e01ccce2fbd19cbb8c98b772f5464df3cf3a95bdc168a785eb79674abdbfc85df9d54b9d82211ec4e7b06e960e7e921e88bc0575bea141b1c2653940;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ae935e3417483639330bef70913fdf8ee1927ca131d04fee693b78f4c0b41089a6ebd0af09fd6c7b266b4d7394ac611f6972d0a8a8894a728f6adb8cbb5ba5fd893a2f49da749a77359f2bd4abc1408182a11402a09915b271ec6ce96c9732628f39497e152726d92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf04e1306df4fe9d90bcc19cc638ab78ade87772c94185fd3a83e51b9021026ef5694150e05b3e0eeb5460ff4f1c90938fdb3a4ee018bb55bec7f9c25df2bd764773fe89d9c2b4727eae1204411cde3e65a259776e3b11320c6e73c3a378cddf88e62561ff18dd039ff;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80a1e84c84ceaf0c373f6e23e5dafa35cac3f745f32e18702ce5791b75113ed221790fa01b40b5c7ecb1597a7194a2ff348897b3cc4651f01f02b5c39300ff64c10fa721122b211e918d22f91aa18ca643a724454ef8c70b9a4be9e6af4e5b35176daa5915a3837bfe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3f03056cb5b9de71c8e5fbee2c2fdedd20f2a4a2f71c4f47e5042e5158639cbf0dcbaba50dcd973577c5aabe8d6260047407ede30e9dce54c461c9c07c62c14a961dd0f1089d557b25f42f2604fd062c7c3d3019b8329d94c11189fe1a7d0c24039eb7c1e867595c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf211abac3e0e549867d6c7aa16096f067acc0d1091cac80de80f479f0fbe1d014537363324bc192205b343de7ea270cc466b373731408defd1329a3286e21f07d9faed13a0fe433a4ec0d01910866705508651417c6a7d86892c0ba49d0adaf332e9e7567a4a1f0273;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hecb1b2a7cb9ccaaf7c19f7a79cac2e0451e53f354caadabefb8101380df2a65423dfdae934b17f93afb392322d69d9a6e463b77b746c6750cde5bdea2cd266f5ecfc2227ca351d156466d685294884e27244108e078337d6af6606cf72831fda6647d23c9c37677bd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b358a213e0d68778acbe4664d4122f225ba62d866dbeaa5b931a09c4c416f602b5956046770d035ca44e88f1210d6ca60dc5c51843057f6b362a1f0ab43245ffd9cfbea0071af013e225a25356ce6b9eb48093690292325230a91d240c93d119deafb8713bbea9cfc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b38932c515bae2f312d9859045cd74497f39e1b49ad1cab4013543097772639fa473d3715ff4fdd0c0c77bf9dc8882445c6eff60b10917548e9ce257d51c8be9431ac6cb10989e0c5798a0fc0322b85e58713d9834be6b70f8a3e465b967a8564571c48835fbcf9c01;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f14dfabb96a372ab4e0e600407cfd46d15d92ac77b2dabda956d2ec563a9088a1a8d0060f0c57bd7f863c5dac632621d3954669a03208e12e900c8c2f5c8ce13a0d0f6a61e5c492ba9723b1d4d95badbcd726720b92644c2f146b19faa8cd8505816348a8cc7e3656;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9b188c986f68be01af5ec65f43669f25c725dd6030d6a7f40df9cfc02830a91cee4b34ae125c1e3dac838f1b06449600751d2c5adfc435d68547b8095a9a13279e3dfa2be7bc642257cb155c8aba02717bca7f01367ba73b41c521b70281b20ca035412d92ff7dceb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h96495045ac98411d647564a3c0c15413c6a7de3e2820d12bfc6a2e9742df8ac87a095f9c3466a51990937de6af84db0907910ba07f6cd3be138ec8a6cad32faace6a03fee1ff207ae79b76bcf98cee48cf0c49049075e64e760051064483d71fb69492103303cabd19;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h188c188b719e152ac6494c7557b7b3cdd9899b8f65a6cbf3c77d66624462e9cbb480f5cbc0dc1f928898513f6c9f5e8c5512c870f0f47ae28c2f974b5a522acc957285b9a172d2a373bfe838b395cf398386138dc4d4aff0f27bcd6f34d798092b33e4f856aac4b78cb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h89cfec79b883d8e82e7716307dd0f57bc36bdb5b8c18e832f40fbb543da3831656f7aa57dd831f5694f71a4b4f2d8d3be9c6100c0157761f86e973daae988c806e34c7a8b31ade36a9b50b427652a78f8b3c3964749d2acd30e7ffccc583e271b5913e4df7e25a2439;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e5979449d2be24e0edee72733aef36ec0d9be4c84f9ba55d326322d293dacfe5320280038ad2c1e43d32a8d4985269fb6c361f6a2b16427498c89dc832be0d64e122e672230b9ea785043adaca38a402b22c7663cb0d37fc515d91e6c4133cf3136ed9eeab79ebc6f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb872b653a89df4ff51b951f24c3d66de606748d13a350161d85a42e4f2b337ab5ef55808241da65e0e368e37c6bedb443a65bee5effbe860461446a04577284041c1a6e5e0b7ab93b785994f037785524e8d70aab279fff2b9a41640b972d55e159fbd6760b79fb1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he3dac9a987c22e5bcc4e2468f8d31107f4e0a29927f6424437c044d1aee497fab63de038a6be206ba0406917ae7d48be069e4d5f542348e5c55532ba473543bd4b0305a29d263ec0e4d796bcbc8d38650dd7ea360b9cbff928a67adb72d68a923453ef53bb58f78458;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123c3f7e3d762fc095ebdb699e8d092b8b3d35e285ee306a088acd0f1c54619fd348b80e349b396e8346ad1aec7c9c33eb881923182672892d0282a4f2b8f48816fac24cd508036f5fe4f1aba6b01d713437c4a0c5b7a6285956a9ba4c3cbae88e3c0fc7d2102835bf3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147d208ac8d984bf351f93cf2316d0af785e9aed79b529a4a8628c0421085259540d885786258fba1bb11018fef82c72212a688af8cdb5f07cd29638112ace45a9dae7baf1954ee61b46324cb5b76ea289a1bdf852cd23be8d5bd54086a2921e7bdb6254f870fa7e0e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17bd0a1270d21c782b2aa0821a26321784fc2e1bb449cd06836f93e6bd0073d80e8d344a328568b0c1c8771547cf3c23baf0a1a5427a0a98efffb91f3aa4415c089add0ad6bd4b7550bf954576897e9bf2aa3cf77c57b724749a355822b059190e4ffb513e149223b51;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16ef2c7e823db2eef7fbae109cfe2d8df561270cb4597af5bba9cd947abed5dcf780a9fb31231395d529ab1b2be6733017716181b8ae5bb75e598afdd885765f9bf2a7e7e7459d29c6e2ba5b38d06fd9c5d76161c3a79fa578ed2843df1820f857d1e187cfed0816dfd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h66d26950dc7f5711b64cf4ef2a45f0184befe889698ccad77a4c18e1d71842fd38a07fe81c68df3903d4461ba5f1b34d596f67f6cb86704bdd18f9246ddebb02a97b3893f5935b50debb51fbd1a2d94b54648001924873ba75b32e61ac399a6f1e3046b713424502c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19131ba2320abadbd5df90d2c0ebacb6eb060efbccfe87e2ae8d6f6a485ec75cfcc8dcc79227352f46f6a0d08df84a6623ead9acf6e18738dbadacd17e5ffcbdb3d9899505ddbc2f88c911b849bc34117ccc1236138915509dde7c2ecd12e0fc7fe3a70d19c88ed4e99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a101c312e34fdb19bc52295b2608ba341b307e73292a3b33726b35082f08462729e62948f814226fa76b0a94605f1718cc0b9c9b4ddcbcc920b0fff93a14547299085043f0c9a19900a836834e0adf4e3c4276415a46e7a1a6e9920b7e7a988b60cae553c70b26c07;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1607a8d9dd5d438a624fe567002b27d3a7bd2d728613d0562a3eef7177453062b4a85393f432b2710ff874e2571a1c765f057034d43e09c1a5c17a8f47181937d542c6e39076a6ea8de9b4f1719abf9b1f2aefdb377edc37b1add5554325e421ac9c989595280ddb8b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbb13a965477e80c4e85e03c192defd0186d784930036c3987e84ae0ac5b40f78a6cea865ee8601fd3ea2c94c925eff39b953f07d6fcea4f9c1a63063917b22425293560e3e841f38a421a9546527c556caffcda02a3b0da8c6c34c0fffc4c4c306100695b205660f40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h452767e3c179ed25db6181495c9fdc340a3f698e39e6d3d2b1a402cfa26a9d6af72ad459fd625647c6826cd1e74924198d1de24da6aef5b1648b1f3e89c15c7e3182458d9729478613d89dc50dbf3797a4ce54506df3f100ae57ab403cc1f5c5f7138c48c78b716038;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ae7633a75a2fc007141204158201a03e7c2604630f7acd04e0e25f7d6fbe5756520876d05133cff53009cd10f332272281259d417dd7f2c3ecbb94df31639ed874c4a4bad21469a2019b5669a5331ce726bd575a773b86ea859dfcd4d7399f151d6b631ebf47ab28b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4783c42add2f3bfd623965dccd020ad6354c6c834a9ab3b469e880384d225f38a35298e36a740e259386d2f87ea46bf6af43d46d50f84edf2b0309c2a80d4777fb6e3f1b121c83c0ce6fd835cfdc37cbfb417bd7fe0606489031c7c5959bbbd5a85aae043242751212;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf6a99116e592daa38d603f4a034011a4ef07eb5b990bdccc5f5b5ae5ef9691da47d508402423d72fd08e8595d30774b2beac584ebab5b59059d714309fe40f28844381b5084bd5d791dd8f7c793ae77da2c31f1847ce4e6370d60d10036f5f57db8b6d9adde17c4e81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b01920b4c8e260c82c8561528f2c56be18f827d1682f3d2377072fdacecd105a5294e117f33679223b4058f31c5a27a99c655cf2a5a6b0b69a07281f1402eba1853d445b418c31bd0e1cd66900449f9e85330f25bdbcc403fb85e2310c5c594a62c4156633e5c7b87;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f8f6c21defc6fe1b4a6ac69ef82b47dc7379c89c0478e3dfd2b6f81297b9189a401a2786ed876cf3f3f56874c6d98af2118b08ea80dc399ba26b0198a0b45d7f312534c648c6ac69f4701d343638f8cbf2aca0d1a9a17baef353ee37b2e21d3eddf7bd0473f14e859;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15a0ded28c1d1b9e0410645d112782e7c503e6d71139bf9ff0cf2e43b28423dbaca0577a096c5236fa74df3608f9654c63f54733b7eb5f1c9f5e4e12929ffd09d3ea376410eed0d6516c01e009b335b39106641620484c35a398bed0f21abde3175fa447035f329cc7d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf42c8faea98739d4812945240e392b2ccf6de0d12c6f1b9950a001a07a0e4cb0fe0d7d352cccd08077ae54861636e673729dd7e2fa818892a2030c832fc38ece2266ff75c50569e559efd124e779d5272f7e30c00ec69985385edf507bac79f81a8d00dd1b110116fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ca14e093a24ea1fd0e33add69a50a7c0a49b1c77343d77c3f5acc9ed06b58e0bbaa36f81064aa7c84be56beb0dade0e7576275d96692d993fc22031da980f3dcb37f7d7f9f9f72b1063ceacf7b932775ba97e4a72415e0b34295eb38032b535440ad648ba9f08d8fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d26d6f552bd2352c7109cdb85208bfc33ce9b66fabed8199732fc36c864e20cfc064cb1c1b7697f60c99ef4537c14bb92b36d2e6620cf5d7755df77e9eb67195df6bc645928ccf3d555fb37643b7993462ba7363e1b20099329837eb372706feda254afc816bf020;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haac7a9e371b7a737850f01bb0cea4ae08f1379370e32d742f434d3a628fdefcd69d8604a4ba6a44355b75ffa1e1a3da60ca892450ec2690d6e8ff3980a69da262425ba5520fa09675659850020d67a2bfdbca9b134e8530e775f05a12c1c097663f8bd51d3fc9b3f92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108f53ba61b408b545ac8e3cd806759dbb161d0682dc0adf079408c58cd88abb319e641f03de69992c668106b3cc0a3aec81aaa9f40e5f5f995a848afaf5ae5a3cb5bd38c5b8b9812bdd14ba92d1490edd6c5c245da454352e7d5aec8a159a4245e12c1cb684e166853;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa994a3413994e2b6d7f7519b4e7b068ccfb08a6c452e61312b432aa7f6d7dbbe386c1ce2beebc4c3059035c716e0548d9a7dc74ba27825843ebb3829f73ec3cd2d6a07fb99787cebd0a255343b5bc44df5d5ebd8cf9411402e19e43ae6be082e000315a4dd0d5767a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bce5267de251fc1a1113d946faf72c055f5ef3c15c7b5fe6e562dfb744557bd9fcb444b5275457a0c26f52f9747e48897ad66c87edfe8a9b1e9d2e4d71ddc3e25a210a1937be4523522ed9efe5dc02905f7da366e2ea72e1838b6d97242d339850afce3abeb841cd6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cad685fdd9ac565fef6a94b6e06e3c60a3fdd067af9465880600febe935944ae3c4213c0e1e0d5e5dbc0fe2a67373ebd00afda47c2902dab8dc85425258df6cd227a651ab6b956da2ffa7532ad104f808f0d55cfb586fba09bf02ae74a9350606405f7b4e84e2d6bfa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h102c5b55e8c2491c52e798c40425c28fd8ccb00ae9b8b78a254bfd5f3c8fe472f345bd8327fb5950869954e7b17e8953a93e501c01076d17951da64354ccb6c84629b8772db38e8570387fdaf40eb9ad9d960bb5c833c8b9093399c25d711325c6e7aba87e9523f5112;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76c683effd46735457ce471c9e6fcd8cc9ad6f0bd1def4f0fbd92d2b09357f3daa855ce22ccd5901b91426c3f5dbde52232eb3777b145c1b227a7946ca9bf7653078f1f243c32f1aa7d6c492c0abcf8bd4688a117d50dded3770d6c4a26cebf1270610a16e6a03c0e2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c3a2bff24b2911e91319c25f9165561be3360f4149b833bff3c3742315d3c701698e973c1384fe84d1c5a5a70e83d3944e5070051fb99a85fcee2800ea816021930cffd97ce0ea8305e9da1a10fb592427663785610ef499dd51ef82e32006383c7c2e6da49b43d4d3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h194cdb8b171cc763b485d8923864fde5621b936162f5ec900597689486d61789cc89c78d961ec84ce70b345eb2c37008ad520fb71cdd7b33f9043f6f93a123ab07466151875dd4d7b1ec933d89909f01c0509b577bc7f99bb12527856965d2bd12d4eebbb053f402c4e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h105084e27d98e71fb34f60407241f04a385466d9984d11c2272af8574948e6f4ecb450c9f19ba4a0707cddcb213e4d04452defc83cc4a1dd90076e0e3ba428e37be226d86fb5ff304d88d5116a1665ef0edb1b71f65854374a8d7638b20b15fff75663193fc9d7d297f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e921764d364a594976540e62b6709f3356e8fa3173365f9ff21ff147f7744fc6a43acfca959033b5bb82743964e410615ace77080cf195c29fc3b3f0ef30711fb1718841123862d6ed556a046ff49e2f462cf461ce4775a9a569fc1d6e9a1cf876370da0b9cd5f7fa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6126bc1add288fe6f6e99b547967be7039390640780de6cff014c588a486dcafa790a7930fa40b0df810708b52de9d5319abe32d5a59da0cf59ea257777ed40e4aab6efa94d3d2e6478cf68190dda06dda8b79b3dc437ceef35cb7d46d1e472af4cfbf18a6476f7773;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h59016c61737cf3c92f0d6c85475beb07418ba28be89c883133edd7cea7e6b846ab68f7f8bc33918565c836a05438a52a643e3922803a1d271a4c42d6c58a590a44e54fa103adaa0ca0e3a5badf03c90d507b7272abc63347e9d48b8622ed38a1f07eeeaeeadeb81edd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be7af53c969026fb586c360de2a388ac9493f128f4f5589c09d6e14a9da00fd257d6b41b83b2b24ade30fbc6673445162597f9d24c2b3672f4aa4d88ac339a80ffbcda09562fabcead1a49eb3c8fcaf0572592bfb56a750e29e80660a4b0a085f82b891b52b983eef6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f81eaea48c471608c713a9f7bfb1c528e346e5b2d9d728e3c286f9e2eff21bffe2cfd8e49be99b46a3f704b95130dc4f20d390b5d06825bda7af3010b8b4405006a69e0fd77fccb79fd2a495affe8b31300ceeef8311bde920dc5e92e6b573336b60bd04ca68d099b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9f493ce33e91ce577dfe87386232a986de4ea384ee2775d2af0040f09a8b17b6a5fd52a5cbf5b4f1eceeac1dda4fbe4f4335488ac358b3d705f786cfb345ec3ef2450c27beca820e7e0a36a06c731e89d1194c752f91967ef288110087d33b5d287d9ac6f8f20f71fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h85304f955f8ef7aca63a0353184ee37a6a1d0425ef8be972d99bdcc7cd269e27de30a9c4d93ad505ff2870e1dac373394a3c8ed115d85189db5fc53d080c4aef996f80b67843111551277517b82a2c099493b9e4ac2f3b3dde2135e8936be034f4514cc29e93cfee31;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h408864e3d54e0dc10a981c5ebc90d0f97f692616edb48636b1accb0c5f4ffa636307f48c7f81a46d2affb64283145a678e2a23a6e11c1d0188d6000b8d989f409951d907dcf8d416f50553c61f9728ea798be11f34a715224501ba677d26763cc599092dd65588a6a0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13babfe7f8ca3ce8e0808124dd5dc586a1a8e7d16cf80f2773692320e289118ac1065e924845fff539a767993052d635f76fdb70bf925736ec8725b5b2cbf65a92ff0bf82f93e439cb1c0d04598aee1fec2075635310f5c52ae385fdb2a5637d9b0082015cc8b77769d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h136b47da1b3dba6cee766120872c0d3f1a0d525a198b606cd1369cb4c24a4542dd09d6ce89edcd9373fb650c150ebcc1b4b087e8c113d9e6a69c123a4f09dbcf30ba446d7c024a4474042bef1363cd8de70f992dd205159551ea60f6631e34e1b46343663b8e6620120;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h88db280d2299e620e4e3cc365a7c50ac73bf6cc4f8071ca1385b633efb29419ce8affe2c21036a1c7776cd9d7b1aab7c12148ff73fbce517788aafbddaecdf987b6e53e20043a9af9fc82b461edc7bad8edd243b26ef199112cc22e3004ccc032bc6e7b9ab6ccbe078;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1071ec5cf7cb225b19d54879e68c8c1ebdaa58f17128c216c38526e97ead3ff7b104b7cdd3bc0829751553945a7d8ffa7ab1bea5777a2095dc89ad3334606015aed9326c74bc51f6a7408dcdc700ba45e611d1ba63522b5a78700e9fcc115a31e1802955a7a650639f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h496f7b5ca5581894fcfecab52e6effa4668a98de51bd7b8209693ec864f0d91689649c8304618c53859c947710f4b6a14d1912e115884ac06fcde46f3b486d587a2f18bcc356203d80189ffd28ffbe7377157824c19e68d48e0ea64371083a0099d2f59add18026f2f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dce00ec6108918cbec99b84446a36dd07c14297519455d0d24005332f36b5482e8c742da519607294c57740d8e162f3be944f02d931374e058fe9dc31d5800261f53a6fae0ffa408256b922def98f57707f680454e354e3c57e56ea1d61646a359f1bf10aafa836474;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h63b0baf2a25ffa08ccfda671b1a33743af0694a658abbeda7d262ba888d0588ba0a3756c108169253a4345e0514c8294e11abfba22c99c7a581eb6d77a67a773a0b2e0c0c1fe9aea89c4a911280988d2616dbb167a38bf59737e6e2215dde2216e71f0f6254ddb3dc6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121b2afc554e209dbca6a01e308f8685b6aeff016d9a4048e5754d58e099a7e03428a4b10277ff865bee4d991ac5694c16a2eeff940fc22c2ba84ca02506cce24d6e5062c768b93411277678c54ee6b8a3ca65404c062de96ea572a7237ddbd787411b97b12302b028d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9432a9dae5991422913eeee1120e1410f444e8aec025005d5bea5ce7e81545c769f03bd41996acd15c45636b646eb5e8e078bb2fedda94c094241ab966deefbf3122dc0065d3d4659d4c60888b95dd4281d20a8636995e7d50697eec46a15f4c5b64d833ec91539524;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16efe14966ff6b453a8f42eb9e54dd17e7da52e62b4003e00fc5e8763c59827c6d87959e2e35d22227ffee599834474a87afc91ddaa1372585a67ea58add244820b4c5e64e2b669ebdd576d468fad20c72dc72ad0f7f4e2dd2011111bcce6d36ac6c2c365bdb91cd6d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192064f79b6377b4a926b63173e4707de8b2c2354e8bbc2f921fd7e1b7d0355d2f367e2c0d7ce3b5feca78912d908c7c2acd2b9b1557697391758b2e30d81ecfc32248b044757fb62dff887fb959cf03fbf00b70d81923da9303251ef2e104a3e2f314d6d493fb720ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h177fb936257e00c11a1f1524f808d1f0bd871b840024e898c106f5e2e98effd3eca59b7487654abe15b634116bc0d7e9e5007c86cc6bef63126b6803464e3c840721de842504f49e95627b2ddeaa9a4dcd8c26e0d613820c1f613e7394cb546134121df1ef58b55bc94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1316bcc75f4398455adf567489c6abb7f9f8a570da225215937ac78bbd0c882e6e9a4b0dc2d4dba63a099d10b7aaaae682a7efa1a0d74e972671f5890c644849fb02ea63155a1789437dec2d10482b150c5a1c81dd891825d16a1ccd56207d9d036e698b59b55a0e78e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1559ab87a9095cca2685b1fbc46746c1f81d9f53fdd918067e0f70c584cd46071d05f8253be613602dc009e5a7c8c5fc75fda7f7ff865f556d4b4883dfb4ba58e7e78bbc164f0a38392d2ca9f9e23dd2345acedfb0a610b22fa3256fcd3115f7f0f8c68f93a92614b2e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a657116217eb28944f2ccd1692cd81bec43ca2b4e152524d08aea961816b736c9568be51c630775db9d66400f7c37d69bd4cef2bb7088b39d5f5e1fbab34e33009a9fa4e37a9efb30cb00a2aad8e87c4a82ab373e612722895d569663e58d209c843ba82fc8f4de4c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11898ddd3c47d763875d80b890a2bedeceafc71d029b2d31889a4f4498196f96ad07ca7c4cbb310049f05b084546ae724ebacac5ebe96568b1a1be422c90706d3f4f32bd364d98f683391b4d6f5facd10725052414451e540eadae7a103ff7cf5e7643c1e880273a551;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e48aef747c5f1117cff7f5fa79f6cbb192c03a7b05eb945f56e6ea738b38c908b4e7c73bd503516ec9393e9d82bb39e86f1ec3f243037ee61847e6310796c6c57cbb520eadd393750a6056783289b8adf014e09397a067d351e38d2d9e06f97a29256d1dd06e9ddb63;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c2fa5ef2206858bf619e04256150e9c1e047285e94b146302174f533cef584ab0a3d1a8495c932540b7409ad8900372e1119054e0963f0dbb59ef4e84477441b41893405d189eafb90e8266f880bb588246764ec9a75fb2e8c01a6df40eb32dd7262f2f66510f6700;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6f35a4d32c5a45a8d3429dd5616e378ab6d9c9387dbda38773926fd9a16024d39d421c456a40d35e3928b643aff41bd24e0fe34e40725cd6183e614f6cc147012e30e13be49efab14432ee9e0d29f9eed4fbb48b332bc2cae8baf6fc7f85f418b4478c8983bf9dd9c8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8206e6f33a0b3ec29f37f3e1680a534fd89949e84151063285b2d0046f5db0f0e056141fcee75dc332cb93460f99b65da7ab55239e14dcebfa1f977fc840694ae60846dfc907fec7639b06c7a7f3ebc102747efb532aa6f5ab5ec8332786ff79204141c861f9412da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h954de2d63a8e366927d556c33fd475c15ec0a63461a3284d601d572ad5c072a42b4a0582a6d9d01cb5612e86ba9265fdf2a8cdeb916b96bd94f81e4c3721e5b087cc91119e329e8092ffd4bd97d8026a5963b18290f06686d30f34625c793f16aaeccc38768d61cf70;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h184f4bb7b36ed7aa635c1e8612278ac863da13a6571720848449dd7dd3acc3ee4941b76d8dd1c547d3dbcc73632e9e3aa5f9de11de346b4aa4b6dd16acbd4a0f08e1aaec9492c1a1237524d3d680722db65cbb666ed5f57a6e7456a6c5817ca2438bb51316cc85670e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192df5a6d1650b15c57c5b6c5b413add8cc8a43edd8074e06984218cc2dcbee700dc6bc1925f65e3fd74b32473a5e649abbfc3ecaf70ac1698a2f083634add693013d70285667ead7b50dabddc03982750e920e7c91d44940f53adab73cf4b335ad9c289bc9bdd4d68c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e242c33e495c03c83a4e9b9482a8328727d8fbc93a6105698c77e01d8b4afddd2cffa4cdc4f2d8d1fe5c6525111908771e5e7f78c04838d5adda22233309b729ce17852b6aa6351618f95702822ee2c1b1ab76d3bfb7a65c138c075d89c2f88840cbd7ab72a048eae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2cb3e5396f5d475f2e1b7a089aa88302581104f8f2bf11a83349e8340956baf08c18a3b913bbbea612f26e25b20cf09cdca25ed8481a58d384c46d7e30b629a0b0b668ed7f3d2cee9ccd0ec4add0b740ba41148b690a94dac1128be7a9e5fe6709b2d6ca09290c568;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183b19f3b31df4a3f8039151ad6b7e3d1238778ff16a06fb21ced6278fcb9de5f50d49508cc6a9406cfda592efc2f79ae1a581c826c1645d11b4eafb9c8298ebb100b92f23b53308a022716076cfd84ee430e2f8ab0ce9fcfb0c04ef5a3b9c6c8cfddaabd95e6b1c388;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27805d1df60ffdf9f812c3832cf6ac8cc7fd2e55868a8046e4a0171a754de7602b3f57caf2317bdd504f167025447420e7b3a95566fcc9aecd1ca85034ebe98437bf29a53122901352b8f467ae3ecd5f01248d11d57cfd8433c965c92577fa18fc94398ebaed5bbcb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12b7e2fa7e8002e2c5847d2043ffe89a66aab525e59625aba8821815ad398d7ee42628bdc9ddd465531cd219cb614c7eb78869611a78e49af12ca8fa4c4e02750c1c1b61a5251634830c06f940ad38b160c54d74cc1f01b56f2d91f2ca7edcaad5199991439969ea055;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h482205b57f94a9e04ec3e09390eae86f57aff62ca08aa13264bc849b51523e9bec1245f7364c505982dc74f75298244a461b387380026eef42aee08fe91cb6aaa0ecb63fb77a7603db7a2a9806d2245cdcce1c334efca2a083b36b9b2f9fe8f0b6064ad937ed2dbd0b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a2fc69b52da8894d8aba735400edf89f8a90ca05a80b029713b97ef1120654b69772a04a5266e41457f0615feadc9063791895c00e25dd1d26750002714933b366f5ea1b0390cf11d0f7bb69c4c6b8a22019ca19684d2185f8c6786489be67d07276b2fd636e17065b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hddd278e244d73dd62ff268345c3cf81f4080cfca31a1bc64d3abcdd878b81ad63ccef2c397b8cdceca8c464953adbc5e09d6fc1c676c640a5b507625f3d61039695dca7cd09e619b4849c5d12c69ea8d42dbdd2c10dcd08ecaf7a843cf6f34ef217b4510937a5908ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h195f668f1006d5a0aa150959b9513fea4d461d56092389248065ab8ff62e9760f23c3803c8c69523c049dd3979452a49b02ea92f52122841d7c2202de9fc85dcf04c644764a5fb3576c7b0ead5bc87bb2c8f07d61eed42842520f7622f9cef1066628a659acf442048b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12cfe15f999f0ef107a95ea71f915c91ecb70448f8ff3977408370a39c04eb4a3256fc1e2483e0a46db2022ff92ca418624967a859677922d6b5d56257d3b48b915cefaed710ad0bbb148767d7ce646d54fe2b11e58a5d52096663fc10abf0ffb9c554521df7b5f135d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79583b5bddaa4ca91fc4d680741623d9bf7a02e19becd1fec6cd3277300864f57c1ef3e93e2dcf4dcb9d5ef453cb4dae5bd4778a7dceda1663a39307bdc3ed8026c378d2cb987064ecfb869974002c42fee54341f12f8115b007b9b31381de0548e07ef02448a906de;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a988ad63e3a9b364f7cf71a9b9efba32b8170a1101a3f584e32fa8eb23d239f341bb68b7c62a0f8910c5e68b2317ff3de2dd64d5de3ca194dd697a5ce49e03fc30ebdae64499f480103b47f83eae895ba5c6a549dd1f27f57da9abcd037021910c7c0ebe7af55099;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bce3db1eb8ae3c78c8c0d66eb769f802cb3fc2eb4d828f487590ba0bae383e88839a5d9f499475993f92b6ca785c7f1248fdfb2af2da20bb1711df229d4c9f7df888a3b55d89cc9465921c0b676af9b0fa48b60ade523430a388c4ae06c2c7ae816c2fe5d670874450;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163ecebaf72b58da7e0456492b0cde9ed8c526bf4d14393ffd82f7eea9b5f7b8763e379ec3b2d3fbc34bb1e1359207f3f0069d7edc41e6b72aa556fce2bee11476b3c7b8dcb096e867bb223746b7dc588ffc9e1b43d0e0ff8a66e6c046d8bb6ba69778bcce81cb5abf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3bfb84a47ce996f97f4e2f424b139287c7332e816ec2350e90253213717810a31c4a0aaa37b118dfff9940404d5c0ef233acdeb3095b27d12c22ea5b4c02c0ecd3ca3b64ba9130ca46b1f6657f30e252657ce28102a79178830083b5ab64b633029fd53fff45e089df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dfe705503b6ec77d1bd0bfa396a93eb0e91551cb7a142336b4f9c4f0f1ad827f7279794ce29fd9a228bdb8bff8a5553940be31544aa801ba921cf9544d5378477ee4a32172dfd2370342bd85e8d9f0b7a3075a9a1736c2659a2195fb60f6893c8eb22764ee29760032;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15758e124e2bb122a8d20a69f51d47575151793698d4dc2fc9f422460f3d269b281dff89f0e123434d8d44eb3f8eee3b57872f1f45974e22f87939d8941ed81f257268d9e2da1fe8be2a43730116b831d1c29a9fba92cff901207bfc8659890f01a986a3ddc864bf68f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1446a9fdd236a9f7ece83c937f65aa190c501403791750997442aa086eea81cf7798b14cfe32b2848bdd41c04793e329e64df29327fd6b004fbba52fe6e4c58a0404eda55f8d507b5b640d96c432a194ecf1611e7744ab83218e697d5ba33265535334d44ca34b5093f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14deaf219516642b7f1d7ca7ea8515cc71545794869ae70113ad040643be8eb6dc25a7c90515df2d6af06ff3835a8e39480cd57cfcb514171d900e6e9d5b25e4ba8c4b0f824bea3995e923ae268af5e55e2550214c2cf67715f25fbbff0f36a39f9ed12d6a4d16f9837;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f7fe40341c3647d4152c88da9f45a0a8f0238775177222b7d43e72ae84f0faf032118720fee1c71bf26c25bb9c9247dec2d9ff0d9fde3f6c505bf39fb580dffe6dc7ba45c7ae6c56fee8411ba093d82c41931997b23559f812ca5aa10f1b4e04a1026452d1054fe37d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ca9906ca689df7f39bfff45d1ac38509f28b95a78a79882b4ab279ef409c3c6492d8a61538996d1d77d7ea6dd85e82ca2cc9fdcfcd086f7dc9e713f1168a8e34a01fb45cce36654d56e70420d6c11e24e30831b723c6b0d56fd2911de6262305fd0ba0885ada1f15b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcc63a973f2be994fd0e13086e262918ff2fe7bac50f60c7e23184b9d56c8ebf583a4b8e45873d236e224c7538ade51a4a9ab51a0ed2648a1e411ee3b548656b72b8ddabc2d5cec629f21d7bd571af4c08251142eb662d344c3e15c5a7deac0eda53d55a877269ae603;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cf37045930923190227e257ad78e223ce993c6a49a58d21d55abbe11c96b420b72401f806620668e54fd746282733ee53b158acf8e58dce839d6a5341eb956268c404797bf558771bce5d87cd21b7295d896c56e61c00d884a693119ff768317c2d5fa439a75adc66f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h534c0655f8cb9d7e1956844c0c0a001d95b15d86b41c51b02bbb0e6ca77bdf1ad808dfc5789b8057fed728539aa8825c56175bb3d0d510e42fe8365331ed3476876c121d4968ebc21cbb3f197c62ba65531c1d76c08bd6284a6876c3ed9513d375d50f898f4a4c61ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heb77d9a28388d837890700553785be6f5d5a972fd5eacb0643bf923e8dc0b7567d383f2a9839134ba34357a4282ed49fa56b8dd5278b84c2ae6e511fc93d2b8d7fb5e2d4f5fdcb2e7325d926794eec3a0604c4adceaa66f6f113571a674d39116e7613379e8208757c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ee9f64a1d37237928a50f0a3c5e0323ee3841e24d4659bd4670c8aa83f2eb81e1c043c7c84a49526bd8c1c1eb4ea9fad5a26e780cf472c6ccd26443e009d4bec036596887d7691bb0d27db1d94250a19c1633020e387bfa48e507065bc66cb0b2059c96856936967d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ed8716d598842417fd8f5707003ea0b451ad5803d12af642d65792f56ad440452858d7937fc77e44978385d9376b33a3cddf1b69df696ff70744256c17a364f80934bbe2f218cbd5cf369f7770c94324c224f72c46a5c4aa38e89bc68b6f19954f51288c6268deb288;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h27ddfb8db20e18eadd6bfd426bf6243c5c3bb7c9f7fe1b0c0950fd75df252adb8897ef6a80b6e93938b0633478cdff367314347e4b22f61385338a4ef72e49a01145b42bb6ab1b5e0e140a7dfc9f910410c2bafd4e029fc2506c6ebdcedab5ceb17a3db9eff2342787;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6061a693b27373fc27d79b4b402d291edd5b87163e2604167af8adc570d497d39884a74dabdcd27e7673d70f07e6c59f214fd4452858cde54b1023b61867ad64e293fa34347f0e1410231f495bcbbec5689df15e50ae6dcd5ad931212da6c9ab14c5301304b284f052;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a57e0f63d245af22f6d3ac681c2f41b0e1079c35ff9d7183222253294b83832dc721000d3fea2507b421b26cd83a5dbd32c47630d5c00ae932d08ffb489e20c0fc89a02e96967c8f563e6f90637e4c308c1b3f3db27ae5f4bee91243d39a3a70e58eb8bd1914a363e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3b6a78fd5f7d022ca7afd94b896f7c7be0f00459da3e91eef29edbc0b12a6d04915c784bcc84a9ecab1934cd38f3a5e8311551799ff64c254ef0923d9d4375ae6d4a45914255a21640cf1a3a76563c12670b4335ad31cd2b1c48c1365972b8c2637876aba1af9e5b02;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf0d663680427a871958a7b2d247ff533dd735277dbaaa92ca14131c323819180b41d3cbfa92921f202aab00597ba2762a2cc1d32a34d36c7c87788bfbc716f8bdce470c760e7810a7ee9363d91197f9ef141864dc52841cbac19a2eeb35402a19c74f30231fa8c3e90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e1b6e80d741bb6e7e72cde13daba502f26aa7c4f203f660bf23f2b38b09b56f23e753606ed11e2a983e764987f1035f99e33bbc29b3514b652fd87e4c819dd4db53b02b81b4af905cabe89e142cc9b913b539f34e0b440e59b96d14ae58dffc9338281f005e0e9b10;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1227551b9e5a333cd6fd8a1be141bf9deed9747a93cd4e4c4a1da7e8e5cf45fce74550ca4765ff0bbf955eb10a27469a7a017ad8a4cf010b0023e89f3c431e2badd1ffdd5bbf4fdad081f708061090f46f9581463554ec1259c98dd840b649c0a3c8158a0fa2c72ea01;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfb8e0ef3c4d6f9fd488a296995709232ad122be5213e8c65bcacb2ce8dc531605b0a235492c5ecec89d56cef8fd9726886ef721a64c0ce74a434003fd7e8f1e89301e926e84ef19e288820a9e7b8352fb49c13a2afc51fde0d25c3223f8dee0730557395223e569ad3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1507b8034db0433b05fd6b863a55ea86ac898abfa79e005099b192e45c17b8663328a5fe62a9b8989d7ce1f718f8f44cfb09cc1e9dd8a737b7f466213221d932b4e30cb6113f996a0b3f25ab427736ade0f00f19b46e42728b6fa4a1d4b1fdb35269901bf1938b7de7d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11ddef141840bdc8b9cb6899d3324f5dc21be277b0eb71e608196918ce4ddbaec5d6fcd1ec3eedb2fb40d862183f38f7a38ffcd66740f53bf60d82abc8233fc9c90c15300021f127592aabfde3021aad73180b10cd7bb684b00acf141dc1d68f95f4e7b215c21d26e06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f57c7b5b0ac50406a90c908229eeb7d55c6d40ca96f9040f84753a09bf653ff842133a31a271b5645642a1b3f5a6f99dd9ff6158d2f2a706dbba437ef6d2942cf4e58d0174f22c7e60d565cc3a03cdd833b9ce4d029b376057db9315a32fe62aedfbc4a5188ff1ae1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0b02d569e3e938a4ca500a4828acfedbb987e54d51adc18eac190b9349e78804e5aa5d8ef7f77b91c00b0e9fc95dc875102769e54de39c66c6230e0a3e513000f41ce21c0ebbc316f64105b4d81a77dba883c116438754220ef1359e611c41ca11c0577e4da9cb793;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h28eed3437b9e3de01824ae349174b1e128549ac07769181b3187d7365012c2c9c35ca4b32f0a60a0b6d6c06cf149fb139c67c1a35a299a67ee55d511396effa6c44640fa726891620fad137de619011f1949ab81c434c827a219b6e36d413e19aea350f6e2354b3f66;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba39fdafcce029f0ebfe588f03dad1fd4a6c883e54e82742ff9aa0750181a11933c907e43b2e6f303be1b4156734454a3840183221ade24c9cfe73beab778588d23e9a14f2eabb894c91a5e4e7d9ec099cf31faf26f02d745d1955c89973f0fca615711427076ad2f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19ec48e9ec5a02293ae8585c219964e9c8f542ce529eead58bc65fd6acff6128e01561cc1618dbd2fe1d18b1a618c396bd1fc6ed8a7414b85733a41a477cdcc9a6dfbd9e9ebd8927ca55081e2092391847db22f0bcdd8f9993a5d28fc44fd3deba59263607b04aafe7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he8dd3dd1660ccfd3f1c5012caea411ccd55d3629a3518361ce3d98206743e8c4f25cef7033f4a822052d1be408cc27aec735dc61cdabaaaf09eb7a06baf133e3a342190ea9ac0b54ded2b4725b675a2ec47ec43ab20d36d985fb501e664e94c16c3804ae8b12970b05;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a7e26c0e49364a2c22e3194a8ecd972d6ef079444f924cb0b8ddd0de5dda0462556aadf666e686a6f4c753853064fcb36aa19dc3f970a4ba4582b95b87a7302d016d893940e69a96da438913a34797ec9514c17b8c6a55908b97c5d3e5124508460c7776536b6062c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17e5133434666ae8a15dadf292db7a2985f3922e2588cd5fd75b56c2d7e94b1bbcc5881a7afc8875987abbbca57ba05800231307efded83fe529649285e21f9825906561c64748c9a6d433947b5aeacf1344083d6b6afbde32b66f28fb0d310a83380bd96e5c287378f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0dc81ab1f1a8f219af6fb3bf82fc12756d60104e86ef314a2b842e69bf7bd686f15c25ba089c30c3c8525fd85a7d75700ce33daf83425d5296f8be935204125f9f1fd3af536407766050159a70dfb8f992377be99847248a751c9968d05c645c41b67c99fd519d736;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39c707276c26c185cecbe8f71f87e000206e8656048de3b403f4148c23fd02d8bc1bd5899aa4779d5b8930a7ee4bd54787ebab1b6323401673bc4d7c70a54313c9c6b7280b22f4c312efa079f2ccc1908ca2f34e6be88bc4871a5d8077e94a14aa8bb8b2985a444995;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h772f673752e4beff2933ee92476b09aac9f1a91f2ac5541ce5fd65ed750bd96fc560b33ba017575560495d0ae264032e5652161038e98db462e92cc9ac8fc0052c860547e9aab447227aefefba0e42ffc3ae320a00b69a42d8bdadaecb74b0ce864d7711f7ffcf254d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf40562b128e5192a184f20b3e69a53f215099c6602ac436d4f281e9a10920a6d8bc19986dea0937a3c66be549e560637096e4ed46ffcaa8649c643ced0585a33cb72d1937710cea1ed79af9d2f7358e3895f6c1e9a591a2d5a1437dea361eee540a94b337f2dcb771;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h26a46095fe49a2b03a9e07ab6788ee7605c1e46d1f1fb69ab3c109485e7470941279338ba06e5c2ebf256d27aa663628250d525776e21ffa7e82d49b7951f836237585c1fe00aceaf7c77d1e01177b7dd7b0bc023a55fe877bb1516822174dd8bc3553a8fe20be6db4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8d60743f32305707d7c936e74fd803cd5179963327dca7e1bf01c7985d4f66dc1df23416982afe9419edaee5526032c828613e70d8f3a6dbab70b99b12581744847477d7ba3a11d1511b687582c604f926e3623b300c5985f16a95b0b50f021713b00c8a5723f29863;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea47395b9acb82493bf1667e968c8a14623bcb11fe1a8992f596ddebce3131ddf7aa2d42726bb3e108cffa0d9ba3ae22b20fa8fc5c101136fc00479ddff1f8eed13ccd68f2b72c96fdb82e8cf0d75b83607e41d3d719efabb98af90bdd1f44e42f8c598dfe41e50998;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72ab6af731560b5936d2916664b56cccc59f167cfe25d12b6ce58cd53145659e1a8a1b8aabbdee544e2ad4ccd4de0bd98ea085c0946f3d91e3449d78021bb306a1e9b6ecd2a5cc52c8d713607d685c8bb250c140a5b07fbf709289fe5d29200103aa797d71343a5c90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1172ed6d9de7d549a9cebcbe25fee98a1a9e9edf9b297a3f9794b7b133e5488f98f903214b569d43535b35b4afd05131e0cfdd271fcecbdf9adbc892907a0d6d48b19632e5daa2baabf35e1027471d7c89c1e9f27c8854fbd07cc8115712bc46616b980de2677c30a81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c8f6fbb5127f410d01eccd20aaeb61db448304dce172a2e3503c4110267f8e31d2353bb7752441fd5c9634be0658cc37cb43b8414456b8c1f552e6553d7914d175b9079d3e6df8f126f5d6694d15f4cb4d4eecbea521d68337dad3e212c1175d26d7b75cb9672c5dba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc28fbbcf8e7cc3c5c356bac78485befd30cad934c712e472d3342231d4ecfd3b84b47a8f97b76a474eb6c81df6361f1b9a520e35273007d2a73bd2a5c2bf42b8d20621adbc52e8edd8f11ebf097a250c8f7a16c98dac5c5a73b556acd1d077b64da657424413d2de69;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15fee05eb898599dec8d28d19cec8c5a434d4141c1a3af42f7236cdef0f99b3af867615703cef166d98a6db8fc194b451cb32a8254ed5695b2f9dbf24496e8912f4a576613d251ccf5aed756a10955fc775a584a92212d11611f84ccec672bb0702f32ed31e2f2ed41a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15f7c936ae336653bc88f560c08da346fb2ed011b2da25728baf1d06bf06ddf2417accb69a28164d5415115fa5b890ca0818a4f0e2c8b54f1a5e20b1d72fbe15b75012ec78ab6842e53430fcff019aa7b39a80469ab8f44b3ad7d5927943d829722310c731443b5e353;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18040b5e71a16185c9bb29b127008dbf7013104cbc6f8e3fc3fb458ce4630c342052892ff06c6a0af6be4d6cbd305be30c1bbaacb5b317ce47f303fdceadfb978dea2f40ddc1337513019b0eeeade008f00f363eebc2f88912f0109284b4665414a1496c2403730271e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcec3672974177fb518958e2303c25f31d4864956243085d48629c62413a16a8f7f6074ad880f6b2cb4bbd40bdb5ff9f19f7bb45970ba4067048f09aad2c4ddbe17c397d8b3f077f17f544011e255a68ce8de3ac2585b6313735d09be574736d2c4c72538859d0ca09a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d7643de6130c308588fb58c38a9b486da6e9527ac31434b20926bc7088bf403e371de7f4f774853ba2f7f16640eb8143be17403c233fbc5457e3c6b6ab672a037b49f4a9a49bfe6aa836294009258fa18337ed756acaddb3936f27d8ebbef2ff7729c87caabf6c604;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fce845c1f20dcfa48e85b3bed3cdf09ab0011e24d906e15d8ad26609bde5aad1cc29bc321b9823c610dba64a79bcc0b85ae7541fbcb6ea9e137fda739e8bec9fe8137f6e5138f9a05d464490e153b7481bfb2eba383f7cb6ea81d4c278a2e062dcf52d78527259d213;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b1066ca44859f36007ddd8064ec9c25a49fbd04982ca72b4f2ca83868aa0945d94a98211e065f766ed36659cc3a9adb93da839fdced77d856b63a399a92ac6ac800c542d0cbc54dad9b1f3b501ffdc38b03634a47f8057c10c4a1dcf951745d304547bf269fee24e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfc505ca33109df4329df6d2fcaa0dcedd3cdab2c7b3de62f8001367e534d5f37219b5bfb0380b8efd1a1ad514e3b46b45a4f3aba5bc11e640a29a394563d2517af9358859eccb93b33cf874c7572ad121287ba5219ebe8fcf470ed74738fc11c1360b63b382d2be9aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha9e45c532770a96ba2aa1b8ed243ecf3e7c43ddb05cfee5d66761e34eff5abd800d16b54e8a281864cec4631579f2ef24cd57a136c1bd6fc242bde8d5641900bfdabda361bff3ab15995f3ec5e90e4c1918ab775f23600f4efab225bf267069b182bc9a71dc440dc44;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6f9b6a1dff9e70d2d010bc09ca743f4968ef0771cb420e90c5ab379a483131d4381f1717d25cdecdc94f3f3d7bfc530c590db33ed370056659cfa8fed2a42f67758b81359ea2f199efab4edc631b47bf07056523df6d2557718da8c074e81c546e15b3fbf82251226;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc224bfb691f77d18159d99af3f4356c701377ddbf3bc22895a4d72a1a0e56df72a130f3b9bf99aed352805b96587878ecc12a1cc8fe5521f26b76e69c7640a6ae440a4fe90d430d143294d5f99f3177ae0892d46ff547ac317a78fd637759a013d2dc850add52ef53;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19eab3e72ffe7c612e1081d4d428f60e3966787cbf4cfbe8061fbc5ac3f5dac8e7d79e6d5c0ebb9a95d465eeb983af93eb4000564119a753b22e39505869b73900ba4b1c3bc0940f244ff905e754ca713df2e871d44da589e9a644f1e2b59bf5ca743d6890cbaf77aa2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11007ebdae4920ad6f8fa66d5acde165f47b78b1e6a59ddeeebe39bb4b6b70297578757f30720b700dd81c14ae5ac2d85902fc72c093360f1851d83ebd3091309b6325000e1553d512ed728f79428bba8278714d1d0d471c873f69985de15fae23ef26312f6b21ca47c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he945c9d23092b2b851fad5a77e8e285cfa15087df3d7169ff5af97e7412e839c9471132e1141a05f0aebbb9fba7c9e45a54dee2641a62257383de80b2d1ea1f9a3382dc47a49f55d694e94f600521b40af8066c0fdf0f191d815c6a5c20bf51e93c38312eefd7531d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1991b37730f9fddfb14011cc87b0df8cfe53469b995a8064e38aae3ee3f01ea17118205febd234615ea6ea0ec46eee04cc62f6ce3df44902f0990f1c8d9c074badd4bdc72e88b2748a7e682f372d0cb44fa2530c78e4f8a96b91e9458f45b40be63f488ba2f54dcbe2a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1bb4a1671399743899a5744e39582dd799cc1ac2a72fc2193e9880e8ee805cd53d89aa3f16969ebabcc9bb012721e9f6c2a4f26afb2b0d7ac462c302f73af1c78745e6cd696ad77674cc3492728a85f6c597300b4be6e33ceac04a28de1a9d193ccf974ea237f815b43;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123b067e34a645b92822d2b1c929e24b826b95fbb0aa40bce4929cd4375f843e6c91c25da008c676a3ed42cd217c06720a7160110fc8fbef3629c121bce367a552886f677fd9f802bd1a73aaed76dd8142e8697482aabaa969141ab8b7c281a026bbeeb7a00569c5999;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43a0b2f85685994d466d0602d25c589f50000141c171957a8f68c02601ca40aa3aa49382f6c6345d4cdd61aae75988599705974a47ecbee56f45e7a77b4083d7992daf189296bc1c2665bfa9d119105c3158f9c85e56ea26fb75750e6a6b2bd1940e45b2b60d64644f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7eb90874a1300d5dabbb807f62ba3408b3092d46610d649ce1e781312a9f32e05a0845001f13b801e729a9a8df52d77faed86f135bd12b6894d99b850963ea1786c0951db0aabd7998d52cb128611418d56609e27c30de9e8128bfd337080e111ee76ae78ed6252249;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha347f9411c1419d20222844aca8062a9c50444866bbe4a907e51676c1c9a13df93ecb5b39e0249135ec5c048c82892daf9c253e5c9b4dcb6f2e1c699881bc7244b2ea4ecd8b8d3e4e6db4b59dc7d59290ed50af0eed63bb55929cbfe5555fec93ca8a09b0602254fbf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h652067ff0a7a8a9416755a1e50d43666ef25dcdb5ffa6e9dea3bfcd7c25a99e5247fe942cdf8ab58f84adee5e31b6c9296b3d7711201672a1fe1d3e576c819b87b2f0a023a8c0643c317519a579b59f4397d1243f4f33624430a926246f4a8552b6593815638abc66f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13419a010e42641ae19f19c57dc48f8ef34c8cf8e4615919e9b9b4dd16817ddfd7b028a933e2569fca10abe134c0633436ac5709f323f9d6e6a7f9a8ea88422d39a545bba1e4b32907aa234848a01e27b2d4b0d02688e8480a94bba77ea2d60000a697ad60ae300ea1b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19437fbcee6f33df4b16d879a4a7d3a89587f0b77d8fb8a44e5ce4d8d712776e884ff407ce484fc2eebe3077ea75caad4242fedd7b091340d5896322aec411e8ee09b17e0773e36a0cae0f3936333381fd6a4c2f4f189235e29d67945fcb5f89d71cf4a2f09f41411a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8db4de6a8fa0154fea38cb176afefe90070931c53ea51d7af9a2b24984f6b128a906f34bf38e7090f0f2d8978ede77e85da4daa79ec52ed89bebbcaaa39a486b982adbe7404e22e1e84395f9890a726b62869f22158f28e3e40131633c249679386ac38082f8837f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e8a47adfea6ced08e8b7d6a43b57c85d757e9a64dc45ce2518b5c2b4742c26f48fe811d4531a9719d11a9c7a1e79cbe4271a09c14a1b727453030fad8e7dc521f8dcb8e65f9c138a4d58d65b399098c249d3f12cf3d08c0f3b9e080ec766964d6b5ff7e8e6214c4b7e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e25614bf70381f9e95d962420c042001cbba25c721924d3f3016b490492c13e2a8f0a78a307b110906828b48ca0cf8bcea530a73c9278a74e65f50070ce3019a19b6576d3d064b3593ad4db055f7dcf3dd681985ffa1aa2fe617fe7621e265f167d95b6ee8d77615e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h496938953bae998129e37775dd72e481f0c6d6c446688238ea15555a0a2ad11ecb9a3dedd07eca09dd7ddb538248baa98d94e001bad40d002e9da01b80104f377c568e961f1bf8a847d16abf5f60fa19e26021df556cbc4eb71406528b624666e7fb5ae8ba033d934c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb2f39ae6b6e280a049e603730815d2811831843ee649c0517078562b7549269705646299878083f624c56a96d892cb7705a1c6b7f979d13e77a9f5f629f4612d21927e5bbce52e725aa51a9d3ace2448a8826ddb1cfb38d2f7dc5d65b6c621908a9c45e854d820d9b2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h813f3cb2a408362f8b257e77e3dfafb434ce37eab1bfa1827e6f30f071ecb9aeca0d6fe483488f7a18ec7db0ea246bfa77621f3da10d7848fb4a74fb7074cc9fe25716fe2cbe1312e7f436edea0a13bac44d239aef36e07734362b9f1fca7d40c02377e478bffa37cc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13c54ed533988ab876fb69851e7f5175b1d82fa28fde7959be1b4b1b7320034fa15b81e1f56b9438529cd017d5af45322073dfdb48389487d600cef55d9ed15cbe08bec60b47830ceea34832d53d96119ceaa86a0b496da28c7dc04c523f144685d84dfd87c88fc6c95;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heaedf0fbece7dd452a83c41f682ed4c4cd165ca61dacbb5e1388178938a402afb083886aa421594fd3ec594e889fd1b19dfa30930b37c150be2a1082cc5aa4eb3abda5808a391eb4b20039ba3e6909eeeb4f3102645f7f50732b06e4cdfda1885535d5d8d1f2886ced;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10797f4eb4234998c31a917a0d3b2ce06725fd3b32801b5ac4c8fda3d2975491ea340f5b7067e5fe0141a10fd543a27c7c77382c8dcd73fa03478daf74f03e2f6efb03bb3241963627e27bcf097216d3e983062eb0895ce84b2c0612d3968b25963b62a8e485f84eb4b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1980e20d57c5ad614b8d087b782206e9b6a9a89dc639090731360834183c0aab2060a1a1e1441cb24948a843f1b98428b3735f3a62eca0297efef8e86ef11ee4920f6592eba63a1a3a5993008373d949d0a093a1326e752b63eb6f2e217181382654a80b4774d5b3dfa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18f46a09bf140992fe22709e2ad026c7b812b5b2ee4f477335a581cd0f3f2a54e7a252cdd3e7b09efb1b3c2d6b28874549ca25fd29a6ee41a8ca1cf1e251d1012d717d6379fa054206d1c517bf031cfa26b73011844deff8e692488f74faf476b575a9ba9c9892c2df8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b53a15fd425ad37a78685011a6b1893b82ec440638c910e86d69cd588ca591f06bddb1e15568bc7c6e70a57f434254a8bc24fef78bf86009afcb1e489815f8a2456f525f5e5bf2c0f954df4540eafb48ecd999d8a6b1bec4d25cfb6aecfaca3be7c7384ba829e25fc0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1967fa0fcb4094ae3a6b3258871893b36b91c5850df554238e6ba394d50c4b9be6b894d6f4425d637df09a9e97edc4ca82367101058ce00631e4d6c2a41f861d2149a8f72d72e2f0e134fda9cf4095d64170190df2a009167c58479ae99299333dd9f7adaf97bc1ce62;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h82f5824f0eab459e1327e54c61422b2a3bd027e78d63d413dca7b788315a22485b0317208cddf96731c8f40dacb45c760acc62513ee56dd8723376f6f7584850dab135f46a19b1079aa8ddc73b6ceebea2ccf098110afe1052d76e5cc0df62428b0b269e72b8752732;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67d8b752e0788b65c400c1ad7e34e5b75b318877e36ec2c4c159711554a64ace05b197b2e20f75b03ecaf13c60e23ba68a5805f1a9166268381b93c1450cbd9917c7d08086bd6cb2e855bbee43ddb128d8b696b28657ad8c721c0910a5340dc7f94892eb92da87e214;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1203fb9c4c463682e98c046f9a0f186d923317ae8e2245f47f9dc5b6a9e7484b47b5a88ce79bb7c73acbbde1950c1a8fbefd0394c0733988fdfbc515d6ba7873acde96959e76e41d5b5f2deba71787cb10937cf2a7c789536a22b0be271e20b1816d78c61d003bbff01;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10b994c0aa73b65a944bc6e665245d272009d891bde07b187d26733b14561c2d65301a83985b8be95b64c63d2f4f73bf265620ab9434e94e928e7d1f45324217454a739521c1d594d7c96a38d606881fabfb9279477838b0c1ed49754ae427beb4c8df3c42e405f9cba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb9ffb75924f0ccfd537e716ea2e3ad7e91e49d73637221fd1674e5cb74e675bcaab7fba8aac1fb28e974efae3266090b166ba979874c4eaed3b30c2aabb9453ced52d7477e970e3d583dae6a55f6313414b1ab6ae42e4ec11421e059d6cd47bca1bb3c62cf612b2d3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7faa20d9aa3c113b34a2cbb6c0d432931a45223e0748dfcae065d10cc74873ced67deb8ecde592ce1dfbf848d0ed48fa1ee69261e9777654e1f5dd61dd65dd3391a072d11971d5abacafeb03211a217753742f5ef9d292d5d2d80166b278b58bb19917d0f3b1f9331b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1258c8af0183dcf0a5114e7da317a3da758dab6c6cd4cc2672f4934ac8dbdb1a5aec5b7f790b6cdd46fe1269aa662f4e5551b8c7e6882184748aa245a18bc8e8d09894c8ff5c4b2deed51dbcc24285dc97173588adb77524f141300dce9de3ccbf47483db4cb10d46f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d0c5dbad7c1b70f0d5cb56a72b93f16d9dfd58944903e7be656f8a9df853546104b4d71016fd6414821638cc7024e10cb18d437bb586d33d6e0af3f36edf66130c4c6281f7b17ed4c21ce0fbda76f7c045d5c8aeb13231add5b111b088ca8abd7e87c52a3a27086ddd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1790861cd5b2a577a7fe8c767c331eb1815005c50353c590dc2eee66bf3c8300b05a8bc0223822771b879ad9e1ed37a3ce3362ae56477c1c8a950c79d40471eab53e6a2ce8e897f746c70ff3662d7dc95d369e20ccc545e6d9657201b2bae150323d260a5db3f792c2f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hce4eacd10e1ce6b2b3d1baf2f76a7fd46e9220e17d2927f1640d703b3f5bd8e76e162ade5c19c2516c7c2821e8b7a5c7d40f69e248e028178ae01ded28b473a6e82ae9221fc0f965b7d45949c21ac4af132b2e9538e8cbdf9b0cd0286ffb583c5ba19ba5bb9055968f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163bd775ba4f20771f2f0d163936eb6f82e97aab698e8b0df9c5641d098f3cf47525a69b7a13a1d7290da4de57aeb671cce3ec73905ab256b8103b77f84e9959ca9358198381eddff09c6114419e5b3145adda776f1639038392c2f32615711118b69b79dfe805c0589;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72a557b9cddb2297953f70f2430128abf83fb4f74e88ef953ee7f2a9c1db7d86fe71095688478cd0914834a526f8bd62fec920f41fa36c38d17cfd573939aeebfa873b1bc67182846244a5a941a4155de36fa8a2ef6e83de1868ff21e44d944be6e70bd45185475bbe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10ede1ccf4e83fa00f8c6f772c9894f85abf3d1774f6da6bd1ee731283f876e5539125cfc3682c86cee81e3dc11b8c2bb1a4c1cccaaada509f440a1b2ee7d304fa2604fd6221e312289d878d5eba0c61d72bd3fc226c1ad0f34603438605f33fc4d7a47181051f1211c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h939236a08507cb401a75ec67afa115d3b427fabf0cbae7d0d47a3c0d191d235e89317d9a64f332018c8c407f172affab953a8445ca464fed956296e68ebd15dfbd280bbb6c9fd2eeac337e4fb100b18f9b030efc2e948f8f84607966e49aaddc7bf2096899b9e7d9dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'heea09352bb44827fb0a5a42289053309215e13910b67273317272e9920e23c177433c0ec4b777b5ffeb44a3d365cde2529daaf20c25c220da92eaad4ae58c7286d2d0e5c1d95d0e81e3e7c0e6683a8424c752cc79e28df86f0c720f8513c85b865a2874f3ccee7e042;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e88b6f9db873822286c05a3c25ea5991e9e89d6fe5254cddf0115838d5cc8fb22f1c52fb0e5899b2c16168ea026fbb9fca6cddaa05ae4ef7fee54900aa62ca93ba901ca6febe895534b606a2e0cf9bd78ebc76b90bdf013315dc7c3229919bafd5af4191f550549e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17a687fa7ad0527fcc52e9d766435f2e404d9207d2b87f43aa847b4990c531f7002685fa80ec06f2cb9b1bb8f75205bd0ee86564eebc90df45424ef158c163d20ad97e9c7819b7b9588b4e1d7e95f96fc9d9f70f2af9fc0f0f663ef5b5646e4d2e617a09169ab6e488f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba717b2ff23fe02e1755c055a9c997717153cb9d726b468e0ec3252eddbbead6de905c3a94ec38aa7fc104f60564fe70d60aca3c211292055a5e620ebe4952bd0d81df3cda7ce7cab02f144d679e352b0b7162a7e681c2da273da36cfb66caa24686be1e8493f910fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16b56d32526cbd3c90a00bd098e3870e3dd488d9daa4b93dc43c95947e3560dda2fdfe6649f98d17962728bf3db87a4e8b1ab61cdeaf0167760e7ebe588b6af17ea7cf117bf0fd80f1caf9144801d218b34c6feb5a6778eb02b350d229d04f1810d3c661163a0bc34de;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161e67c4b0c9a703b7c800dba6218260189970ec66ba86790db3b7597d7c88ca3f8088b6a4b200c10017d45a890be5538f18dbe8a23be0302213ce23016a09223f0c92111fd25ff0cf6dd92b918a143c961e9ade9ea03895a63dc978dbe1efba3c79ae2e3f530a44b51;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4e036cc14f49a9e797f100a0b0eb308c5283a01de5ff2a0e5e34190693c6384ce0e75afbce68f3895f1862bb289e4c439afca80e49770a13c35f4c50ef04a6d443e4e48329a13f6383c9e43bc6e4ca69fc68b0b033657c6feda9b49e40b2c2caf52d4b1968d4099337;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148eae594ed44c00d3a111b7099ced37b101bdacd0faa113ecbab023e41b87afabdf44f969e840b7d4588761b9cfa2b6694fc09e92db1575f9cf8e3bfdb4574d775f2e751362647c166420696283efd23769d621afcef547a4595f87d8dff943a0c5b28e0e5fffdeca6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4b8eada22f9ce7b6c178f09bf90ad1b8602d53708b5d65dec8442a845aa78bd3507b0b718e674a7d9db1602fc4922d776eb63d432a0a474c204b6e422fe68765f407f06c4e695251a490623167a184b6b2d2aeb2844384a5ccf2aaf3a82de67a759ef0cb55fe9e08e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f73d10f6cd4df27d4e8ada3eb390278fff0b3df1f2de0846fe7bc0a785eae54caa20c34181399090700fbbfe123b7229da0723de91a34c55af74755d9cf367e1c6a17373238ee3411dca32c5b7427a967b25e1e6f4e87350845e906412cfc8155a9f3690fb6ceb523b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d082d944201251f055775f1ce796a4d41872f6d883fcdd51a0bb788caed7bc523db39d942415b3159f0bd54cfbac7a78e68acf1cf2ec9a04ff4e7dfde3a57d4e59ec166532dcf59f5c56f8d232ec1b5580837bb33aa2be02000efcb1c51e88ba8e6be2875841d706f7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h69630d48312bca4f1c76403b6bee03acfd0bce836b4a0dc389a6c3708c9bccfd54e80218b3ba0aefcd7f49b11b23ba5770c5ec5f3614e5a7d06000148baae99a721d79686c3c8e1d21c9cacd77fddf1a527e0cd0a09468cc5c8a55254b47ca500a82a0f360cb080539;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5922a5e9a570d250394bd0706a2276a500e714f49ba8a801f4a5d1f43402ffb5139b31969cf14c5de202059c829fd170fb4d02ae20600518c4682f12dfaf2c83553ccf35e673f69cd74e4c66c7b9f98ec3788beb4bb8ec993c443ad54fcb523b5e0716026d851d242;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h72ad1eb1e55080126053a81483935e1ed582402de62a1eb3c5229be02c0ae1acfc08f238d722f67a9f80f5ccef98d1d6a65964aea9b341626d3041a4a2a4aeb6ed3a3daf2fd1f5a9ab940e030a22c9546b6191696ec7abbc6aadc64a727deae1384a840ccc56338d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126a71e2d6e19f2270a6bdb1837de07ecd618fcd265ddc95e091f82d29855d3340ab07c21e871fb4acd3cd58215c2cbf00402b6ee8cffb4cab7e74b5905513924d5e0d6216f096697f4aef376b296432357a9dd95c97a4385757b4e07d7af0971a40a2f2266baa08d21;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a3c0f152f8aa585150e317f18f72b1cf7cf432bc8dd3aeda660b47bed6bfb209c68ef5133fb249b1944cb16cef2d5ef0a1ab5280a5021d83ac8b243c34f8f1fc1e50bc3fa37e8aa3d083d9b026137a6e0ae0ce9ca3f817130838b90e64caae94b96df46725cb78f15;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15127693beb8db52dd12e86a0a918f2768d4354f5f0372911b08fbd8b9108f9ff0edf1bdb80152027efe69a92345686b571c8d701121ba066bebc7c3d033b8c078ef647b0eb2c372e09364aa34e85f6a7dfaccc6ac2bac704f2a2b631f043d4956b56ee0a89388bc1fe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe39288d3ae0b363f0bf10576cf67b13a9f72f1edcd4d0118a5a898955b117a40b23cb56ac6144a8f24bf93964bf189aec5c7b9682b55dd9ed2c80cee27e0197c750fa67e86be9b56cb8ea9365e96307902ccc2d215f34d27902e8bbf60f1d681b2855207c96a6b130;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbf58bc3f9b62719e40d705b864d2ab20fbffcfc7629d3d423e96376ad2ef4d3d9d02653dca75eb587980bec5137732ce769937a965341430c69856bb1bf496ef229472b508032a6b04f0cd543bf46f13d8f4f24636abc3ce2ef2d774ec9643ab88815a085f46cf76c2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc44cb6cb7072907a6585a9d56bdc1b831990f88b0172bb6faadd6579879ef0ca14b1a78392f0b8339993e4b73a206b8f253aeced24c82ab2ab6cafc1c3bc19b0032488f02ac33bf9547aff7dbc40e62bfc91aafc23684e067724d55a6fa355daf572bb2d671215055;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h947ff50b9c1b56cbb1d8030c6174cfc5ffcd5ca65d025a54590a1a0876a10d9f19ddee155f9b75402888f158d99a0691f63c9207c84d83f637d3b93c4129964c69d7ba8b9671eee36d19a0acc74aa9f66210356fc6abbec64ca9d8acdfa8e77eee9a44d95ea19f1243;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a8ff674a57665dd6764d0518fabc585ef00f36bbbf7a3c0e53dbbcfd81ec06c2ee9ae57d1323ba6adae00ea5060839fbb8f9e68d059bc390c9059724b7b34df9ff523761740470326ddd3ac41212b7636caef265db3392c087dd19c9ac4499d2bf7546a620e35443e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7371eaeac208ffbc066a3f2663dacf0cc7b7ac28873c6022aeda7f7f907a030ef22fd6977634e838aa27217606d08b508134509a91c15661970b5f3ab62a31850f61993d3bd7d84c81dad0e2b55482d1516e7bc91a6c61a71639573a14f54dc031337ee920fd34f1ab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16cdd2b9cb2aa8d22bb711003c72e51937cc5179459d5493b976798333466868e039da2e261bcd9724987a7e5b7b417b4ea31a6ee896ba6254496ad3febc582be0d6732f70b4ebcde9f06295f72c2bb68e13003665ca7531db4700a6624d8bbcb226df9198a9a8b4a04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19322802129891e0af242e96d24ca3e519d7c640bf48c638d138b322cf5423c88d91ed9ecb416d33ab1da17cfba0aa43e6dfddb8722823b79a88a12d97b2255cad7b2fe1a570e1297766dddd7c772c7ff02cde5b83de9047dd7ca70adedd21ca258472729889bc3fba6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16e341f21bc0d14c674796d7edd0ca4e98e2d743e3f31e624462cde3ef152580bfb674815af7da8eb8f0ff3b6ae7409cb070ec3feadbf776603549b845dce0adfb0da85bc102c653819581c3cd7d70cbdfc975246fbe2922c4a705f384328e8e58801327a2734d3270d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h21737d68ed7ee87349720d0618a1d615426d6fb1a12bc6b900b4f9296ca40a21e67e1cec2a2e45f10892faee6203f5363c170fe1fb46be9512c04d9a8b0012f53fbe5497ca8b32a5d8e7fe16523f6f3477cdd7157001e39c8fe80d7383ba9854bcd384779700002c46;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hca5274ca0ae13edab28c422ff0a12b5a0e6a0dcc3f41146986d8a77a3debcc39a764149df2ff36a3cca22f570acae83a083e91707efc9585bbeb06239038a511c4e6452c0ab7e40d582927790f427c52ba595507ba55823bb428ec9c4ee158e34857f40e6c713a899;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a5e333a7073ac6eeb42875145a66097bb58ed1edf925040b889850743e4fa531800758efe3d6bba5b89e6ed4c131160e502e26f403497158b129b7b8435f20369c504b92ae9b3f32d699e11e1c74cdba943ae0a6505a2d18b53c351f32e58a637dcc3916ef1bca0ad2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14a48dd51f55e70a2484cb5c3d5e17a5e6a45dbf4977ed2c5d7ac4cbfd05dd4cdf8c5909ea17eb7cd0a0f27b547ecb507c133fea656737aa92304b3e831ed321b13a535b1378f95ec99a7a73be3d329f3bdd2fbb556ddea3ce12f803ac9a7d825fb7f79c713a8812655;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h108eb928291c17f2069ca66f0b5fae48194043cb7594fe3b70370e37ab352444fafcd71de54332ceda05f1835e285fa51c8de22b8ab94688c4344aab68e4062f5ed53aaed24c37bdedaaa0e3dffb82a4ef91b068e0b25923e6b36f5a04a69aa42505145bd2516a5aad;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4f27c6358a59db49324d475b283045d1489dabba040ed743dc6607573f80863230e1cdf922810d99bb62b54a55d7821f38d87e928b710e41e404fe9edf2d9055ef1209569479ee92614fd5288a1f9084aaf8d8d92bcbc29b103f74c0cb83eb361090ecec579ef494b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd354e50a148045d70b111aa5626385beaa6f0c231b83bf3c7fd08bb66445b36bec3ac38032d8023a7a58312417cac9d53e92a12e8843209b6f9afba26da046eca2d65be47b92c6653ff8676bd20c3e73c46ed2bbfa699ea2f7492a9f861e5f3c5ac6641296594b6a2a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143a6993e138efe67d5e9a76e744e8e3415dc70317ea64812c382d2c95b2a3d3f1f395a07269e882efa265c46f52e0992714d264801fbc5ade8e2fa1156c3ea513fc243cd2de7046221cd97ab06cdbb7b39cbd135a3c34fa2b49f6999e098af083c3419598c17c26720;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha0412689d5aa8588271b236c79e2f83f4df78924c513d713a2027c02b885bf4816026a63df0692737edd1001a9053b624524f05deffb23c403f965a45915f52062cb93a88194a4672cf37da70e608aa5eafba913be9d8b5f54ad0596a3de156010658e1d24b4022ba5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h64f73d267a0308b65529b0ca9e3c3ec53352110e5c6b270779a25ab67a78113bde1c75bb0632a439819648a1e70fc9851bf3bb01ac5cedc7463c1bd5f2cc85697cac8b53f20bd7d17d48d3a9b27006c95ce72b55bf7214b7c5d70cb02a6de6f9213f44f8fc83d497ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6c18fae4d954f1f5c9e65cce62e82cb35c55b2626f847e82a7bc5c47d2f3c16812c50df99cbaf7c60e67a2a77ec6a5168991049c5642698959a853dc216aade21fec479754ab1c108428c6ef924a51901f3169ad64237eef5bdf5ba080dc23f19285b57586f9ec0375;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e90df96f5ef2438dc26c10a22ff2859b6c850f7a8975da909dd3e3fc0a87ca04a0ed70b76827f2aa3328d5c24ee4602e4a203ea7b079a4ec0da5cc37e83f307c12f3f0283beaab838a75ce6cd5e90e8e52f54b74a507252c357e4baa163f40b5664d7dfe55a84e9d2b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c0416153efa06efc72e3017166df669f5ec9bed5e05b042c1a031b951ef719b2b198c329c4f8fc3db88d60d1019a0bae8bff5b188e75441941282310bab5f8cad532be29c20f5ccc18c32596294909b5b753d95de8c2964269db60aed130445f43fe12beda45a3663c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11463e08a4b8dabb4a26c22737328d2335691a0cfc30984c09ffc7cd951a313cbd567d0140fb860d999e523f4a0cbfe30dd434cfe4225fc44bb9d8b2dbd1cd367e4e021547450f2d176d4c67ab29f6200b2d62bf01df419878e3ca4940d311c749626ee151352135a40;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h99f36cbb19f5dab48ee0974e627ef58c74adfb74403681d59a96b0f4ef20f0aeca3f289cb5fd112395ab658c3a49f2332729419e578706178d6576776036148c7af2d0eb653258fc44b31dcdfc54c065dea87f7f174e7303d139191bb502cb6d156095da14305ff5ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f880442ed1ef13a2d7d914ec4d32adb878599cb51a5e8b9e25cc87b889ab9e94b572ddc0226f2ec0fa77e0685dd60f595d0066b94fb61d7b5dc66de25c4e893b5037e5454cc10e6da7e899ebd049cc3359e5ec961a07990e943f6f9a497470ffa0bad22e7f2a2864a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h62ba51eb370eb87c5e78130ee9f86fae134609bdd6b85f155681bc642907023eccd3b6571efaf289eb58f0ca120c78e4b1b83347cc869e02e391e479d7e1f45a50a3c8b023cd5913efb7a562a90cd3540a92ddace0f1520374b618baf8de87179be2985031c604a1d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1555f5f5fd10c8ca4c316e59cca0c26bb69a179a6da8f6c5dc4aa96aa24519d8cd6b222a2f227d3bb237227623fbe13cac88420b62c7cd21f2bbe1e9b62312c979adfa15956d01b955e4819776b86b8dac58a564bc03de726a6ccc0304c15c75fa6665a9e2aa5f2805b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ac93631386087e274b5fc59c7ceb36ceb2b77dae3e2ddb3d675eb090cbf2b6c3efa886faf903669badc927ed219d1ccb84ddc2c89a0add50935202769bb4b1cb7404c1cc06854549e7d289a07655b28f771d0a9bedc7d52af169e0efb256017812ffe1bf34593e90;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfa451ad093cd7cd36410d6867d56ec5033d970ee08e7a980cfc340bced32ee7aa126da826e6cf819108390df7da0b14aaae73b056fb04d9dff44c88c7c7e40228acb54c756987155eba1f82502ca9a8aaa14096da54c013292e400fca365d28f7c1fffee346813408d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h101490b6ca553b22387240eb052ff1b8f98d11b1626a816525ad058258ab449bbcb319ed8f781bb90b80474a0f9d3c2ee84bb8ecf1f6d32df28decc652d63f632b98d5c2a27a8ff36fd0931c4ae71da315ce8a867b631e292cde8d589e5e1bfc6698477ef36643938e3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1196abc4b9d2abbd1f7a3a3761b9402d437c1cc0638a8c041d787aa557aab8a0c01e4b9372a2e89b2f7380e49429ea044d193f5c4ab10ac48b2e1ec73484967012f9be3625306162d4b3d094fea085c2ee4c9ebdf22df1ad4a81d3d47dcf3d32ed4c52f8193f4680f88;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdbc2bf26105c49b15dd254ba8216b58c94f93180bfbe29d3c58155a5eb0db49e99e8bebb8f860c9346fd1a6f5244b68e70cb4bbe5f1f035126f9f5a57132c76299e104422f9f8993f90af72232741e7ccf3931813b388dca2b519d8343ca2358b917a83342e2169ae9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7a3bef2e02099e633e75673bee857d19c8551c8fd179ba51c3211207b6ef7d5ee5d5c697df47f68cc1fc801e2d1882baa763d63e95929d58813957f3395fa81e4e1f84d0a18511af721f1a6eb30df339613b88041b8403bc58f6b060e6a28b11c3b69f624fc9eee3ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcbed92302ee5d5ad0c8025ee43c2ed768be8ff79a8ebc48bdb2eb2575263595349f64a46109c877fceeaf93898189893b31802c6f6427419553967e9c5cc9d86101482d6bcd4204847d2a3552b833125a5724f1ce4588d0fcf68722a295f0e0a04d3e02d6846aa2ad6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e7713ef32e2f95cd6554251282f0691f9515cf1947e895d53b6fcf0148881eaf91a9ee43a972d1bc89e4684aa5d8c75abab1603c8980f11692dea92cdfdcabad7081420c1123a2cca6ec17cef205d1218ae4915b97c39efb65a48dc4ad6616f4c9a1e5a70223a2216d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h40197614d7c79bf41b69a896ae0b5074c7ea0783d36547d0bb13a9c1966080c40b90ba0cb03dc58854c6cf0b20b37e23a7af76b3390b70dcbb7b3cc557637d05853d7e2146df33af40803854834d5637d9d477acbabef649380377bbf9837b004ced8750721d70bd99;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd46be1fa08ce4e8a604eae5d295c053adb18aa65957a889a25d0e15898bc217b0fe92ff233a43e01643f40453cf769eec998b4e3c7b254ad08d3321236fddfbbd52064ac67ea0e55829719fb52cc11798fe853099230d52d763ec9a133fc77e32ac6acd9718d9e2fa7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h197903a63d593265edd56d24a0a18f9a189419190d262b445d54cf6fe10db9e0723d1df45bd61874c5c9cf13866c56f907c5dd9eda18e004d2ff1d6a46c9ade582c98d48938e8b22a4ee9d456b6f6b117ed54c06fe460bf326223a5de7053f7103a6b30e29fae37bf8e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13582b81a78dd3d18b2914863d9b0e02709c28c921ecb84da3597d1935ec743ee1b171f840585d3e8574895824c1d814da65f5c31e21d4c5666d114a418ae2d93bdf75662a13eb56f2bdb19db8dfda5b34f5a2998ebe9eced961645c488500f04e33560f5e870f78263;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c5a926155a537a274c675279b40af699f9afdb7771ca27b26136b9167c36a4976023750f26d29f8518e82f9b1046c09d6405981b85979d919c31824d6b7237f40fda5193938dc43b77d8260b749fb8b7b265349746235425d39469e6b2f583086c31844b298148b654;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4297d9901512cf014b42eabac2302946c38e396c2da149879d65c6253be3624fa61501c962ac98801584c530900d365a89545055336745f079a908595e9f3173e17f128b69fb8a777a01772260a3c30410ad88cbd4f54c1e4b6cf8cb3c48fee9cacb2b40ed5ba1dd06;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4dd27c44537601f6d5dd375f416efdb2c19bb731157acd38bc2fbb677bcb19200d93e98eef06e1f136def6f93ac3f505677b1d31c43e823a92b9bc8065cf338a8c18e4a207ac7607437b49ea2b967bea405745f4fc02171d5a3a9a841b0b831ed1f53ec9e9603c547d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d35d83f53502232c8bb51808c16e4bd9e830c44d596c6db56eb1a88f67c845e30e485091369877f7ae756739d8e967547c0fc0039008bb88b3e71e47a6ee1f1a144474a2fe37ad5ffafde740ade6ebf35c941588bff5d1b3188066c83ae0597a690319ca6cef7e53f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10bb2940d8b024a510cbc5634b53fb24df2a54c6c04a15f2cd35cf282e46ff530d0c13f7cc9938d67b9ed2f78ab72f176151bea5ee1b2ab000b461bec70b84109570938eb7bdb8f7cba15cbdce4924fc834060db7bf7a301c50a92573bf596939df7d654f65c9d384b9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1132137a675dd6d57e928888f1b469f95f06b89e19fdf8272e875948d6b650144c3441adc805f75965cdd0792f5a6fe4bba53bdb72dc420145250135b85110bd2d08311ea130d22030873b2e69c6395e622ac20bcef267f6b21a5882249fe0e75bf1488de1f9d75ecd4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ca1987f0fe56d73ff8e0e28e10081ecb4bf93a0693ec3cbc7af2f085c25b141f62a7a5476126d45e1dec14efbb779b258c49c0febbab12d286cf908cbf1c93a78302071259955a8d5138d619d4772c5243f33ce42b5d6e4a7b32dd5ec9f58fcad6764b690f169baf1e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126724060f8dc41f27a53377d1c811073d42f04429c1062e5b42a67333101c0026642f035c0e2b1bab53b28af8e8a0a905bcfad05a1e0a66759a53912001cb94609aac990a22be8d3ca9f0d5c8b644db06148942eb38348f945e0b9afc7986c30affdcba3a76d3d7cc0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1de7d43090350fa39a7617e3995a7328d2f0e0fb437340830fc43f04ef6b1132f99421ac5e812600fcd4c21e9dc1cade89cac6f9bbe1dad6e6c90621bac7aa528d662ea05284264a30a8ab04dc78f7be15f0079473a3e9f893591b05dd8441daf7aa941efc3a1d6a679;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f620d5dbe6f81b08c74d660d71556c7b44f1179c3dcfe162c605b36b5c7857d1b18452aaeb0ee44f154e2494bb5ec640e57aa6edb910640c06a45f09e19ac63b51fe2d564ffee509d7d7a885e00ecccaf11e4c18303534d92201350dd082b13d88302d70f3ec1c7edd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13cbaab560070ce9ddf919e0e903d46fdfe7fbe3fe2c063d2e8324c6879b0c1baf7d8c81de23166096f8a8c3fe0fb0a01711a54656946712f102993a36da531681c29aef0665a67c92933119a653168b835c20afd135d4a93c7d54689e8e05ce0ae0bd0f85c38b00256;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d9303360e53b7b8ea1bb3c068117e16d6de87f8b75c2d82f4c52588ae1b3afcbaed0798c45291f5a399ae6001249d4327138b2f939c9836743487306e3fbbc6447fbc7468c8169ada0511d6587db807fddcceed734ee573d7500d35fbd12c4ac15a99c12fa91ae70c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hde012c50af06321f9ca7d732a4ca19e628654f74b88271f77cbfb8cc10f49249a320f5ae69259e3d47e5aa4ee8e1cb32f69c6f7fe7c3b609a91001c32f5f12b1e6956473e803ac0662a203e8133d650d3d69931ab8f3800ae55355bf7ab4a8145f20649661a6c36466;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8b0ebf79234bdbf8dc3c097799c6ed1e3f6fa724124e263e4f5564d1ccd3d5207f6a02a702767747bdd25e456a4cfaebd194f699723af0d5453521f379dbf83fca87f72f4de9eeaa1ac79f97247fc1810513b30b0799701aed48155da6447b57a55ceb3e9bd677235b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0c84f917a3f96fbf4006a3f385c00302214a7f410880371eb8942f22688428294ffdf0848b45fb2ec402e2161d6acdbce346676218544d492282e437837d2f29bb7baabfb664d53a08a569d7ced3eecf3a40692d81b6c09cf541b316758462c28f3db253928875bc4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd0336b7ec32aa555dd974e0e3ef66ab6237e86229528c5d0028d5e6ad769a112c85f4e738812b6e97c4de7fd9e7f9e64b3b459bdfbb75a5f707bce0479009ae519dea07d35b235eb2e8a71b31b844e474d3ac70220ee78d6b0f7955ab012d332e9a736583bb53bc21c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f2cfcceb5bf841eae412649d6646a73aadb04bd5e3f32eaaf0b9f8bdbe7634931efdbe8ead33ea03e261ff718acfac04bb08558cec186c8731325de90818a42b42b20308b4540fc1fb919f612cefd75c63820557d63390030b2736c46a328f5a1b9b674d4ae588f3cd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b512349d25364037bee7342a6bff9d2948f8334ed6dd22ac942f37f599962325865dfb2644f2aa7bcf5599cef3f499cc5b1be2c405b2ff4a7098304ef15111e9ec56318a651a0bcf57f095c8b5e06e6e41d63712c37663da078a736f6d2aded5f443cf9b0c9e5933f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha719b259cd85e2a9a6db04e490af67d22d61b69d49576086aed850bc82276f4b0ea595deccaa93d4026a8f8741755bbdbb4c1b345c58d95524422d4acc64007a03e1f04d8f82aaeec9b88263ad358950cc7955f2b8c8f130414cabf6664c0c1138e42676ef2eb67bb0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbe2e04c923d1fc4a98a315cbf592b64b83c566a117eae4f0b0fb240ad0660228603199969e57ea55b760b87b270319eabe853d274755101763072752c46086046e61adbfa0fce2ac21354c90f62b6c28e5a8cbd802e4d3a445ee48133bad98396ab589e1917300c2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h76e4b43ef4e92e500302230db43fe116ca758fa268fb6afcb8c0b21fdacfd3a971ad1f177a3828b155184eaefff0a5af4a5c2f62d9e50c227ba7b58d91633b69cf0aa6b5d349760e7eb4e172f42e91f122a82ca6e3540287c1101f28708d23f4a9ed1381cfe28dc592;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h413c60c61da73d4cea9c7bb3b1c2647654f93b2a69b873ee03513870595299ca506c851a116792d08a81e7684019d2f9aec57fce27e73de486fe4df89178e187c4b088ed0fdf5c39d8ca78662943f980ef35196b5b87eea8fcb20f50abf2d6bf9fabf54c90b6aff2c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he991e45966f4febfbb1700a2ddb690ba9b694e73a54d466948356f7799ab63fd071c9524ea07a96b57b5fe63fc1b3f888cf07f8ae088a2996667c235abd1d19e73fbef7fa00f7c01b4d5701b11b786fe280664feee03dbaeee9a317d15337f4b24b50c2a9a972f1da3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1319832030cb98604ef127f00d247a02c6ce2436ad70f6f1e10161276d01e8b2307574a9f53c01f329801314b9124fa97fa1ae2eafe0ac1d40304323a8de4b3d7d02e07faae16cf50ad79d9b10774d3983e811b9cd7f294b016d0041513f38f9d5aac602d27fd24553a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138a5db8770b489d3dc720cee944942f890c40699f316aadc55b60617d30e13dc4e861c75acd74deffb834a5532672b17ab7b2fecf54a39fdd07029e7bb938c0fffac4bf5ac5cf6c5cd3001af2bd046ccdca393cdb7ea29a8e0f533e6c34dc6dc092f6d729cf45299d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h511fef13cd99d8834a934808a76fe3bf347c0973168d2a11d1bdbca38995c794899df8fa22b7bb6534c4e58b175aa3fc6aa53a74211687953f7effe6b1d59af70716efb230cdf82aaa839d54a8dabd564544b14e70f1f8160a8865bdc826aa9057e6167267945e7d28;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d8ac83faf7925bdce45ae2f967c7176c86c7b1eca82fa4178ad91b1a611b88dbf09c81cc8a59a16db81ecab74ac81dbe6e1e783ff8dfcb746b205fa9a12c8562baad2da1b5c3c93368dcd12e2543f01b7136d12e08f612d0693c456b8b6ad363057b3f145205e5e71;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c4ad153cdddc27600f299b07fba617fd58fbcc41c149a6bfb26effafb559856dd6fe4362d26858158952aba2ceda64e9ad340e0d8641c64ba4606c25a7fe2ffb0b3488a600fc87286a099956d91337e5b8b1f320187c52e44416c3da791e0186036be227da021ec48;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c45752aa508ca38ff8f71b4391f2ffc160f4d5682bf468438b4b13afb73d6b2b3b2b31cac8396c372e5a476d6bcd7aa4f3799e1e1a4aefb412a4276681c7d8c16588ad8df9458275b02a17db4ec114e5eff997981758378f5f3161c8e960f959e834e91d02e65df7cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h41d5479bc1c38bbb6661e59c6bde6f996d6645478b807cf30b53df582e9d790591423f35e6808e7b2c0cb7543b610efd46502e003498cfd32327909a708b3595d938f66f831ede14c6ac222a2cfca014954cd7b62028e23cdff6be196ede6fb75bdfea171a446a57bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13f17c182a0555d92d957bb0ff5e2e2bdae6abcffe8943290157cd2ac341b6bc3757b34a4d0b64806b2a2855f2320fab0bf9ac05ab74905f9b39b278f95bc595181a436507081884d462d9e73bf184426ba4a68e80cf5bf64146716d8a2a3448128e44a629de8ca4c37;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15d88485f28b7267544af10c66eeb61fa4db7c994748736d9c148bb9b182baec3ac58db00f47e4296e7a0007795b319493178d03c69c8984595e40c9f6105716270c7a5c9df95cef3c171d34b8981646f547ffd7d41adde10e20ab1705c66867ae8b8c075dcf2058328;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bc89ae4c722ae051999d0ab4f5ae8964742fc547973208fcff1a5acba4765b6ece88c09e49aed2f02ee7193d21e9b2a268c0503453a7bca5ee3e2dddc65e89faa9e4727d62db0c7df9a12ebf8e7790e677c5fb1c317f85341baffbebd356a1c4ab503a5af4ab98a64;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h58c2ff7ca169790c6e7ac22d38232862e8c944732747f39fdb764c174fc1f209fc802845015d84c3388424a03654f7d3de44611672f5c0a6f5a6ae5e4a8a1fea78f16cd6274d4837b1e2ab75326610ecb453dc863cd2cffdba06073bb28afc986362342dc88203d6ae;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9ed35040fe7b34eda6f6300717f195bfe8f31294ff5e56d321bfa98b1d996b9ac6c919c06d7af24f2f5e5a9d32e94c278c7b59a8a43fe53e4bb36e36ee4be8a087d09fef41d8d3a11a6d7f23687d88fc773347bb0612956ef0bd48f2a1a99c628fdadc7ad68cf8f38f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12636a85bc98ccd48ce232f653889c56fc070a1c7962b1af06a76f94bcfd8c0b39bac90257e2da605572468585e5b1d00d6dd433f59693cf0d1111706fda62f11ca661fd8b239bdf5f3168774b761647a56f3933df3f72bdfc7087691b113bf297756bbd7e9e24e8fe0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h169c8602a02e4e57cb29174a69bc8a9f765f517c1562f9943bfc2eff570fa12fe9356746cdf019182c86552a8ec35b9b751be3890f3e4ef8e38f655b00d9890aebb3f905e5dad7465b2f9b448cc706e2488e45a141453d666b0123ca064c9c62552c8e70486e017318a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2556b42e6bfa5449fc4dc5800bd8f06317fd0eb8caf6202d43da0168210a6c36714c883dff99ab93a4ff4a4014135e1300f6b9531ce3edc66ec2fe91382025f168a7580a42e48f3c120fc0c1bd009ac8895ff535d3927b18651552d113ded92a675fcd4a00b7447225;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h39bbc47fbff0c4f4666869d6ba291fadd5aff478c98fabdcbc2ffacbd3cb5273e0abe26ca643d9fd6d28a9868d615e0dc6a6c1e8c0c132b0ee49ba7e1a866b862aa71f534e0297fddab18d8b47ef3b427715d0ca2329bd0a19598d2e35da6610198ed72d6c5ba206e5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d1fe983d55fb2ae0b44214e197fe1d60df765ea151d79eb3b645bf4d647ed25bfa077f96069d4edd634f682232501619f8ae44b0f08702be3574acfb5e8703bb303856b86af9b3f32cf39dd28b2b64050c0c0941a6bf677d8c694ebcf1763a2fb9ecde81ecfb09cf8f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf725850f2528dea5c849ccd1661ca31383091cb458ed5486a9f6dba82f674c6ee4c05f05553c9e0d0f73021126ca30b1c0189111274f53bc855907d5a0267cd8a66333382a65bef644ce89adbcd0bb9e0692f3df5433fedda6b7347459f0299105504c38974d9e1255;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5bd4723585cf9a0701c80c5d9dd50b79c2d9fe6c708d292a56f68defa2f8fda01f69b74b004688200de4ab5760f77e6c837dfa42d6755fc6375a1576b3eaafe2bed594b843af4782b4618c3c06ee25cb72faeca71e29bfef2a42c9b2b1abd7233c98ff6b48d05ba166;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf7b6d3a3870d3e50e382982fa2159aee7036719242637607596b1113bd27e2a443b18e34cde321d6e860b41da914e8eef11c504691d4c97c7696d7cacf667db92ee8b7d5739b90286a967d28939389f61b139f5c9be546d989039427431cdd3d9e1909c0328df7cbc9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3486e246f6abd2331b5213bd66e710f4213ced840c8f6fc7f0df5cb70be555b42f9321462819434fafe2fa8b17a47decb26c58706b47ed0d2915b17489fe84984dbd91539d62630420a0857354bb399277455a8aa979e0dd3547636342bf6152636f6a9f1798305975;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h124ca8d7ddd44684cc748a12f01c312542805b686bb27c54b896d3a9df844073c671740156b140c5da0dc208ddc8bf9ef92c7b93e93117b374f95a6dcb0440e452dff50df7045784e3540cbe79a937de5c9dae72ff78af87c46253caefde03851727167b90756436488;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hba0869f7100d24a5e8b544fda74c777bc0ccddb359dae771d73e2362c5d80d62d5d998ea9d2dc37149c8ffa9f58dba0596da5b6a7928f94bb3db173b6b0ab94f620189c237c2ae32d4d33dd7bd2159155bd423dede35dfb94cda195a2ce40555b68752e433effa9307;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5f0d01244f949be425e5b608f4ac798b3eebec55f1d402f4595aeb1ca82567bd1587a04a0a4c5e10447619efaeb712fe3b2f6ac46069c0b87e65dc90b9c017eb6f4ff86bc241f4d22d11640ab3b1171424c614462445984ef1d5bcced5e6a47bca0d4932cdb952dd19;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9764739e5e63526343cd21847948e54edac2107707bd6d755857948f481cb5c4f373b4efd4baa7d3b842cf41f66a30ec3d11518b6cfc9f7a3658fb665b73e3b1dc9b5072c8367c692fea94284fe44a2442b6455f0c56e7d6d29868b753f76f4f0ddce45699beae99e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h53a415338dc2c5ffc6a36b9aeec54207dc674a7729ad2143cc9774e2db8220b1d3b286625476896116d446c4d9c3ca05bd3ebdde823e1317d7fa0fb015bb1bdbc3bc4f2ab33b2aff2725a05f8329d857088d664a073fe8ae9d689801d9ba5feb754d20ebf9bf245fe5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6a0c5f731d38a1f399777591762baf14d84fd08a5fd0f4268ca6f714ceae52c22f9573470a3d35faf1d4dc521d620282c156d8f4fa6b18001724f79810e641741c8c2b142251dbb547993fc2736ac355e8b8adfeffcb250c4a8ccc51d6fa4f345afc511e88740d4acf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9452512bf3ceb8020333be42347ef796555c3389d829732c55aa83928b75c71d0fb936099b7f63a72b08ce3518848b93b0116995e13ab5c69f16f14d128a80c7ddd367df9b586b86932dd628c248b918b96b0769a0c787aaad2efc513f3f9ab4f903a2ba22db091b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1faacbbe3c8bcae8291a7b83a33ab69dc76564387ac745bddf9a54f08e548d6aed20e97211e2b88e68200533672dd62717aaf7997cea4e8a77d5df08c7c1817d507798e71fbec98b8522a5c1d43d7ecc09d9cc3fbbc7a646ab7b6e6d3d88cd28bedb1390902e5daa049;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13a53b11f8b82d96a5a10f20cdb99e6c8425a0192b1f38120703c940e0747e48ee3bae4358cc8b235484cb2f7859184e8c88fded7c6d10f54abf0e08eb113d53b3c91a1282b28d6b9ff2528ae6d7f349cea7511cbf01483a34c7d45daf9348f255423491b23bdf2aa91;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3e1fb40eab803adfc6fb709c25e2eb140dcc0e48c37460fe562c86b029e3b11f1fad5c16dde65dde3e2e674a47ae01f78c2dbb55bf51371d8431fa1aadfd9725022425160219a04b7b04684b7206b0ec08d55e62fe7281349234d02d3333f12c6edddaa55fd010ae9f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9de3c9a67949617181db7c87888bd5456f803f364652c075c3faa380f147f8fcd62cb13b07b09cec55dbaa3661a64c2dd7395cbd2e4b4b379229f2210a1fc73a7ebfa12aa6d8a5f103200fea8ab21106e41cf7200cbf4ef0104ff636f0032bdd8860c2ac3193a945e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16bb39d99a78299c4dcd2d51c2ed255801d55b586821c5a1ef15c57989b7ca19c2eb58c451d6c8e7bd24c8316f31a3f24d9e1a0e9b31a9517ce4ec56b09d9a0f77b6867a9a0371e7c0a6df4c184d4518bf111708d98dd65e76bc71a58066f96f2360589aad6810fc2ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161a181c75c32afb7a070d328f4dd16977f778bca4808e8e0d3c905c3250ccc30405c14a3139241c15e6990610b5bae9463718113d9154d1f5472e526c9fbc4b610e58134fdfb03201b359110b01cfceaa1e911ffb0d489e6dedb07aefbdfaeb4d531952d156ec0add3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4dc9165d035aac7da2b4d9a2605eecb4e8204ba144d8bc5be88f58b098efd3a46db769c83f6e23993716aa7740928cf33401573c2f224622dedce5a95c8fe79776cfa9131dcb58fd5b13c44c62e8bd9abf372014280dc466ec780947766e32f36f5dec4dfb2c375005;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c8a2b815ec706050d379b9f27a8909605c2ab9ea15da999e5792eaf66ea9c43f382239e15dfaca820c818b92f518b6599170a41e11714e0d828d14972dfe0521a30921f73b3e824f55f21717f754d5a2c319995d59ecc9068bb91c624f8f788765ca0255e255f7618;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2a94405bca112bd8c80031666265ffa062a11b68dc12e2a96e97ac1957f20f9313746d52eae52c84b0c2813e86900cc80d08bc0bd226e7c271aaecf90a3a703f23d0a24cabbd40673def5f8303ebebff48c546e9a17810e2472a1c087d7c3cfdeb6c40dabb79b32ff4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h126d9dd9d2c7376ef5eb5d6ea86402077d2b0ec6038bd923445ced0a8a3601178ccd1548ce60bbb468162578b1ccba66e1e2d49bae6e30c78b2b1d92941ad6a1e0556b6495e621700b391b5ca147561977812ff289f7853e9a21841300fac588599f224d162be1af74a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h429df132f0c2e21538fc1ff50bec8578c925b94e3c92304c358cd3eccd66f28c6ac5ee13a5c387495534e9e30f6e0fb19083dfe04123604a6539186dd863e915bc197d99993225e1efee5d2e4ebad00c201faeb83768e819608cec3906b9ce7fc410df6620ac912e0b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7e2393afdb7ec3eef28576e8fbc497c71431b3d869e2d47b2656c32e2fda17d7c21abb97a7e38988fef7c63cc8d7a6d9feb19bf0da10f41996509278350ab08ee06e68a7943abae701a8e34272c1711098a85cb0e84a76cc2dd821dac5dfb2f375bc1f4b10be4bc501;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b617b335a2963b0f2533b1286c1f12d21b98cb6b2e8c9eac982a80da0810704399f7c9e3e66b7eccdf94601e14c86df8e0cc4669f114726513fb8bf4290784e17800ed425ebeefea7b2a67b548d33d1be3a2c0a9b6545df8ac5f71540ce4cf5cb8e59f2ef4f8ecae64;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha0d2a9d466995dabe55cbdbff51f26508b9f7f24c0ec4db96a782b14e3a85012f5c080c5fea68eeb095eac8ec8ed2ecebb29823ef3ad99c8a5eb01daa4140eb3558f019a0040ffa76d4993c5d17b08211c8a40586cdebd27176b7d07d33474d2dad1524705dceff738;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12d0562bfd83ecf96d8ae8839966b057632473b4daf7de329f3e5cb5cb661847ebff317cb026916b31066654a2d377d97ae0d5e1ed23da144fbb83b80ad84dec34846ac7af5628d26c72dc7a3cc775f2b9e07759f229cf9e57429278d7af09e7c207a5b1febbeb24fa4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb898de6e117db2fd961a915fbd407c558ee14c6171302970a675caaed601498a1d8b769622d531d3b9fa7be3e77ef2a0944de7558803c79170b52355d579f3391b81fb3dd793da1c9a84fe9f4278a03cec99fbe372ad8d89fa5c39fb9efe1594ef4d825b511bdc7c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14172ec62e28e1c2d56c28e7d3a1ca1495ec1052dcf2196eac8b8e09b7f3eef7f49ec0e0d7850e2b15bc533ab32ac60970eb41f6067e13f66869d8acd759878ffc87038f748d9cada910ca0efab559edad6fb25c355acbdecb1bab99ac8369aa7ba78bf1449fe683ece;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h220f2a66b74ab0dc7b7b026d34cacf87e46169dd0211303d8f73f15758fc60c49527ade01c4692eff383310c5934f0350c36a7977b7579bf0fb8c7aee7d2b4ea913e5f4ee5f918d2df2885ce0ac843d61f9ce42ec5671c6318d75b5da45c2ea8190197b657e9f108a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he75d32e783819319b52113fec729efe3dea4301fead9be86907ce1d8202ec3839e44901167123023f575f604066a825f5b602583e4d5576b5b6729a373df989df156277354f35e88faa7dcc026f01f494f85052a6177963b41e5d628cb4869c2b1df849fda607e92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b29eaf914bf7bec804ef90212300f02a1fce8e41d420d412e4adb71e789d8a3f3da7af096117690015f766886f299e53d20b62d4830b69b9a998d3518cc93d39ad309bafef49cd66f3b4563deca02fe2f39a61583f3e7d3822a26af6a350785cf3ce9f031d43d10acb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h497f6ba38329e92304340ffedb15ad77267ba647d652445aeeb4f6c2f1a8ddbdf584729389e5c03c794abb82b166bab8d97523a083917ec07b79a809e5fac49f741cc5894aef6e6ffe2f21f3fb97693247693990440f94b4f73294cc99656e49a0ed8d6e3966433963;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1380264555019f36ef7e87cfaec268def60986d1a683c1029ddc26e1c759c7ae39f5787ec1fe36d52421c83c9359b007b29c0b6e414073ffe7c4d3531cace6af0842a1a67d83db4b1042cf401d2284ccd484046f3773da508b023b8cdd17f43038b3ff0bde0469313a9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3eb43e9eca368949dd6bc2720b67800b8861b5ee8dbb24d82d6f293fd356d54bf2091b94730bda9aa3c0ccb254f27f2b973ec1a8062fff542a58ebebf5f9626cfa8982e146bacedb4f8d9677cdce65b90b15f194a2c9ac843ed3688f39189d3f6334a3a54b79bc9225;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1451e18434ced25859753c15beb6746b679e3fa8bdd1522b36c73e32ea2c2e38870a9b7527a3023200b3b3dedcbfcd72280797cbb33a516e7d5bed3a98f7d5efaaf793aa34be4e3f89997d015ddb3578692a770aebcf7519757a81d8bd9160c23c24745936ff0664df2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he621d6f3bf2d85485dee2b71dc643fc4683076b8f148153c36d142bd8dcc55b6da48cd54d243ea7ac3a5c392016259e9025e209e4a3a9379e81f16eea2ab3060e0cc702ce1e52c47b4f26f07188371f04b82cfd5b73450c2f8cd5e663a1ec756f92bc1323de6f4d7e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h174a01468554cfbd29ae34751c77dd142b296bb466207750b3125c3d0dca2e0fb0432c5fa8abf0ede51d25a65b22230dc42ed7a934adadf7758ed0919d4a947d792709ad9be63ac136441202bdd27ff9fb7786c9ad7130b100f6e898208530254a279f6efd9b2e6327d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4bc5cacbc6eb9a04f010e1b13db16a2e484e598e93cf1b6273fd894b8b313798363b9f9e73e1ff19bca5893b6eaed010e20c304e4901011000a79795a89c2202c21f7000ccba51da56d239c79e19b91c625947b0936fc46ef6bd880d6d303d44432adf3ebd72cb936f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13fb2043d2a5a0a8ab7b07e2554f52cd53b412171421d35dce8b7c4bb461e67b377df994dcbe5fd8c7fd08ede2a76731c459b13f9a76143c9d891ec65ff0489bd2a14435d12db438b3d3ab6df35a8bba44fab435d8f2168a32e5f49d7f535f3085024573400365a94ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hab42e89a98b5df9c162b6ed3062f0feadee88a65b621e6c7b9b07ba2a9b803b9cbfb7772a510e8af5fd2ec6a11d489c1de449d8913d3483fdf5cd37e55ac278b9ba0041e2f7a734ac2844c55a34619f66846a43fd0ccc4e7fa84e0124785667543754c1fb5f2cc7397;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18263d77ee0dcc45871ba67d46470d625f264bf0286c30ff09f039e30a83fddac18ccfce1d22b474bf68fe75a591fbc3ceacd77b002226ef6c3ba8674766532ef7ef0d9690a29753b195cb660956c976763cfd06416d809cf580f73d25588beddb7a60a3c64ebb6141a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eef38dd48a98df3779455f7b3a14fc54437c9a0b86818cd16b677b7d9ca7546dc5ddde58d4c1af4c5e257586bafbb19f2a61c7547a5e62cfc7e4e8820cb60c2b6b6853e1fadb29ece3a3f71020ce621d3a0254ecac1bfc9cea319907e61877ac9eafa2849d7aa626a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1505abcc119f1de5c570e9f8867579d1625a8e8f1eddb3e34e509533c18e15d200d899cf732e11b94c72527b73dd4ed604cb1f29256c5ad4baef9b910ca6d7f703c1beb62e261d10333fd2afb8dfbaa647e518ce05120fa68d570188394b435814225624527c1df8ee1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17b85b256ab2eea7d478406b21a84b1d48974d8a4e241793bfa62d0e1ea8e848d6d978fab326789ffd1ab7ba7c18ef3b5a82ad37b442510a2f71625f809ec5a260c0e5d99993b7a220f1bdccc376a6999d5f04cbfedfb030dd0601b84a98d6231ad5963e2c3135f346;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb51da864caad37f53dac72941be074ad7c745d388a09efec26dd568f529b4e33af70a058e8e0ef97eb6acdb88530ea73e8810395df44f6d030c63531ce1ac9a99bce1e697ce3d99250a70fe0d245a1ef7ce1fd0af5353a237a78e16ea23159c26d836eddc073757f3b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ef5f240b64b3abdd0cae05e449fb59e72a968223c44553ea71f7e2f8bdde75f9d42b532ca22ace25493c7fa415d50726c6c93184cc93b7fe0b3efba7e12740bcc4f712ca8c32c1505a2faffbc8988c83df66c2c0a935ecd34fed8b705ea77fd61454666f14032c3d4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb76d0a5e31acbbde952389511abf79c20d82713469c4b4a4fd1264b54c7746994afd5ea450ff5b2eb9867d8c15af68b17ce96a7e98e47458f9ca3bbe99bcfcb8553fe74e0a6020f84a1f50d0293b92f00fce11918ad21501ebc588f0a29624f3db0133a9bd7fc651be;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha1431193042ddaf8ad134820b97e5388b6e6b41df27a3989609b9eae1ab42ecd585d010864ed70755a470adf3819fcd1c42d749902d7294d2404b484e26dc00323dc3d8aba89f42b937e59e3da446c57718590045e7d4a54a47b99648f3f9cf636aef113bdae036141;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11296a4b0a61ce0040a0da7f6f34d305da37d1973a1d5616c790c9b180c33392fd11ee3015831a66300e8e661ed1321fbfea0d265a8311e8b1d2752afcf77c613c19ad81bf1dc5353b9f90f5078eb088d1a6d3ebf953ce411d9f36327dfc702c38fec1a4eefb3da329f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h111fb14111d6e58db4a72e0fb2cfb9c6212dba1dc3d248ee300baac9da060d270ce82c16d5dae452549aadfb85a5bd84b0e1297b2f9a8cea34499f1c19595189d70dc3b03fd34a4769743ceb75d95ce51d787cfb04488130522d7e72324ac5629e9fa073f592faf0fcd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8e021be6af31a7e2ad10a6eb5317b1ade5d38b6f2560bcdc79b2dc453eb0107c5572b242e9940bc6d812aca74a602c52b88371629ce7c00af609a6348b14d93b1522dac8f47972e80da79ba6fb031ee21bc262dd7079cf51ae2c4e6c8b8c05d94b45119a9fbb8dd438;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8add852869fe5a3f294a74851a9e6074ad0c4ff18d5be076c19ea3e67a0b6da5b32acebcf24ef3cba460aab2a561ea6851e82925a7807f226f503438b3357cba59f9793f0b77dd94c60cc874289ab6cceb2c0a529015e8895808fd2cf86f852440251f29d75d6e14cc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b55e98faa66365b55de0d50b4e682de1c357f544be56b70518efcd528531cbbedc253cd9ed71b5597ec49f61b2997566e8d3e10b134367a158aeba26ca86703af00a379682a290c0d7bce1dd7a3dae091da964471da2eb2b7c47910e2929163a9e69ad9d139cc1fafa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h122f20020eb5e074fa54569b0d2c873e523baeac613e387f0d509dd8b10aedfd75b205cf5aa4618cfd7645b6dcd8f08c5c70b18ad60dfe0ffc21b62b59af0a7eb3676776e3d631f8484b48302e3f73443075e6be5a3f6512f58fe0630d3c0919fb9e5dabd0a677f5e2c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbbb1cfabf81b626125270f39113d449c3944c787000c5376aff29ac1f1c514d1ff60396ca853eb78efabc1037e578ed22da8f6e0bd8d683bd7e5fe89bd1c1d452df1009c8b1cda01ddbc2537b4c370b6799ec1b679f874323d5117c64beed3d8952eaad2ad0f6ee94;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hefc455809405b3f1841f120397659250171a95c14e0e572ebcc038ac008648e66acb9022e430c6884ea3b521a0e7108ae010a4862ca56bf1799745feabada6bacc16f3c28a81fe549fa2b55f701faa91350c9b3b065baebe7eff64f513b2f04546f90093af9f4bf98e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h420094e79d75f9f7459da1597a8c9a1a25a7aa47a46dee2acaf844d3452acae86bb454d616a9b7311c1e489a56420e19f63cb308b72a482dd30fafd550bdc04dc84752625903ed496e366260350706e035b13477d48ba3c4ec6267e31104ff8a40086a7e653678d07e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f835f092044cf3a06a1db6c81f8f7ac54bcbd1c28a154e1a59300c3b1df093165bbe74ba54d59c6f2983ded2b2a57a775376b87851f9878ce992564416be1266a4a867832e3f11490e6c670b8606bf73795903bdd0ac24e213c4fbf4ea91f3c1be6556d8eebca98aa1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he32aab7b203e03dd16ddc9bf0238736a7620efcd15f4e1bd87dd7787a173ee4046ef67132627d2605b75d0355a96a35a2f3bad68ff71cea626a869f8226725c5687b89bf94b06d121430565cf0813bc1c4627a4c75685aa5ca84124eb9f0a0b60068ab83c29ad73b56;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18956d9ea7c1caf56afbe760909bf16edd333264cf4349ae6e9147b73d1cac1ca8aacf24bfbe2692551e38420b41329ac02e3a8120628830c8f52a3e77b2c12dc6766ce74086e231cf354586d05397627b079c38ba79007f2ef1d4b3e50b0ef6999609bec5661c940fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h181de320182eded2d4badf8bea816f31cca6f0c8d3cbfc0d7342351fe04a0d5000e943ef438dd3adc412dd4cbcd9c97876184c474ac7615b1044c772dbcf57345d7f4e0fde445648e2077efb7f8876ba04b3d974f4c258a90a7c233b7c0008f0d9ea13f84f8930ad16;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7ad8ae1e05f2098519b107192e72a9f1d9eeaec1ee1e80555a55b2bf0fd2271ffeaba5d401f1d6f4306f2c7154b9c161ac5eeffb9b79ec2dbd6418eb7a0257275b17672285a509013e0b896ac2a52a0cffe41d89362ccde70b52e08915c7fc1d8d2c6f86b90899939a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf0c8c522041edc94a0dd1896760c3053ba0477aa0e0cf3549d32cad172400c8c3acbd46057e0d16d4b72f9004a06ead2a5ac0238be7c1ea02689bd626863fd4dfa385f56914de903028d875e7bcba2a756d02b4dee403fab10a807b14f372890e40abe595e0f91ea93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbca203852497433cf0a47bf8e342e158cf11bf9929436e1f2ae39e691083e8a5a5f0bf51d0ac78638eb5ac01fc57e32014e4dc78d1c941f1095c23e300fd5a9dd05ced9a8fe91d4167e4ee170046da47fa7795c783534695f92077e28cf235133bcca1ca62bdae163c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12c5df0e929f5972c8a6b9f06f2fe8601cf0dc57135f2e92ecde58c39bb0af42f8fd4cccdb791c61b8afb7673678340e1ba9bf296d5ee3c6fc1b9cb3a400ab336d0b91758a204c12f75f1456a96c241f21d82c8fe4a388a4c0b3f9033e97fb6863ad9c888019cee1cbf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h165463711f6229de13ceb3f0a20a2680514368fea00406be260a326fed9ea8908c4421df5eeb0fbe27bc2fb7e7eb54a849bb6e98dc26dcf1e6e9c03ac7263d82bac6aa350a0e903cbdc51e5754343f71f6197957a890f2a4d9b79f3aa80ffa4ece3ad58ab743faf55d6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfaa859968ebfccc1073694d7673c6f7744ec9b7e59b5615a4c767571b0952f7216cee5edd689602e895503ab3ee24ed5315897d3daf2fc7ea83434e71ab3edf2a1625fc45c560f14889117c8dc6adfbffb43a1fef97cd064dd5f10990cc22cdfdf3e0e993f50d0bf4f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdd8bc684cf5fd47fe4422a0cb58fe764c324df43d6b4ad0410f0b8c0162f49042de15d0f6ca8f1f6f638f85d5efb6c5b656d102fd9368b7233d3d7c975d393eb354867b93118737a4db6b46acda2c3a63f1f2396b365365aa43806658e7521719fdedc5b38440f57c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c347370659557dd1d936536c610cc440681b706b5d48c1dc6c566ccbc1cb550741b5a63f21ad7e0c8f9666706d28285149c94fd095e8f28182e27eab313b7c5c7ad0d9053aea0b781fa7222e03ea1bbc111cfbb71c16938651cf56b73cd38eb3a19b6f663e3a73553c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5204bfe03edd7d9ad347b73b7b1cc80fb2b59aa96a3ff215b0e04f343f7c1bf827dd7fb96d1010b0fe7e3409e41428e7fbe9fadf579a735f68bbd5f31b5c786e722005a3008e5797d84ea7c6cee9d78cb4bb4875ea352f7a898571dd7b9ee6ea25dd380dbfc92e4bf9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15ee5c4a6f27a97da565e4eca995e0a6d9e468b5d16c5b58bf8151c00314cbbac317e2a297c4c1ba80e2ac56896fe5b01fdb22152ab3d2e4951f3361ced6b7b4e46c60d0256ca8f6efa0524573e84d318e4baaa80ef9b76fefbc575d7bdee6bbb2f2bb46ac06e0cc996;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1678b075544ce394bc11c146e11e0b857c4af8a0cf924102dc99e61466708f6c5abb66ab65e903002ed4b57943ab9fee4fa5176256dcaca26db14d111d0650d353a22855a5fe9b54fc84df74d5ffc7876c0e84aa8d575606d5a8e2e20a7976857510cec5ac251428039;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1813ea5eb405859901651af270a3eb981ae21019a52e2470d4b4c80d91cba13d8ccd05a1cb0a31e392536fb7615bcff4dee35f00a42c3b764ea93d28acaa5b0dde1b7ddf95741193d20ed956a18d47ebf491b33f60d0ce95d68d269c9602afd68e6af4243db126c13da;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f0b8faf1f8236421caa5079e7c263b7f00ae6b75fc09eff2d65c718f51441239d868a0f341413ae5303ee1c43f21b740db1a56076082c349789fbca2bef7c8c9b494209bd31271340a5e283396dde8550d263f347eb263d09277a4da683f8beede8cd9ba2a61235e89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h15501f2fcd15082eea4dce385f1d4240d28f17d900c36af9d26fa46f2455aca2f689ea0f0b377040be132b1dbb58653f55047055ff61c74a43c914d56b56f830ec96c6c3d3c70c6c9259e9c97193643b62dda4bf349b7f5686bc8693f873f20c653799d11ee07e8a83d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h117bf8c9102023dfc7dba174f92f16568a5e5eb6b0a752af58ea63ccc1373c6fd36336a8a9bbd97007a1d78088e60acb4024a47f5fd4cde19fa3886022ad5689e1f1a56c721a632074e46975239a8f2fea582235fe0ac57ff8849f7cd3cd11c4a6f53bbe8e56f9822cf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f56e5c176a3c847a279872bf785663c03b15b38cbe9c1790ade8f449ac470645069a9496d2710555b92eaad681cf6937939d7a7d7f8e2e6ae4a8f78f687454fdf06455ef48e0e989d7cf9df4886c61b9745f27d4ffff6e67f80aa3fc07f77d536b0db96077d8a0aab;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ddfd56e9486f9cfa458c98534fd88f141e3f75e80dc3bd004d193f723b16d28ce9b2ac03464cd28dbcaa03eb949e9b135afa68189b9c13b53fe711f527d2f52783644ea9d49604136411f01c8451e2d62bc3f4352786d5497e866a801d7e1c29e3df2d83250702baef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h132176cb1e8d5a537ec46d7f8fe1a542fcbb7b14dfed0e5257115f9ee1c27116c7bce654ee69403032d38fa12db87edb98a0e81303f49e16d32b11efb138c1c83b92bc43ba3f307fabd3c2999cd83a78bba60c6b75fcc8a39d4f6ccdc923c124eb3b217c3fbe1688c86;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9110aa51986038f338d10863ac92dbe2b7321a8c91ea15a9ed8dec4f21b7f10c7496ac317d5355e5ed22d97064a881afd45346732bf40abf0f7058618d61eb785ea0a56901751853484fc5580023b9b512910fb03d5a998a36eaded85a4b5936f00069e153199eaf95;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h138261aca71d2ad2bab657beefae9cbd72d72928fa4a4aaf971cddaea61b7de23eaba6fe2eda09a4a6e87c4d5291af153f44cab1a2c3d69efad03caa290a837e7fc26c0d8bb8c9bea9b59e2f15a8637a96c3430603a4ca1378ee5396a62ab9d62abc504759cc5b28649;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6b4c49e08c944a44128b992091e059308921c431c5c386a215906edc59bc717e51485db254ef659562829f98d63383d473ee4c3605deb48b0d2dcbf8d0d5bd93193fd74c3307fa01363f027aaf3b8102f9f038413cef29b514d699437a8edc1dd5f95e959a76921762;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3e7dddc74bf6ad7d5a4058af086b09fe8099b4081daf2a92ef0ca3e167c294b9c0baa6c3678381e0051fc2a0de1387fd1f1ab3618492b3321bd8a2d8735d62eebf48f2eaba9ccdf2c6cb22d5e1733dde5c756b35868765ff208c9ba193b807f31d51c84ed4f5ef4f1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6880df422690a719eac06820ea694416273242f20e4a7c8e3bbb8144174191d0056b6f9b0f265dd6b37efbe7664cc2bfd54c6aa8ebf650114903b0e86f0d80ea8855a2113cbe510587b958f23608390ec872079b8ab8de2eb389e1b2f29629d462f47bdb7a5fe0ab6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1949e994a3b8ade72e868bc61031aa92c3b988a05290331bdab93cecca601dac8c2c9070f48e81336e224d025c3dfe013518a40d32b5fe510d45ae0f225d2ab073519d4a200d5d52a8110426056c43990c08f4c3a7bc6209862995616d62de8fea7a8ddff64f09af2c4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hed7b825f8cdfd0f3170e41ae88279e74686dd7d6a914d82b34e2774a7ce56e6abc529915f46abc74f0cc3c891cc9db389e78e6cd0e86eeb6280b1673cb5f6037cf7c40ae5a3dbf4b1e0095be227ded04b1131018cd03d0b21641c68c8cfea4096492ce5bf033842201;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h160a2905ba5cc5e507b45a57a2e9527b65eb19a1eca5d5b772af70013242f0fdc0925f2441a2d4304195dc7b1a6ce76fc3602cd087629f728aa8b58856148b2d780f56978d68620c7c5a158dbfeb1f74546969df2ae3d2f1609c9004c5676bda815d7ebebf136a3441d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h687d60c972794480f080f03626c4a549c2383a36d360ad80ebbf1c85c701f767f97efcf174e20ecf61efe57c14b278b94e0b788d475b6fdbe2d18a2b4b5761a567a489cc3fc4e86d747955b70778c02216222c9ae039106a73cac55c0740e4a582b134ab446aa96b5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h193d3b89c8c117d5709b0573643fde0fefbccaf5ddaf5d56451976bacea5a22f3835665b5f97c3fceb101a312ea5760e65058ec3bef19f3918d15276bc13b08ecb7bebe38e37676d62619ee4fcc87e708e18142d668f129a39b749d23a3a2ec00b7d702a4d8e8288446;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d3d300eafb79e794c520287e7c5901adbedacf26534ba68fc69551866f6d7e87868f8464be31b547c65e7771e4e3907670126a656e9dbb8859a38d9a7ea35ef012133a0e944ec2642dbc443cf1a7f53861a884680096ba8b5f0babcaaa590da0e8935fd7e7e66a9c6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1497b45560b22060ff7f9d388dd6a482001bcd70074809ac4b11a6708ed9902a43d2b0086db4e62c3da7e2fedf50b06e13a5244b6151594e57658f3a199caba6b222a60a1eac82b67a2007343c54d8d32b778be54b3a4631cc3caa19cd845a2ab8941e12bf3e9b360b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190d893fb1d56a70ef7edf23a1aa0c5727e6b404a0d856dcba9bc49f1c6997c22a0357d214582cfead0716e59a18ba858ab334ea9d37b299872b2fc7ae7773f4f11ab55fd87c40e57ac3594072dcc55bc757b21883341f439cebd53591343dc77f335517388ba09d50b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd775c93cdcec806dd52069cb5db03c8e0a17151197d97e1f797418793153b2edab139e1c31ec9f53e2ccc78bc12a2b0c28333f4ae13e2cec77665a9eaba5365e9d5f72177b3d2c786dd8ef251ff6d4e213eff68f9e0c10ae2ced667664b7ba2129276e7ca12df63cca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h155024e8cf759c0f32dbf6d5210831028e5bd7009669414368b9977af0691cbcee3d1813b3cb901e055d552d4962726b1c9582523b9bf6ba3bb6d2dc140e9a4c083aa6fd9ad29e5074cc69e72f20fc1d4501e04c0a4068b29ede4661e3c09e975fc7c693be0b103632;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dafe3796b6951e571fdfed4913ee947e61d15d856adb5d005e1290cbcaa894a11a458753db38a5546da7e74075b35589f63c5e5174850881857a43b15bef5e2586864753c192f16a55f0a04bf1d65eeccbe335b00e1a7d7c0b707b95c7e62db27f5f71392ebfb40cef;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8bc1531e71813e1d7c7027ac17648479f86d7602445df66685ef083f104121c9c338ffdb99dd82c8ec8f2fecd97385737ee187c9936982cb0a567a838b8a8bee4496a81fc8cd5f6697f8769d2522e149cac56247916a8961a5318e45d8db6728d7e4ba93d0fa41ae22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11f172591e7f394d08549dfb72cf374ac617b2a1d63eca39ef5f82c9d047cfe0ef49ebc81c0b93ef2115786bc92f342abad0ce076f8128344119a21cc5364716e3a0c5e1de2a5a1e4c1ed5c1a1bb14b8a1501af60b1cc9a0d0a2d4afee2a99ab71d4063b8494ec1488e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4f755775401cb8af66c98eed61acdc84930086dbf8a2a4f17e14054895c3e91e2572cb9d86d7615998bb84376ff4dc9754b303a5831c25616af08b6acddea484d6588c449b2d7df7f649d395214dac4125093cf60578987ba60487df79e3887b9132452d848f2df7e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h69317a5267afd3cfa18823ff0172c1339f096296a62fa884acf2754171a3910ba75dc1e2fc89ccd7efa2b74e1523493a09e544b650a3adf1e1ee007a1e54eba70d9aea796ccb0062cf7ae2898a6509900ab9b8a9ac8c19239ba7381b96cfd06d9ae193047bdb2cf85b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12e7542169c7c564d1eda5f5ca4bea4de893b650b3e55d4d882b5e21c8e0d433983c99210437a7afde7f5ef11ac1614ec3f2b6c1a0c7d322273e61b8d60d0add9d3bc69fae55732861c8959ffb7171e01a92931bfbc9b1c4730664c8ee1d06eed6a5e4e4ffc3eb16d7c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d667c957ec858dcc3e54d39f50519312c21474245030ea56553f750ebe382293d9ac1def5a4d5916f211dc3fefd9b9fc2138df78a45a81aef099434fef3c742e6bc03ff02fed63998c2e67d72497992ec3b72022b7952806c558b5d5cf663409dd53e6fd3e28c5ed2f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'had3cb49e0db6a241e1c6ed43a316b998fe71cdf16fb3fd9b3df25793f13a0282241ea9455224f844d9a8a96444c67345acd3f5ee5d859dc4f0ae9f79a06d2c2c878b1bb7190dbe4038177eae2d5ec889b8bb75f9cc431cb3760fcdb73080a17d241f2e2bddd299eca7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h140656bca38e114879a97231c433f7de00fe765aa295ba41fc911db6bf64017bda245ac3da6f03ad23d58cf56b4d8806cc380c45cce5a2a5a27e88e4130e91e17d8be727bdf6b9c69376b0b6824fbe8f65fe342b19a9ccb25240834fe25737f65d94ad80859e565a0a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha31b1bb2a544d662180445b82bac9f2e014d36d3aff1a2d51d78b738d356e1e0b68cb64e22e65fd44141d3a83e1bddcb72ec82022226a871d7e55d0c5886920195b6c8d0d3860cfa510091a7f1273c5f1effdd57f3f44a3baa59ba2e966499356eb844da0740476e89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4d6233e873f155ae21f598b939dcb25f70e674c8d6c11b32d862073d55648f05cd880058c577c40b413861117db7f81f6a52e6ec57742421b4f96a3cbaafc2d43f1258c304b20d2c89ba29383e6f2b4a7b617df44f92bf17e55c214b649555206246a8fbe385804c78;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5a8912c40b495dda004a7b12daca5daf1a192ab4bd8f102c04e5457d00db12f72c2cc9b56c1a75c118cd415fd723e2077dab73a14ed904a9154562a444157db09ddd763a28d0b0337740a50e9c9b28f8fec272eacd23dcf8d68f8c0bb63adeae5fcccb08b9f9664567;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc89341e8bb45d2a5339bf2c326134f4ce92b1bb0dfc98c7ef6ba8c4002d35322df2d1ed4bbf2429d8a02dab0e3e2477cc564b92d63babaa82130d9befd3fc7af75db118e5f78ffcc95fb4bea40b62505a04ce5d82bc6920feafa5d5e1b373b7641cd98d3ae4c43bd61;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fcbf88b7ff2cf1aac0c3bea577caa3c9156e7c7f6462419980f9b5f4796350f0303a9097fb865ff21d3708f798da7868a22e7f9225654c8bd0864135c0a5241021a8321e22aa27329d9fdda796f06c162d389535bee6528589c2ff9783d27a74020ecd724f257b554b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1efff789ddbf9594499e085667589a859cb6b5dbfa691b39388240d2c417a404517dbcb6efa987e831f7383be8283f8d41d205414675fbf4baf8e7d4c5d24b07ea3c4bde81c390bfcdb5328f0e76b5fc1572a9aeeec14b32e892514492ba2e9d6fdc56320f4d2178bdb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13ac4abf84142755c17d693fe28f3e3e96b5fe498c21e4ea1e67b30036dcce44f95d099faf9f44c0cd731d090e8a005ba5307703d449fe29db99c6f9993bc895d8a037214e4f7b101471e8d0491d158abc4f9054f411d4701cda6c926d5697d454a7378e514d7421ea0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf2940a59e13b0f8693950e371ce4b1301f24aecd1456fb7daef20a3ba58f33f61279ba020d52f928f55a96cfcecf60118e2d41426bbe7b95bf9c5e6a58bbd7edd996d3626818108813666e0bf44dc951733a95c37895aed797aa9b324a274a3db93d1ac9762129a6a7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h79eede387342b06154f216d511483901470b860488c8da54ce3ed655ee367514b4bcb371f1564f220c6c9294c4b791948b4c5347100df145a95f27945e0d927decb712035e4ee6f29ec1edce52825a6158588c1980f160bd1fc1c71cdf646e3c2a56551cb127eaf7d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1186e93672e06912ede0ad16dc2b281f78f9314946bd7fe78d84173e1558cc0eef3e9c04c35f1d1089b22663215864e6f37351b7baaa147665cc0a2f679b57ff0192b395d0f3f7a877e61fa6383262f0487ad477d5348ddf4e6c99731d34d053323cefee0cff0b51e7d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1424501f752f338cfc00bae4a821370af99f30c050617aafb300da33294b499ddde40c37f0426e9f5d9ed99e22101a00d758d0c9c30641ca95f9a2955d2e86478c92e0dea334ae398fd6aca55aaaf2966fb349109b191abdd2a78a01b329e716e490ff23ad4da40374;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h9296b6393b7edc08315486d89f9e4f5a718a074296487d320fe2589ffb246e15e7b630f80b955a0cb22140fc45bcf25917838feff005f00c6d5b4fb2816d1f1c3084200fa2c97c00bd16ed5121e58b0e639a210c429b90caa4f7a9e18a4062a4fa49288c992cf18dce;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha5fea2c1cc6dee2dda4458cad1707790ec1f353c900dd38b49e8acb61b20fbf183d486dba58c2a3a306caa8316f8623b951714c8b128fa547cd08e72de9056f23631178ff258cd84a41770f6c0d386284b1feb5f73597be5bb379d705a467f0d06f7cbb7a5ef22cc26;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d343d042494805f3f98e5c45de68a3964bad1272e3034d1437f28a977aa208778ee0a456f30eec3869a8b8a8142aeaf8c4eb3c919b01190000fed0e1b0f617d68521f0f8da02e1644dc7199c81138fb687bafcece129b35a55ee64173b97873b28e97714caed404d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h186dbfe3b62cdffba299eef594688ed10d7e75e7773b6bf9deebfccc938b15fe77f2ffbc3e76cecc78a0e079baa34b3df22a3666d0de308b916d85d3ceb8e1afa0483908d0f39379fbb2032c73ea3aaead6ea6b45a1515e5016b4989e3b41595be57356e07701f30d89;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf5626bcd6c9e9c253a035c3889bdfac3c0065da28c8e2a97f2928af5f1f09f5dba9b4b4cfa6e2aa7824951846a8557df68393498ac12e7790c547307cae879d1ee521d844c3799b5fe31475dd518ae2bc3635bdf366ba3fe68af1ab21b8c53e21e240ad8f860bcf391;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e131dcd8fa01de3b0390aa215e90a8f1fe9136119929949338b4d8e6bf6e33684e7e370b378be034789db75b93280b1035b46fa0892c12bbf0119185df462b6f18ec922350fd4223355954a042ae055548c083f64ef13c5a222ee706ac0f5cf189b6fa9b93c21cef1b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3a7983711abf1d32f4048eb64d2f4abc715aa33908c38b828445388cdc883cedf9e6cb3699df633c11e8b82dea9b793422ca8cd4e9b4f08f5b3a5b47f41d07fe931a5c4d525ce0b7edc28e713c40893d90cdde720a55825d0468df605f330a60210d987a71239ec4bc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f9ba694ecdf55ece801f9eccc1d2b12724ea65154fedb281354a8d83d548299fa8a7b9ba596fef4b6163cebb449a306c3f7010aea117a266afea1ba986c7c8aaa211c334ddb9e6a48c005c7ad9eb6a6dc53832a417042aa07977f704e0a9fbedf2566968ff702d5f81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb76f725f7e7fe2a09a2bcc4d03727e40be1b134d37ce23b0b991192366af9e0c76225d4b55d68cc7989ee563ae9397eee71ccb11bf0390c3f0330c3038c2b19241a6203ddfb2891d4154704c0b13a48bc222d6a7ce7abea51c05f7b836e226b3000f463b5ea8dbe757;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h780ecd805b3f040486a0b817a4c2b9ef3d36ddba1bf336d07450e8d8c1bf4f08a4532a1bcc8616393bd14e5102f56e61f9bf6d3c70bc3ee92b75013d5f946720397e1798b16b32385a1a5886576def1266360a3daf5ab4d04978284961185bf4803ace416b2915acb6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c7781cb9d0af59c38ceab2844217042acf853c02daaca9959410f0c384c5fe133438403bebaede682e321c03a273cc736e534d6a7c5db4d0d8c47640217348885e3a31cffc41251a1f399ebebdcc5645cbe2d5ba4d01fb9b19ae5d443590772fd1f6c905cd338db331;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc61b4e3379d822973ced50b4458b8ef44ba4c685b8e9f22442be79cdd053f3b7c54282ccd06b49132d9f3630c92c77ec06c79f5d34c5d17df575a0f63332f9b66dc3ad3746132a278dc685489646d5df85ac89610e9e181d0b8e98aab90334cb1bd9612bb1c81a9b4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19d4854a563d2f9b75960f00bbb361f17cf469a09b144dbabc3172c4920e99672544fcd59295398f7713535adc7e4cb785b034cb4c8fa08207c9149c8228623a5142cc0665745d15d20223d25b9ef8bbd220b2c47f5ca28fe345c194706113bbc2d0c1ee5096803e231;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h176b8dfb937dbcb41490f05b7662864ef8ae939f6bf3645da0cf07cbd1be02f9eee7f3cf6da5a4b2032f8fb23b18e94cd742983da7761a6e915f5dba81ca4b10c9dc2b8c20ffb62f1fd94167d4aefc4af0d33896ef4d32e25d18fb465fca2740a358a6fc2bb924ceacc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h89c565eb7100dc6a8fe63c3c2c58aae1caabdf53985757e1ef7dcdf315af2b4821b70b485c22ab2eaf0d83f7bfa4bc2fcf0d3dc9033a0e4e0d569c3fd01297e363dd2827d0af5dde1c98ed1ae6016464b20d4068cb1b770ee2f892de4db3c6f36714ae8eb84888fd38;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h12864a0b397233e4b3eba8ef8f8fbb5a447cbb10f616e3230b41db4c2348f42cfb1c76ccf5a44f5f58ebb81665c3dcb891edacaa1b26805b378ed9822f122a6517610e31594b93d43733d017ffb169b03d5f4d173f8c48ff5d51b55d355bdacb4486061bf895032aaa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6809b8643c18c432c422d8e490bf9b09443fc8070eb4d078d0c3fadc88802cd6ccec00ebb43dc7191ca0cb7d69a546b26172c94a31f05d421831cf2efc84854a7f0ab04d2d29d80e271f5dc876558f47857c78ce945a836ef760ff91ae95570a559fdb8c9d060510ee;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d4fe28cf82e1766086ed70b541d4e7c54cbdd5038d15a063d82f69480c6676a81ef0054ad19c9a99854f6f1ef1a03d735df13f8cb8804e708805735eab54b4b7a1ef1b65cd1a1d0554501f9c448b8e1888c82b9bb61fcfef8ff36c1ab229e99bf142c90ce96c10654;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7c446301d58cbb04b3dd45c23a4d352357f23b171152cb645aa7d91379a187d01859a9ea2aecf6a6971dc686b924576b97be56045821b3b20eca219aaa26d38e79fed5aac8beffa929588b1d10f1a9c61a4e361890742475d8772579ad4b7d8be6579d258aa65b7cc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4efa7c9a418b7a48e4a395b370b2ec3be5a1be79456035a5030299e0683a8d5066439590db44e892267569428f0b9c022dae48993332618b4a819d1401c048860c27af60bb59a30dcd2869b8a94f43e423e6df1cc1659727e1ab8a287e49796f01d053f444f5b4c23d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1335832863b83a18610d2bedc8be582755c011d4d3b8f3dd6ff9f0116dcb012a0cf828e3edd3426b2d38e39961d5d741e2791ac73c9a50b87f9f960cd330d06e4cdea6f29713d390b026f1985955f6ce732bc4a9a9a0e1982f038932376303a77ba3fb530c36afb7f35;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cec5044f1262d446822c6037b9b3daf25c7bd7e2996fbf0a312734aa24de39b7ee3e1e9c62160497d0145e762930c32bf77d5c29e1a8ae61d6168c4083164ff43647f85e5aa9012826a7caa169047e90ce8b46883d740bc049fc583a0884d54d1efcbc02bd5227dc8d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1087e6b32f787782122376ca4aba238a559144f6fd2f797aec93b2645ea4174a5314631c8c3722987a3000352d148d40e619bfdabeae255ec4af0cb2ffde46536181427f709c745a451cbaf21b68cb3fe53d437d2b382873fd463b67c5b19a469664025ac2a68fef3b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h65d187939e99ede1b1eba062712c239619ac82cddecdb1cd118ce9b936b0dde923b8849c01763cf352502c2f66144eb2696ed7778497a29aec6bc6bc485a71fffecdd344e824b33d07c805b2e49559ddbc54b3527474514471f3dfe2df614fda52657f4fc00527e3dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c00cd899a02368d514ab77a0afb53fb29980d289b984583f51124a5fb86b344c767142c71444104e2245935a21a3108e2d4fcd628f06ad46246071a331c2bcaf61d0d465ee223cf7bf6584ed9e2a0523f7328cee55f2c8797bcd11ce6c2d2ffe4d5e0374d755161f2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h46f09d9a3262ca45a065968909a2f754e2ecddd9ffe7ba42ebb0233fa29d5f7112f12f34295590cc40cd6d79043aba420d7b00be67f8d0a275ccaf66da74278e3b4a9488c21937bd2c9d2296570f3d7589c61d1e36b4966ea4cb810046369cdcac039a3c8d51a16a55;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha76f3e8b9cb3806c7c2f9a6367ecfe51f0059e24efc26fa916b09d1acfc98a1be02d36d8d1aa57db63fbba4d86f1773abe61c74a3f4192edce065fcf52d62b6f6a3e047d3ca9672889c3b0f4b1b913149f39755b59be5add67bbf6af53998c0b852ab2cc11a6b4e0d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h25f99b1b296fc9958e99f49e441cf980d36ebb839b19e93abc9ff92a26c57ae63a1121928e225e3ffdaf434778f555b0ac31b0045dfea5943b23920128838baff43e0f3a82c13a0e50132ac8c38a5062d0fee9d58aabe7bfb8f77d7262c6deb35af1b81918bd692ddb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c75c1f98867c9470239debcc1b205cfe812aa4a16b4c834b9eb20465fb6efb7c93665e5d695e152f4a5b7fcf4395d32252b4cdaad5307ef254e6e9cd3b44920f07658b03a688ef4f2995bd873c2629db81be0f12a17f04e1343b484355ee644a3da581ef518ad6843;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h134fc052a85a0f64da9d26f2b18cd96b046b32ecf79fcfc1ca26ec53661b86c6ca718ae6e5bf25ea4c5887d09e4e0872d54d8e1eab71e7396294f17eb98319600006a5993424023cfdf7528f894f3f28f2e641ce104efb137a39ed2b98d3926971ec7ad7d1e81eb49cc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ec6f704ceac93e8fc1354eedb00dbddb7bb5664e2a811685d56f52b97e794d59eb2a7f3b07ecad5fc0b57177e19ea10c39c1fb6285f3e4ae442f8d35202dc4f3b2771f96522f52577d403c30881721d3929641c96f56393c5d92a2264b69d77beec469469536fcf7df;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cae4ab00c0af6a09cbc3a0331591c09312dff91506a2fd1e3a0e6f6500f3bd25fb3c06c8ce76d7ee6f90dc70464ccfcf1a7624c23a46c5544dc6a072285d8c3944674b6babeb40856e86559c258619139a5d1f0a9211581dcb808bf0dfc6c02d72cb0d03870b732bd4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1011f4ea6471836c708bad57f37e93fe7bd9c98af6f744904ddd19cf786125661fedb69b9401f9fedbf6509ad65d30b1b957e3a1928f725983cabbb50a14ddc6109c84e3efbd37f29dce1b5cb42332d79dcec1a69a16c70719d7799e6ef8fd6c192ffaa6fec42744407;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h31d56f0f4bd9ddbb9497c9d0c8e8459e5047d51557e2d5ae181495b4ff399e6dea6151ebfec765ab91b0cd20a8719c7e1f3ac421680e1f29a6ffd9a7a6a563cdcbb3d0834ea535828d587577317c9a9d20dcba3397db9a2e1a0a2d21abe9f8886d22c7bade95b54a9d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h148a788e2971007bb0ca5efea3da55b96c085bb789ac8032fc4d75d40c7d41770e5b862168af60d05b837732e37502bb7ae21943c71b59e838a1bdcfc132334f699c2e769d1def2cd6a8b1171f80069bcd7ddf8400d0a5da5b32a8a143110893661d24843f30330a6f0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe73edb8bed1e60ffe6620465be7c387a10fdf40d9bdd8328d6b245c1686c3aa418659e7986c5841c1e43fde3c6836b2e0edafbb28a4bd86f7add08db1ff0f7fdd28f7d65bbe722fddb09a18cc32ca5e948d391b4202b65843fa3e0646dbba543cc5c01ef38dc1cb0f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1894bfe21b1d0ef45442a79e1db7187d8f3b615fd0a74fe28e7aff7c9c57d118eb32dfcccdfbe8ad0c3bc5b6e7913e08cf1e21b7c2dfb3809b8bc8c3420a857d369c6b5783f8af949185962490b12c4b8c31fbeea3c21f0ccbf568bf0b66489ee177b0f3a729ed802c5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h91f34028fe8bc16082aa735867d92c4d76b44996c25c616651321b85bb7014a049c02a4c1b7d977a6a4d9ae0a952c9722e7f828266a7cd0b083367a4cab0579d4eeb1abc411c225c69979ee2473a4f7909e0a0a11c300b51a78fb69b08e102d425426ab9590c89ba69;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8420fa0ab6c81aae7e7fdc5f4d18460cd02136e1665d8410a09cb876ba64566e5e2151594f58a5708db04bbe92acb7edbebc3862fcce7aa56884ed4c6b40d3def77cf471000c779bc8ce8b0cc2cb4580b551e96b7dba5480f4c414dd41dc1b02a9d3d371b2ce1e7e81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h156258fbdee1e17a58822c618074edc7a62b00e20549546a1274101a3a208c62c3744fd1d789aa754153f422a632fcd65108f857d30574dabde93968f7f1a5a367923b9fdb0a5f73c8e551b64b78e98857213daecc4846962182b72d6eb405deb87f385cfd3d744d0fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he3c17aff94a3c8efcfd61138afc1f8a033c43143a1b44a25833a61f6a86278ad4b59ef92c659c38a75eae4b522c7adf4f358c1f1f49d8305800c8cc4fe02f6b7c23cbf821ea7a1728e51ad2e350f1006b24d3aa024dd72a7e7cdc4095a76140c2c24ca062170f98da5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd90788bae8d4f6e3fdea819c38abd0e6521b15385a1306d141276dfe1f20ae45499136b00ad273359090f69fa198c4a180446d9ff67903d0eb6c145cb73d22ab484508899bb57ebd4df05fe0a8aed16ea7698689ff0ce496705e703902ce06559639c296d2e272fc31;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha046daed64b3a634ffb4ca101ac68a66a4ee272c378124b8626a3f61872cb38eb9608b0adcd75e5abd82bc449a9f8b4604f81cde9636c60238f370f3305933d0dc98eea50e046770ab7fa1e9ad821d936c211a2e1731ce423d196a9ac0f66af1cbba3f82163a452217;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2d921688776447b2e7727e22af8644415df99b88b86d8885134190c7b8abce21526d7724d43c4da5d3730e5c7c9c389763905676cd6a4c5f5d86955fac836dc7e923986674289178216d22bba77895e09aa7e7ffaf39c84cc8c414dec9866b66f490fb57048e337808;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd246810998ad3c1d596069f2b615105c2bfda1d60b874210d2f86efb96bf9a6478869386ae6f9b4449a09f26fb837e0ae5e294c7510f88b4a287daf5365e6a068489727944a21f9e2520c103b00d3f6a3a9bb6316ffb1bf86ee9af6635f95c4407dfd8cb24bbd871ed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5e1369b1e46743e1f24d88bc0ad3874542538a5a72e51e61f62fbc65a016891bb9d5c5b91c3bf6667db517bd1f859d38c2fd3410db69ddd353f2f9908792bafb60def892b00cf35e9cbdb9d4672a39763be7bf2c09a1ce8d41a0d3b498d5827e5621120412025795a6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4104c3e5d5a17744d01d99631c23e05815bdabf24e3776e582fc963e6208cf03a877d1da6a035cbe7572a8ca4f55e586b72ec4b58ecb3089ae2d5b21efb1409429dbe8f8b2a5570d9edb10bc92071f159496d86cb795030980346ec1c8acf65a018e5667c5c9cf2223;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he61bbc14e63988d5501f4fbc5d3ad430ca6bd3b5439e28986965ecf0af0b4bd3527c70825ad4236f2f83cd63354e4cc8566aa7f2833dde46bc7f7b0fb7b112d1f1cbfe719663f527028ee2925959bda61a07695db43224f97d5740e8e45e0ee8d12f09eb1b67a76fd3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10c04ef4e6ba179b8a864fa7f841c602c3aa04f12cc36465930c9476973d6998efb8ff956f731ad7672a6d4f017d87cf13e5c2efc60e0ea7b8bf33197630f517984e483714c60707cccb8ce577a84dc0e2081af4875db03d4190ab49681677b4c61e7306e136de53ed5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e2b67266291333bfcd1bfe0a61f0527ace098e20364f8faf2772dba7c5f49a020e868f555f870ac4eacce5d010f1b47572bcb2ba8404f0649ea3c6559b101dc1eaa6436b1202680d627d88f8455f3f739b81a8b79772b094bda03e11416e99190be8eea376d86adab6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e89d65e53ceb54976ad26b667f75985933549085081f2d5cb842a13fb377f7905b30fbc11ab18dd46f65f69f28adbfa18792e238c5fdc2da9e08f3d2253cb3f020c4b41d544bd25754146bda5804a13800f5d48196f9f5cc068a9cc76e3a9c943a606712918a44d626;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1adb3fe37539c08cdbcf6164ca445a17a48ea939d6794510322b5a4843b8af4929465564b2c9f074b44e6b1ae10adb6d659fd07c78f8ac7b003410ecac4a3c958af10133e7842b4a36d3071bcb526c96b84d06c7944d4549238be692afc6af9b740df02e79768fd39f3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h47e3ceefebee26c68392af7135e89979efe3fc5dc9db1d3ecb5611e6361706fb3b8108797716eebe5c87568e587ca894e5f86e23e152ba03d6ee4d82befe73acdcd2d28ee194fd1b23439ad858db3df98c47855e7a88bcdfee1308647134dfc77faccf5e9b9afe3ddf;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd722c565792264567ade02340d9cc21d3eb3cf2e70cb8ba9ada3f95e267ea89558aa7973dd21881cac611a6a37cc640db59f27ee9a2e29efaa7f99f26bd73ba4ae11e116ce4ebcdc62a58f4eec0b8ab8146168c219b96c3a6e506bf9383336eed47de33fce0fe6149f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f4213f46bc19996818e08cc4c0771c7d2076ecc74454d93bd623282a94200a19685b19669c209daed6395714f485bb72ca7c1730d2422451a1f50de961d2faea4812e239a5dd0ebd35c856a29930b076ae47f5e8ec49e559299ad794de64bd70b11c279b234bafb0c7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbefdf3e8f2c5e1b004b34f2fcb6157ad3a25d496ddc6544c899780377dc30f9c8b3a6168d88a7e571b44229b5312276ca3da211bdaf204b012babae0de0b75a1f55b8abec8661f64cfe17fcdc74c106f3a525ed1448dd65c3351771eb628ad8b5c8f491da2736a5830;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h98950fe28c57e472146bbc756491ba68acea1e4692460a2ebd8f5122b9a1e96f0206dfb20a06f88c2c8efb448305dae5a43b041cef0ed24b2b186f40c423725126a490258249a25cae766856b3c24ed7038fe9704daabe94907e657e335621713251208647cb30b66;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d386f7e475036919fe03c238f6b71bf324fc40cd0ce31178350e63b3829bce0a59efb5084af8c65fbced843b4086f863c054e12e324b233a67cc95385d99201e595ae5bb5703c43cfd46a1d480b8a8b5afa2a64e60e1f3a1f495ce49eb07ddf19fce3da884fbb15940;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbcd919ae91eb652645433d3c1111b7ce380d215bafe397cf20c9ecd3e3a539d1d96047facd743fe6ab5833f6a1dc4f04c768974f293c9210dcc654393c1b9edd04d2a666b21582c80852874e620a296477a9928b41002a0942ea9ab3a06a46667a8945036a5119bc04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h192c6d795c37b771e199e07bab3ff6e82c9ce33969d2eafbd55faefc5afb2fddcf629d7b22cd96b16e2a9d2dbec84be7642eb2a5ff582ba3d61e3c12a1f21b9ea456c0bfc939e36137d961bce10ae037654b26b274ae1a5194dd02c5819d2335472b2f87af28b3bf3d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8edb0bf9f7fdca6fc598281ad6b8878fbedc80d5374aaab98cae81c06a443e4df7f5911d4d02600796e75640de3cc6bf8e8ef6a6e3316557a464001e0f9b6df289e4167b5802a87dafe4d46005302ddbfd70be6ffc552542c3938e439e7404b7cb9ed9b75cf1ecd8af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h121901e5fd9e5390e5156fa8fcf46ce3e7c3ed08d076542e852cd088940a1699fb75ca70e5c34a920f407dace6c2c89bbf819a8698a0b99a188ff6514b6426700a17cb23a71141bacd5b13a42f33852af8d0e82eba1af49e9e9e870f7676389f9a8257ae1c1e01173fb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fa9a1b0df6644bd5ae170db7770a5cdb97a146c4e36fc03ede469f328879735fa7c6277a6fbd93750f75cdad2774db058b63f858e287bc5c37f2ce02ebd4e0ad9010360d88920a62cfcb5c53980d9b65194a3ef6d4470e44500e6dc3a177111a2eb1d462fbeab5e722;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d4ed2773f99a501eba9172b13cd3c5d147e5c03e4a61705723b0c2c20495c357aaf3b4b0213b750edd3e5023c5e87aeedd2b77237d7046e375197ebf3e8d29f79dde6b36e06fc3a06ea4a261303faa2093885239e55b48d34117099a75f9fa3d3f9a4e008dddc61a53;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h156122e1cd4d3ec564d89116e52a3779ed8c660e262b71e487d048fdb0d2252879afde4d2ad3cfbdb868afaafa71b0aae9c7c1425f091359bacc02c7e010ecb2219c3fa85fd8c069f622d450a8be394ac377bc79fea65068d01104efea17b44b87200a864feb782fef0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19e2601b66868f8c076d421ff5ba77ccb689ac916575af8a7b596938fe88d176660856991b7bf407af27bd976f6d828fc42a02bbc4d648cfc3d0e43ea71f4ed0a86f8cc4e27690f4b29268873cf861945e4ffdeff44fe7c09fea59fb2a064dee71ddc2416436157c4eb;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea5f62bc67c84ae99e380ef6a62d476a2ab3bf276dc7b7d6667891e7526e06cc423b3781530be291aa858d8b1cebca429c59356110ada00d1acf44b915d26320e331c3ec6f6cd9dcda8d986035c1dc321f9288060f49f3901e5c751a7969cc7fa221b62873472915d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8435074dc42b06fab136b7045c45f7609b078d326b47491ca3743d3d8c56e6bb56f03f1d86116b335078e5983d778b64c2e24d2b52ea367cd18bd9bad41c502128c265d87df3ba9b64fe79dabeb6dc3b41f178d41838ffaef73d7cbf41935b5216847d61ec3031eb04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he101c3e42707c351f7975848cd42d82897c9f71f4ea133fac046afdb7908c63924264767b7f95943b80f593a78bbd3d57717fbb0787ec1e75a3b82924f8a87ef60c8505f9ce7a5ec31fe06bb8945a41db96f75313400b2671a0457fe36298c8be5cf07474cc6bbe810;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18ccc6efb66efa0918069cc44cd793dfe973d4d7a2c8aa1e20e515dd0600cac6823b992b5ff75c93da76ffc4d8fdccb20f125b6a231c5d2cf31669eacb50d485783ecb60f8b5e0d804e9d9397127ba1e77e116c77a2ab19795e6d251776cee04ae7a34a0a944242d301;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f560278353349ed5c7c7618d75735be01b9c4d1044be86dc930c70c5386291c6b772fefc3043dd1074f2b3c0f010d9e473742eaf55165e091afe67ee01436aa843640e95d38c4f06f6d0eed3ce6fcd86742c0d3e4c760906f31207fb966068c2c76059d1765c878b88;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h7b22d66a368c9d3b0ad79f9ced3cfffcae7c71fb611b2d65ae4b99008cf2b4aa740b65cc7835c2bfa9ab2e5c5812643dd522e2e8aec6ef2c0070351a3f7bedfb91d1d6bc35a37a4d9eee06bd817b7ff2be89ce170348a0bb370adb4708f79495fb279ed25ae2ee43a3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h884aa008c09294b336bc4f2ec351ee45ddcc59c2c14dbb2f66f6c8e242c3c94c7098d4a56c09dd7489ebcf4ec2740750e40b98437040d9b94d33f0ba2bcb376e148b89abf88037d1d326a0c4b2bd46a18042985c0d34c6e3abe24b2f2b6432084a1698e4901a216e32;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha31f211f9099a6a41524452520b649d178b95e94348f68024dfdc2d91a0b29bf471c79aa5bd7748d6061024a7ea3c35c56ac589bf2328f632fb95b3c676a53c40dace3240b6a047a8b6196d3a0c2fa2eed5c503e4bde42c4ee0654bbec510b6623d2c0ba98d930ca33;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1fe934a5474dfe8ca855ae3864e90e91fc8aef3c245714faca81ec4fef4b46672e2412b17584e3898111617ae25d7b06009f0180521ad37b37f1888596b7e64665e495a760f2805176c2cf2e86b8d905819b337d89470b6b856e335b017dfae9613221e3951a0a319f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1449c18b4ef4e2a959e11c26d57d35b3b3d4c9e89f583731331d25a61742bfd6d7689a409622e08b823581de32e7fff30b5a869220a634d4fcf302888b91f3e624fe153a5b5584d18fbec00df49ffdeec3e42aa98118068d2641046f7660cacfb1b657f5966ff664aac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1364889d1998308d87b79d0593431a90378e295498228bd85b4e81b36611bcb3b9bca0d1c86bb4069d0b0bc4fe5509085dc3eeaaddd7f7151d21bb7c86d546295e4f6ba4a2f4fbda7689b8a6f7068ae06a5871213615265be6e5e1f981dae01258911a1a4e3f9258180;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1dc71f42c47c2088dacdf16e01350a33d7427e90852cdaf5d0961c80197bbfae266b7d684af9664002234c81f83a05040476910a7d3bba5b76a1370dd7d2391b447966ee20a23de5be7f7f96f55cebc9082955c521aa906278ce3b9b39b0edbd45980b758282cac3ab9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10f962702826ebaf641f31a662036926331cc09a086e730890abcb67145976782306c3de1ba3c672904a97a792de0a5841dee6233086bcc954c3dccbf9afa1349315fc61134ef50995e5e0ab6b5120199365560d12f364ee8c87c3716efe3bfcac539d21122ddabd6af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h698e6e4f6299e55220bfa773d37db5c1cad3ef8c472a6fce4f1fe626907449adf547e964520d9e23c3a368346621fc9be5bb07b11a2baf050e6c8b2e0e7ccd9c13efe3ba429652cd6d0c0836bf6ce56dcd488ce7b14d2e1f8e931983137031908c024cf4b49374be39;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54a2a4e8310007ae870b24d6856b76238ff44aed5e04afe2a89514c8c056d41e2d0a406b950f8b741e95bfb415e1edee377e483bf58dd92addca3b239344d9ada4252165249f2df561b3c5716aadfa49a20cf6d11c28ea9b8a56d783f07e1f31b162dd0519d390b1c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h24e8912160bc5696cbd55cef07f36ea7c9e1043e803d121716b3122dfda66601f9226d91cbd8e72edeac009e1ac3b83ae5d3372a96067406b103da46df5707067f5021628d89977bb2630e9375a1c712147c7eea1f6af2e1486ee419dc5ed7de9cd01892fac9564b1a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h597771d6256863496b8fed045f9f24a684f8cc98e267981de9758ee0dfc4b96ba85b6a87f73d39f767fec2898e99e65ac72f0619cecf7b7016234806c9bd564e11682d4dfecd282fdcd43a1f9573b5fea8023e8768f45556014a90c1bc10eb22988788b1f043360118;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h81bf2b692457dc58b64602b1e53f00f459aafc1518969499ed128c14ea87933dbeffdf1d1e095ff1906e97fdfd129b8c3ae5bebbaa7e92e723d7bcf84eb16afc723240ee3b8a2d9c4de9c54fc0a3a8cba21013659093d9bd4086852bb63ee075843a1b10e425e28ac6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h161bae09182fb841bd7d3fd31dee999e68883f66ea944a879a8266ac44ecd9201a3db8372a1dfb0db89dcb40974588abacd3c07dc7caefaae3c0065377d926fc43b0199b38c28373c9ab7652bf1b99e6803212915278c9bd1891957042e58a08f665fe1ae7ddc223c6c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b01a1ffbfff11e5c1610d944f7ffcc92a11497e3253a90574dfcf072a63ff836acc86290276b519305175d404ebeaee4541ee17a0bdac3569a2de2be9d7a9668f7875752ef858a877550ea501d9e8c3fb01561cbaf0795eb416d0ff771a51b9c52e3c2b3e37e823b81;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6d8c85af6a6bb2e256456643b4d83bd56fcdb939682cdc1a49579d61a6f27f3f3f388281f59f8ea87c97881f73a4125174d45012cbe7582180ec0d9ef0656ffbf1036ea2f2dbefa919ca2735586747d5591b146f09f25145e58b721a0b46b3f3aa9f9067ed8e6be14f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1be3230eb8427648697b439ab1f6f47ff049da885b443998ca2b5c5edfc02f69327b0a1a606663569cf0aae05da6c6cf9ece04906215cb81e6f97059d82ec80d3be94031bdf44f165c530acf157803e644c75cde8905e49013b21c3bfa5aa3ae573a631bfa4a5ee7cf9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h147e05b1db4ba54605faf4395179132abc6ca0b9dc2fc388a8296bfa321319ca73f753c35d3f243dd919bbbb50b0035a1db51dc3c1e89d1b1391e61eb8aceccde5f314a8ec00e31ff10d5de654ecb53e59895e757af5670460e28df51c3be812305139a578c07d638b1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h123803c91279c2486eb84a72479794fda73ed2ee1083ea7724774f67f9baeec4d6231ca087b5e5eab1dc4fb7ba0bf22f0c26b602c9986bf0e401f926b0b6ad210df7de18ba41bf543d567ccbf306a3f54ec3db3718bf1ca947c77633b7fb3cb64a55f8b1fe3e6c7ac9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h190336eed3ec610ade47687f87ed11367d770f9ee70e66d0abebde5b8bc802109fbacbbddfe3a6f3469933e708dd7464c2c3d976fff4bebd234206339ace5b4e2975730299a556aba38d1f433feb4d325e3c4d65597d0160e7d81be6e637b6db82a91762e5f5a34f60a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e6420b549ca74c01a0ea2437d28c8acd255156433895e3281aefe4f942f7837655449fc148d80e2255d1cd4a29de2826d867631165c59dda31760b338052e1261fdf30129f81620278e99e9de1fbe130284a581c99043b9a001f97fc1c72bc9cea8f74ce8e2975616b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f51f5bfcb4456bc1bce567cb492f78f1bd84793b752cf557e8e90d7c536967bdd5a4778d02515adad75b995b7244ab14757f6f3334867e31eec3650e82a75d7b1b64238adcd69c57769e9eeb5078f87804c74b2bf6c5b2ca56ef15660ad14b0ec8e83e66562525d416;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcaf65b88b3bbb5e1c7e55bd790813770f57392137562e6c4d60eafda641170e22b37228ffd110570c4d8689089fa7e6f7418f89fe64426b4f99b0bd8ed20f16be675530d22078fac3b4d8bd434a0dab3517dec9b012a4cc139ba82aa85dbea2f348156ddc8b261a3af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h336b4f7020760347d35f122c63b0719e3cb9c95d48a91e44ab31f6e98d0b5ab9371e7df610e38a4621b9a06f4c87e650d0ecd989773a1ca65430f4405a0a59e8b29b7254e0df03ff709ad6537293916905738a3508553246801cf8d2638eaa29c915e7acdfef1ffcca;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h133bdea89d26d8ed3a834abfe0ed29ce21d42c34cfed7f4d874d40c982abcc5a58d3a7fc5b714909338105bf2bbdb59f6bc05b13aba17324320cb17950990ecddc78aad2c6e90c601c9c462d11d88c6050e7baffacc535a0fccd887102a5dbc687d3dc1d60bf46da427;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h43dc6e35d5617c3610a8b76e9463005b3ae52f315b3f8c37259e1be3c06f8cbe435f682f858dca54529ea2057f1c4ab6be6c326abf870f10969a3a227b023e9b317625ab440cf41b86daa83de8c99d8d685c89f25c059425cee5b0089c553dd5e8351c86babc9983c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e3f5d42c59451a8eb208b71266070f89dc702104caf4820c1a0d66d1f72b7f4c6e804c9a5c7d2837e654a395d7b11d01a7e20260d0f79f457b364681663a75a0ebfa68ef17c04672e21a03487c4395bd7048e1cfe4b9f680492aa0d078d971a2846d86552e5cd26302;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h277d899c4de0abbc1f081650aa2a61cda276f4d599f0078c94cb66bc6d9142f7876ac891b3a95d8863ffdbf800d9aba9828408717714dbbbdf431706f894ed775844bcf86ccde9dd4f763b9bc2cc7ac50898a96a1c044f3742ac053f0d9a29c02801f39f8a7cb35233;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa85078c286a62fee03e88b2e784f494522d20d4c2aea0411f44b26f71227fd2735e16fe79d382dba1296dc17755924657c7ef4a67aee673b75592d28ef56b009d4627d3bd24fcb4fbeebcdef3433f374e31ec5efeb30a2ff995b5f050f30d396f64eb83dabdc1ac3e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1877a51f646c97b7dff8ba419de931ef16c754f874075b872f9612eb3cc7ac94716353481ec19e4fae970e054a72824265d18639b633bb9af7487b737c5fef194b6b0f97bdaf8fbbf740e193043ea2fc77cb814de2332d1c14608158094ed5ea98c8e0e00d7eea9d165;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h54f91c93ae1ea165be31cd033c5167080fa0894e0e6513dd4aa945ddba92710a71982e7aac835dd51313aa542bed435bbc57d91fb5f9f4f04418ca14cb33189c862222ef53a05270483b9e69d4d594eb277ad25d957597c3a81b5e176d48681eea9cc4a0ecbf79f17f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'ha793390a902ef81fb2c798e3f5a056bd4e9e38e5b218728b1dd5e326976141dc32191fd974f0b53b8c9872c48e09d286f587035e397f025f212be1efef330e4cde5c6bfaa19e643b4ddc78884b626065a21b141b43edf84522684b102660e6b268d37ce9ccd98f4ce8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h19419cc1c2dcc68881955ed38e988a85b042a8219d09539b5a6ec76c57ed19834ca29831aefa430d57afae63935e2db2f0ac7e20c12b12f41d920c6f42f5a815ecfd88c9449faa53aa932602992f6e837efd9b78d69b35c302a561c60c0d4b7c1840ea7cdf62f6736e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcebe74258111f70e9527f4b41308864fc389c9dfdeac43af899dd5d7cea08ec6dd1e1e7bce200405d3d109d915248be7ca56cb34659a2b84378903b33fb92ef290d92123b3d6d6b72e83fc3c537f01623d7c0921b7405cb835baa82d83d591735b6e9b3fb422b4c4a2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf8054fa65491fa0bc0f4561ed3aec710b69810618007715c2b0281e44b153017bc7246507ee268f0bfadb8cbbc53fce8076b897b8e5c0e396f57eb26ce3e87697b09547ccf98f5f837f22f1d6d820c215d58947f79f59d4881bd5f81511e8a2f85ea19e2f332efa728;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb3f70f2f42ca776e1d7dde83b829f1c6b46a21321c46cbcbba626b447898545e8d7a246b66fb8a21eac68966717778790606304fb40342c2d74c2a7e8ba88939b71ec926dba3ea98378bcafa883d62810dd6a0f2dc57c3a502a2b60e83133a40c9031cb44af2087f34;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h772643488e75e219a8f8e06281110eadcf4147ed75c84a2197796446048aeaf2c57abfae345f7af6174c754089b6cb83a3d0408ee70cb0c40d7d6ee748fb70ca254613129f571e9d05c5ebba2733d7f4f7c6ef7df97dd7b7ffc2d4dd32b9849be3aa56ae20f7856faa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1244a99a3e20819d1479e90e919906b76ea04f518c4562371de28a68e306061d4c4cdf0a79e0e10e7753974987b5f28c360e7b3923417568fda0596bbdc0f3503137a8e65a7ab221033fee9ad8a574b10101def390dff6a59b7f5893a9ec525d902091219f7b75daaf5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h67fc48fc13fa2367eaee5fd400f5e088e64ac2cbfcdf58b607d24993913caa4a6d9b4cfa4874790c7580c149a03f690a2cadd719ab4e609887be93117174d878c4bbdabe9430ad4000c11cc30ec8d225cc559fb1a34de7698c32d5eae9baa522858d04f0b7b5545f91;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11acd0d6df65304cab28a7996487e9457cd926dbe9e88b774fd7a0030200e96fc153e02fecd63dc0af278a98d19c333ea464d618aabf91f2d6567c4765bafcb6aaa6b5a2908fa4a495a504859956174a25aca2cd9c31a79ac31fbd76847479b69c3313a8ed1dabb8752;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h5c267459a4290c3bd69441bb6bd9741221a262cafac6a99c4cdbafdc746f501851fd89ffeb8b5ef537f0d8ab60823912b2aa86dedc07f8797e27711b420ba3370082ebb4188b0c10715626a9ec5d739d101bb482f26c51baee017fe817ff9c299f356fcc1f1a47bd9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b130ada8da4ce49af44598a7e9ecaa26d1fbfeff6b8a56490a992d87e9d4822811bd4c0b1ef16dd44e733a1d97ab964c1d427e7bc0ca08bc3495087092c06ed317f51a52caff28e6c61beea55de89fbf8d8ebb901dfb9a297f20aae514b295764f954312d6564cb08f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h80efcf56ff342965d01a4a41442ca6abd01ccc0e8ff1967709ee92cd09937f79705f0c8cb0b260d50144f187525e31f6c496ca1934657e221731695f1d9426d5c90aa94587e84043f66ee8c50af3866b3ab4dd92c89563739c25fdf6ae647756aa8966da8e5ee1e6e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16c5008a9a7233dfe1fcaced43536a2e4ba74330e0a950230baed9444bdcf1434af06d625d305f34ad91b2021f97ec3746afca813b168deaa7fa0b87156f84170e15192f08990830ebaab5a79e52a664ac9fdaa4642222159a4b98d14fe11f799550234f2d909a9906b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h11b041d601a04013836000ff5140945383d8a93382edbaec55e123de9c0bf16326ad834bdc2177482e853da168b728f0639aa1a97d75a8079506250891971f405b06a626f9fe2f1f9a1567d9d424f0eb531efe8913e74724d845aaa892ed5b777fbc4cb49ed767eca04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h6101eb8151c5e524f5f7c091338da68315d6362ff8e0929f38ce9075f5a4686fb15f89d19936ba256495be9a1d30e628970d984d02ae5681e679ba21bba773bfef02d4987ecf081a2920520a7c4f9a18273fba18f94cc0457cb1065c99a133a4745e12a02c78c6cbd5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haaf738e5152cde4a84b577d73c45ab1b2b35b859813fa30c9a16d4999a448e0696d8f309fdfd5ec27de217b3311c5a709a64345a6ed4daff8328c9fbca02f801d64503a213276a6aef0994574fc99a9514153e71dfc21ecb274b9e5b9cce9953f3f5f45f1e5baa2799;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h36e6d1db00661ad88c284bdc3b70337053021c4d38485f09d6639dc39467613064af884f3a261221711f2e18c69c6a267ab8b981bcca2ce6a3182306f117bd5f60572b443addeef4d65b5726c92eb273f745dd35ebf7f3e425faf34ad6f9418bf78663e6f860a41234;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd594958e2b14c105ddbc10f8603a08a2f662f0a3326f6c70ba009a25699f1c6d5885b141db9871111d30eadff9f84a1926e3e4922f51ed11420d1a47cecbc7416caa2c973b0bd44c3f43c6d3cd39099414ef531239fb609732456d3d26729d096a911a16f652111a13;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ded2033958ffd98b0d2f41484e7e6a42fa959c719c047dd587c002ca304f2a03bf939ea08ca2a792eea6404b0d0436b417c913c04c7c278d441a4a8e14a45858671d3a6a5fd09e05851b75d921d4cc16e612e618ac1727af6b46816708d30e1d8348716702bf96c380;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d932e2cd2a9290cc3410942d5670e2634897696f35658225033251ec216b2877bb6aba07478b818490c7ee1838e1af01049d8e6924b228003779f72a2334a66cdde666d65f0afc079db05d3ff4f8bc796afb093ff2b7093c84243fdd3db0316031589da82c66cf9e9a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'haa8d8a523d213beea4462ba824f0ddd140b51f2cccd0686ebdcc2c4cb8a2e8d30af887a38971739515476952bac250514d8268ed34a21e871e58db073eaebdf541dba20534abb47de908fd3f4ccf849fa579641f39380e9738183ddc489e3d4d820f0336faf6f1cedc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1464dc7bb2210496d606fa6df368033ea3a0735e8ea63a4f90aa3a6b87f950a2b2f4ecd39e3689cb503c9cb0e52af6b3019a7f6db1f077e622955616cbcbdbd0094f52c21ef0bc3046ca2ea4516b1dfda3adc16d2b00880d8e3f1ff054e18a2cd7aa5dca21e840de184;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d866c322fa0a46ddf5c2e32f51f682bee8f2f3a48248c3563024ad8da881691d9a42ebb762e76fbe28fa14cb1cf25d0e4faa88a00a6456cd2a30667e1a8527b032b2d288d3f4f8585f338105481801f250ac8e58f18e3ab1fab2c35e6a2cfcaaff816b30a7d65f85;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h143f5398ff81dc6984146d4b389b165a8c282f7c2dbc8948d0712d245e4ea5e8619d1442a8e44a49ca26481b31cae05f1dc88b98948cce598b1361bb74323019925ddd7b4dcef3dbcb356d898962d86d3dac4ff40e0b676c94648eb6110cf57348ce39b143a663f815f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16d5ce9d2a628c89a472d2a60008c0095109d1c234bd1c32ab99943adce55206d5f508585e5554dbcb50eeff17077448ba57c9fdf6c23eb4b0edaf3d28cf9e635fb5d29712c838eef9e197e173f1e70a023b8858bb5124d2b01ef039865957e492174cb1d890462df42;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ef8fa19468016a09507929e07c33f37496d660796e679f49e658344d0055218c21f227dfcabe6104e9d465511e1775eaaabd0df1ace46e1727cd9b0f39335596370d6a4c5e4b1f8726856bca4640ff8330b0dfab1e6b8e9d7c6d9f0fc9b125508541e7523725174d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f8317af2d3ce52ad5615713d9edff45c5a131c3b6b8b72d5f4ac733c254251ddc659e77067e0bb6648e1f452b8bd7b199d0eb6d50136ac4fa29749a7cdb9c193ab62115924136240325558cdad6a3395c12f4c41040e39b63751bca53a8a99887b85b7fc79807e0103;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdf387c4414a6ed07911fc960111d2db6803a0b9d0da158b0e8d82f350e0e66a345cd84884fa728e97f064b8b788340b5380f4c610ebd6af6779b3c289f107d3458b17fc343b70266bfd090d6f66e88a77a20e26ccbc982af05b03f177ee7cba7923cbcc5d339bb03b5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h73995a73d5568260a5b2cd2911446371150d285a9ed6ba2568609a5679469f4868d9131f838360771ea63fb01b2a6a0511f67589f9fba3e7fbab85efb9e09c761d97df988bbd9d5fd59b194fd756913bcbeacc84d72c36ae932332c7b11bc4658240964d1469b2c08f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c4157da1991c2b5932c65f9b6db7d8517fa4e59495ad47b8f1092370aeeb56d07540425bc7c4ba1f69df77aded31e141016ec4a0c2130a2dbe2962e6da15f5bc6dc32f9dc89c029571c75c65950c79769cbd5a1ef9b68c15c5b9b5b6034d6b280b2878b1d3be018a16;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h75c1ba92d63f7f8c810cf4e763ece35ab1921dfd7865414193df195924fbfe74add28534d661fafe011d812e1d4cecff5eaf7be89866363d5145422bd532561b3e14cb8719591c17d1ca59a7dfd9497d9349eb506b205187342ab1ab741848317706f3690a48fbfa96;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ba41b4ec02d560fbb2fd9457cddd79c33f43ab84f96d35aa82f386e23f1e2c3242e1ef61eb29cd5bbea2608d9de2ae470d646316eb529c35006dcd3e5de29f168e6571aaa83f89943bf55ce1fa9384b9eaf89e1ae527939456d3b6d579d329aacba6ad95683851c64f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10d79f455e222189f8d7f9c7c86d6f96e40a81555c2317c7fa29c34f3e96b6b64008cb70986302c2d71992e4678dccb0d2163160b41447fd40d474ba9822fc73df82f1bc65ecdcf9110ff3e4ab7cefffa99539a5867bcb4aeab690ef524a2f230f896e6d3494acca90d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h119040e70cec37c9b4439c27887fc5c3727eabc710bc089619d38f167c2af8edc98f10fe4c7c031965b095386f2137fd37d3c66b67d96cdccc7c0f4bd15f4cce88a67e77efc6fb82b2ac9cb85cfc01dcb307ba2b7b6ee0ca0b42c6aac47448cd08f39d3ad4e44685b9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb908ea2bdfcf504ad17fda61258419537677404995cf7976e0d700b362e8980d092128da8b8d2c60802f9aec1d6f8bf995f3334fe8911c8276b26189fa3b010b3b0c6ea2c3c73189256e1f87ed200ea57c88dc2b7a0048f318e30de4f6a098ad2f8b6c17626f3b30ac;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc2ac2fd325ca5ad7d7bf6dc6a2922dec9a610a0702d5ca5ce095d331d1b9c01b9f7d4a4629d5d1b53eb964cc21ebab64416e113d18b46d4021d8f22a0d65f4bcb8af00329e574ffac9e26b18f4254df9edef9f5e446148302fe1deee2d40d5740ffc8c94c2be53c7d5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hcb31ea97b04402ef945bc7af7ed7c0274408cfad1a96d599e8ae74ab232cab55b8e62ee45a33b493dd2662c749daebdb193d4c288d55dc63b5245ec6ed77650523c23c1ed68065b44705c994124255c4f49e13bfb9a07f5fdf9868bc412e0900a1605b33d60f25b5a8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h809dc1cdb685546f6b99816d49419c026a43f252dcdb5d468ba4f246fb9b7aff3d814b1b27381fd9052246b68ea3fa01812a6340279972de95dcc21ce3820416777dc0e5fa25b0d539f489d3f9fb97331b3ddc01deb6c05635b11bae4f551938947bc296222b70d903;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13e0e9d321a7e397a6940fd7841c2f0af2a8b766eae2732c1f482d58d43bcaed7ac8e939aa3e7af7e8852ded6c4cb807d7d2d060493ee227527f087adf74045f575ad7c32321d66ae56ce85e9928c12c48f943a37860a902e7a2c4f1b478715a88c0ddcf8e649ed69c9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd496a77b5c5807bca1aad0fe3af24b73e269a66e31a18ce5e84e7d39f4e0445ce0c4edc75b35877c51b5a4ef24999de1b73495d5e21452379c32941afc9eec70e867ba5ce14d9a31b9d1896f65e581d17add2f6cd0ac43af01f94e49d902e2860aa744c2f5dc264ced;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b1d2667f36dd2aa1f1079caf8ee58f8c215f5c9a6f57e7e397f9f548c7090d570e2984c7182c26de6893ad9ec3608244653eb2de4b1a689c3aa101de91b3d4117094221ad6f62fcb804fa13853baaef6fb5e8591c5cc5ee2499723ea90c6812d1c008d8b1c9867a1dc;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c06dbe8f6468c541fce76139cc72c8359552c0eb96c862ae68d8dcc1af10d8f2aca69cd9e47ed1d9611d32e793afa965bc34d8e2dadcf596d02292a35ce2e4a6c09eddaf24d3f86759f0bce5fdec356580147ee2fc3a167270d9285c2c3fe5bad1a3440c7924bf1390;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1d8a606cff3ae56e5abacdb6ca6f86e9b7fb29d2edeab145da054412356817a4cbe721333fb3a135065842e6c58fbac01eb63ac0f3eb658a1e75d4522429d6419d78e7a027f124deaabc042e9d362751f83f703aa3dd5d8b638f90df8fc001478f0c73fd024f79adcd0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3faf4025aab2ece919f5e626f4f2b5806606a75d930034e25c6f09fbb883d5644b7b51390f58c99fd1698cb17fc747a7d8bcb232b55115639d79ea529836e6e0249526832e4061d536793a93dc8ee17c4fb7b9d063312aba871a32bd105dedff0a7a8df87b43a3701;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14dda4164929c4c0a8f8143ba3da6410b4fd6e8f12ca1e3ea4fab3664ebe6f4cc80453c7c004fcaa24225c1aebc8d0f10368fd598835f918c18b4129341cb312d50868ada67ac5014c7981da3322ce313d00c52a48a1e674d85845d30b695a61038a278f993b5989b22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea8f0e3f8eeb7154c14894aca0c60051f84b9922da8d3426676887613d8b3dda4d6cd4ca6ac8bae438756cbb6a105b57525f71aad89b4c695492977dd9e87d85e531b7975d824ffa1f3ab857604481b7f94d13d155961cf414f2efab4e983173401e8aeee301533c7f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c84fe5cc304c1bf2dc88c7783f31ffca515186c3cff613013416f9b29d96655cceeb3fcc96e9c20138eb8b94b44753b40b691bf7f5ce208fd7d808a2819a878dd5f89109c6d77c2e45dc66526f6f333a9a403dfe7e3637a64531848dd49f3fdf378d24c6715f27fb93;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13728e1f6e65cdd7943270c92e6968a97b36eafef028111127d0f8aca2c05502e8fa00cf5ce3dc2f0ea6af1b374fca2bf29d3b7f4b3fb90b315a4f12bc541e2dba579890dd2d15740dcee005791e06e1569a1dfdbbc08ea4e91c63129fad1728c498a8df25a6fff0d9e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hdef98feef36bf345a439dea0a76d0208b7d3c07bac3cfc6c0909973408f889c88cbb87e81f2794b6acfb57825b31729f6dcb6b11a3e0ea3e47bb2b647b5cac9d3e90605f9a941e672be1ba3e1e835acb3783607c521f59d169ffe49cc30120e3ea7bc48adcc21728e1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h88b3c5d250919d621e8267473c2536cf6f2cbb7291b0ede3cf63f5129db5e2034cdea080c655e70ed19ba9c4695a7e6b1a58296272ce9811196fa5252197d314f29ba7d0492cd0371e1d771089b7b8b0bda81c99bd6509693610cb0cbd75dff1cd377a738ed3b177d2;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h982fb333985e6d02d6a2adbbc53990a6591f568a217905d7ab0f7f88c67f16cb5d4abc93f7f8fe8ce829f38f302007fa50ff926413d03237460971b55235a5f1afde891d486e9d785207b1c83429f042c8bf4ca9332989c7894855d9b5d637c190fbc2a4256afebaa5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h13816af399b485625302d63bb4a07026f424ee33b9ff3a7a9766babda9aeb94a4927ceab9bee6d1e4c7619cf8c7825607790ca5b94da9439c93bbbd78abcb8417c535d26acf39bd94f3e145abf404d9f4437e54d99d6a3338e569708b8d9c523648f39147a9870fe6b8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1273205308efbc3afb6c6c3bfc6d62365961e002c70fc0c7cc07548fa70142a873aded8cfc1a37d1f8c7724d16748f34cd80be39d1ce062fd42a68f0318f847129231f91ee601c5e94937bea7356c8ab5045b5bf2a09e9168946a1da0ec1c6ebd0e62c5f2a132abba2f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc0ea58f9e435cb861164f1295280bc38a68ec6b6684340349fa8aff5afba500b87ce1ebdc9b77c16b78ba12fe8cd08cc8724f7c363ab1718dd0d3fdba2e8decee03ef1eb0bd76320e3e67c5cc273a9588829f7072e1c5c72f31010f79ebc7f5512863aa9bf0e0cf3f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f15281b1eb398b5941611be862fe91618fd0bed78afa0e2fa9deaeb1245fa77d103c1e2710927cd848e940f850855f4ab067c65613ab8f3a6703287025af371c9167ef230cd1b53b693ea7ac627d1e91fed213b165fe682940207bcdf5345a90d79aa373f705e7b41d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2c9bedca173e2dac0d21baaeb3c141886bdbbba70450ce6a1614179f3bb5b892ab6c8e94f110887553114d6982a1cd155d573733e4b3a6aebffa905d8808194677946a0b3c9b87bdd752ea0bdb552882862123047e16371d20623fa60f7f974e1d63418b2c429853ec;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h125f3195cb54ea59af026b32ac9d246b8873b8975a8a8213df4e3c7f260c887463e4579873e818316ae12da20582c68c90b9bbf350de5ee4935cc1fbfac7aff30a7d2c06512ddef0bcbacb98c1f63fc82da4099000fcc114cfce58b901f759094d53e99214adff79ca9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb13610ef00e811d4011378cf9f6e4fdd66f61a7b1b0689319d1424b8e58cc7cdab6b5de385d8e8e40e59cbf10a77e921be612b15feb97e55ce51d74b4f935f4d1872dcfe858f04edba446b899e98e1ea0b09e52bc433298faf9447d32695d23c7ad2a7cedcb92e2629;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1486f8dc5198a2db933102671da1d23137e11090b4fa3a6db80c6b663f1ed056ac40050e690f07200fc69d1efab41cf531761c50c1e579d771852451d00babaa104a3a16e749b9fd69c6f3fa3f61a87f6b1c1910e4d2ddcf3154555ffb14ac7daa39f4e26db165943e7;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a0284f8039bf2505e2e3a225af8241b3fce98fb748411c0068c94acac7c5b8d2283a07308685865c381d0fe1a89f05e84a0a75124a208d49a71f645c622bc2c03b113aecbfac4e403ed3e6915f982c3ab678deac2dc7ebd958685f96edf31bc48d19e4d08fa2936f04;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16899e8a8ef8874d33bfde71f38ceac40aabe00b3bd30f42c8b29ee9983cddb42935cbd9a41c996f733a2c9de1b14e783fb8b6129c35f26dd56e3586869d619e54c11227029ec9735d88e6bef95fd1a479f4da3089b9d05e6ea79893cbe1a85b06f8485dc3e33352cbe;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b0a67db83671a6059e853b74061a2fd7ff3915f96541802264862ba099d48167e5df95b7cbdbd868a6b7fb5a038158f53983d33b8d343ac301343f787df569363caf54781c412eb8086213710ba17d150fbdd08fcc59c413d7b734ad9175a695b9b756bb7b725027c0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hea59ddf0b460d9a3d51c2185523914e2fbd3f10f8372060e0e5e65c1c6340164354c01f88844e7b4193b37849a5fda717ad053f5d060f7067f6d9880a3c3afba2db3ebd25e7cdcf6887f1ac57791c6b2df4d7bc6469f5ff5f1dd4559535dd71bc0761e793e4860dccd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1681d24ccb24ae76d5d7a073418eab6588154217ca64df45b115aef7275ee99f1edd0b36d3901d65ac94d47b6b3d74fd266e2f7cfdd0f9397c2c9d4b4fe251f445d516292bd8bbe24281b50b38c8d651fafc9cfc3ddd3f08e4cc07a5c5d44237959e0c6149d93cfd7a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1c1793f5f99afd0a3bf34558550b7acbb577d0d89109c03add77823fc45c938955bd192cb5f5941dcf0b1e9d78d4abf8e287d84ac26ae0af09a777ca76b39da37cf16908fda7a9bbcf70e66392f95e904f3bad8f8050001c1c2c5ccc9f1e3da5444c9ffc32744e3b5b3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10a2554b5626e9f77ecdec1400a78eef4dfabe44e673f5abc6aa848571f1df832a62d17d23c0e3e95ac0da2b2f538178363abe16a9942d7e28d17a0667145c79518ec7ccb5b30979e0854f47a879aeec91e8f69310faf97b4e27d776f46d155bc927820192b5a3f7e79;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f222019437de8d8bb12db65ab780128389e3112bdaee3c328dece11c3f2742b48d2c6da712bb80661565ea3231131b300d280b1e19721484c84291121ee6ce513acaee939641551107cc9b965c4013bf484c22e073df2d6c4b5acea8b4e373355403345c8dd2b62e4a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16a86177b413a671b53afbe9dc5f3765548abb6bf28edbee4c030405673c60d4a01e740ebea97049d482deaaf4e4ae44851b499cb13829bb4bef5b0db4bf45cd4b94c6e0852efa765fbb97b41a9bc185e6c28d59e02443e80a01e4f59503349e703a2aa75d60be8461c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbc8fe7f950f9c5a8a24698af822b0f736c8aa10ec7c3d06161740a8c3accb998296d71d87dd57534f95f9db83817faa9d7a18b3c46e9688033d31d8edfae0cf9d787a7d8adc878e8d6332f4351dd22538b39e5b5a45ed374c0205a18ae2fe863ed7fa8da3b30ba26dd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h182641e54c83dc46463786fca2de3263bc67ec6bc2e4f46e511a34f12d7062adf636b288f9a619e859068b56ef0db763f4eda605d42c274d29952bad48886a623c5e5cefa039e4cd0960ae6a72faa6d30d3855a33e200e1d042d0d7f1c76eec6b43b32c23c58da5ee53;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f91c300932bce58e0c894bae062d41ef135ce89acededc0ea4f607ffc25a213e3626d9a3e8443ad088275f0b364b3a570bb521162451cf46483bce83bf9d6b724fc13b649ed9e56a7fb4f01ad49e46a494cbb2814af5ed00695abc11a6f67909c6c87802e28107f114;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbab200eef43d4f97567a1f5920227a94cbdab08ae4c4c690334a0f857fb1bb5e286c5424a0ea700f2042392e64ccb9dd0ba36d565a9245a1515d17f3fcac6a9084ed73e6f4772bd6f54f31d048451e88cb91cc481f0b2baefc5ab31d66e85668e12cba62a06954b09d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb7e46dd9d7ca726f3bc90be33e5390cf14baf59f77d92f768b7ad297af5e9e580aaa48d69fa12fee9bfa9ba9b303dc709331e2717ccf4e527ab7d87ae04901c0bbdf556eb62d75e396d38e972bb53074ac06c82fa898e890fde1a06e2ad61b6c383097daa0ae66bd8b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1005b9d2f4bfffa596f21ee56a3e2cf2bd9bb729173cf8d4793e4416ddb5e6d3f606b47ae2b390434195c0daa0df8c600d01686173518a7d15aba77ff4bd765a13082d38d91d7c1eb8c325dfdac0cc4026279cb92c69b51055f58beea879c93f1175149ba6827ae686e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hccf037f2039631e81ad9209928f24eddc83f45a1601f4539fa2504d1238a04f91ce8b5039a5ac7601728075b1dc197c76a2568febd9cf91e2cd4e41207bd1d70bb2b6be17627a6ad113aec303fbf9e8e8cdcdb334a8a40d413ced38812cf0f1cb158e73e64e86a0b22;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1cfbb3813fcfbeb82a478e7896519fee6d6c66c701e93509797b28b59b5d5eb95c901693e4de381417dd9a1a6b69ead140a146592c70102f6ba5fbfc589f1029335ba13aa06f32967433b7cd721d2b43cf2532222cf225c679a4987bab5a854120aaab28366419d25f9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1844374e99d4c6a7e98df839a46d81bf0584320307042dcb7735eeedc7d7dee50c08b88cb2edaa5921675a6d02ad7911ec0dcb016065c42f59133a0a32c486090655c600ceb260d0d711993263a0144c8f584cde4b9b353edc49997619841f56306ae0c153faf71a0a5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he9efaed3697ba5fa98007593b181caf849e9594d589b347ae4aabf5e65a36df1bcdbb13b4aeeb7531d412578ec202ab5493334d70d8c00d540719133566e4882c0c42052fcbf83489ddf5860b49c0f2c7f6330f75b885eebbc63df29b30a9aadfb4e446da07a56e876;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8457da1c48a460cb874107751a11cee290901caeaca113d6d0f9e96dc77013295468a2c3ce977e7d4bfb08996140c7d6a645459e3e22f6a3ee4b7059d70baea81c200d3371faefbf52da8ce71178dae002c5e6e79d0626c49906a4c67dfed4924c8d30e8bd39096a92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h2f91948e31f8c9484144bda5ebd208699bab31efb14bb6b25a70092a7c4dc97a4ca13c724c331a0f07031ac75c1d669f1b645e022e547a15d7bbd3c3192a20ad6d0e00ba836902b98ba8a6a34219390c2a97e1f24604c6e7bf1dbc821fb264b1bf2acdc1f64e013e4;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8c9367508d658bcedb1ff291197bae811626b452cda244777e733631e5f767ea8f9f88d1eff10393211c04729016c20e2b973006fb14d45142e39d7134019ee9d8992f2d2e256c7a910da82bb8f08c29bcbaff491c0dafd3206b40ab0e4f0ac780e5be20308680f89b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hfbda2e5e40dc125837b9ac6ee0f32069145ebb4af14f3407ee51f911092c0f3e00eb2eb882daa34d173243003555c1df431fa4b48e2bb36291d3b5b059b5682ffd0fd9321d716cab6d043878f8baa570b8dd3a466be58d8c1edd3a04335640238299b118ac0cae9099;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h16199cd33ced785786f9d0262a024dfef3c97da8ba9156a87f7bde46e3f24c70c899c4a955f8aca87f40222d467ae8f69aa98909c7b65081d79ada7049854d6085950ee9f4d813fe4fc27e27f4e0172026e1c88c6a10d9304284fb6425964dc88f372570908c4a5604c;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h14d980175276f21b83b075f84438538c4e748a607f94cad8e97ba106e9dfeee6bbc55a1f3574a73b68973c2d765070a91247c300dc109d6f567d24425264035e4e7e8cb342cca8b1126801307fd181229f670951d285c2628962b1372808b940939fe0f0916c20cdc85;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hb55a0e0b56dcdd2bc92d2eec3b2168d7493120d5408aa6a8a382a646bb62208ed45fc03c4fa74ec2a3df47bde9249a500f6dc2d00732ab6f48c4ff4ceca263a1edf6279bac9374a0481128b31fcce772293cfb795856e02bfe654ba613f0e49121db4a37c029b69f6d;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ea96643e625fb16d1a372d47ee1c228e77250c67a629c5b5f8d73e5cfd7111090f9fd735d3ca2e92cad1c5af719c66a8dfec286209e10904cdbbb67d2797f03d927e298ecdbcfd841d82240efc1f3f7287ffbe4ca987e6de39023f88c7076946eec64a4f72c9944552;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h105fc1f65794be0279130dda17ae0c28de502ff03e87d03bcef4ef3feb387e1d4eb688f7c0743138fdf82c64fcb07645ed313e5ecf3d0ba954d07310cc545cb5be9b9bedd40952616af165a1877794e2d8df127053a95f8339a091c6e31031e0656fa8fb31408c334e9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h633d4bd45312c0bb20a34e6b0a6d9c23b1dd2ac9a2f2653b576ff757fb277b02e057081296c0ebe0a77e419e6092c9ce423bbad581233114a3f54ae6dce783895f47466670245d5b68ed75d7b65a13729d43fbbc5deb0641744f1e4304c4ab28645b9be2df8576f9ba;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h183a210c1de64bad59a7035b303d2f27c31712e6780834b2bca41c97dc5f21313dcad78e49bb805500baa1f2eae4eacdeb917d5b45614e70c7bfcfe871d14179e14358f5a890ed247626468924bbf2211434e5321270095137d0701e64e0cb00ce414157dd6c03e134a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h180435be4012e06998b372d72d38f4012fc523d2a8b76e7eac2c86f0c3e1791897d07b3ddbb0a676dbc85c6ac18c20d7bbfb88ca7025f099872fa48af730128fcd81c5e7d777470b89b34e8d0029c56fb27324983c1fa1d46585b7d5cebb3cd22ccf7e2b9db5586afe3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3480b1d9d357564b3695c169dc986f5d9c8d4bf58b7765fbc60dd768b32add25ba9cd90e7d091c5a40e5781af8b57bf93fdffd94b713001dfb551419f66edf85d1a6750fbe5401e6490bb0e681f6357765730957250818a02cc08ac082516da6461ea00382899c7343;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h163e5f2d8d0c0ec0dd0b7a1f42953ae8e2773307224a8035befa6385df134efd5c4fcf53dd61df8a686be84935c6c14ba75902a533d09865020771a859ea8c00ef1715bd52f5ea3888d574e398b148b7a209f0c86cd4f2537601ff2e6dd37c1fd9c3f76d961f9a3223f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he098a5beaa953e3880556481a9c469ffb491938d71ace93673a5f312ac94e923426063fcaca78bcd6f7ee08347db83df434c6ac3cfd2560527fd72a5527ad915defbd417841c36a166ac599a4c46a896316022bb8c276e99313f3909c72c7e9ff01af136271a63160;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a6c867f86c159854ae36abcaaa69173653b522628cc60e692aa1e5de2b904cedae4491fa2f92ea94893b3280438e48fa2fc6f312e13bd92715df6dfa403ad387c543b7cdd889a62682cdfe614e9c4f6e79ed93b0c1f9ad555918346266316424f77b814ba113b34e4f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h17ca30c7fa8ad1dc294d54cd149697c73462cb839ed7ab6b2338afd1f5b86fd246f7d6eeca9b90fccbf849219d8ef367a4f7f1e23f81e505c4a236f12e2af6c329561428e1bcadb18c86eb31fc266f3c27cc766085dc55200a97c3e0ed1932a1b0f6995503454993457;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f3efacd4de95621990f405d7a6187ac9927f84fc8923a90f2868318ae4dba06e3b731b973c0e7eb67381c8154cb3b42045a5d9566bc84f1240bbc9ac0ca0d844305793b0fe89134a795c787732ca79da1c922981afda3f3da11614139165d9f353c86d99a5330eb191;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hd04d2e5450979e21b50e1ab521af6ae87dfa0a1c3204b7a99f5a15ab0d5dc42f144c0125f8c5ecdd51446cf94916db81a163138fb7836dc0b4981f376afed20ae589c13d3ac8dbfd2e62e504824d273292c83c76510070b415dfc12cb6605c5204ffc351264b067059;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h8cfc52500244bbca6992334457cb5650fac0fc8da7e0d4b5d8ce0c3e8c962ed53466a837f808d9ca7037a930a6947c715ed57908e2698b8bbbcb77a257a9138e97cc1054996e447f5c0e735329e28f0779bf62fa79dca8f15bc2d071c5416ca1bb4d249cac3bac517;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'he624e155acba006dd807851b2cc1c8c06c87c5044859c21babf188ec3c26081146e5958205f1ecd1bfbeaae345c7bc92fe97e439a1902b0c0d255fed14a30eeefa0db7debe4b3068fc3e65acd22b54dda88f5b4796d9cae3fae6a0d26599cf73013d10e9864cb4b61;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hc01f8282b0df4aac4b1a5df22d689e8c5917364c7ed50344148ce152c81149700d0a149a7671c996f02347c9f9c47b4f3ec61f549b5b6a126fd5049ac77d8db0a890570a05f91b68d4d565d8173ecd1a394bb5046edafe27bec69adbd371056674afdda4ecef298639;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h188bb3770c7685b33729277ecc89aea5d70172fa80f8cbdefdfcc928d3e5199f52a1151c9b101b6c2618b07629bf58d05743eb1d5481d9e7074133f8557b1e72f7d56db6313e7c01abcb241b40bcf568a6354ca09ce31b231adfb2aca1ef18928dbd7d199fd88a6b97b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hbdfb23b43429f39a2974a85e7bd8c09d5a4b6b7627370e2adbba896c333c1e0a23575ca709617230532b83d5467e9fb17635db1f9d507ebd101789732037ab4f2b4af5b0cb9835ca1775c881c47b5ad037a598ec58eee3e4302c3920727fd8576ed48488728b9cbcf3;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1af26d258a28bb9b04a8eb269ca035fca5b954fae4e518e2136b2591b0018dfb615c4e86b478789cb929e94c3832a55684cd9b2655ea76158912e4092431603794d88234f692899e4d08414ff81e084212f4e2030555b89858314056ab0b8d49542ecf844fd68d378fd;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h20893a2196b28e2dcc53ef89678d8b1cffbb681344a63158e1d06a083b78aad9ca9792e7f893420d9f6c92305c98fcaa066c9bd6544d416f9e76df97a383ef8bc86f425b913a11d75f476ee3af7878564e04411c3bea2e695d7dffa1fd323889e0d2dcfbb424d9e48f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1eb1a6b7dc3c77bce3c3a64c1e6221c4893ea74c28273cb7cb28e673677cb8ec0b4e456ffbebd7dc4e3298772f8099b22931514456d39640b9802169deb69beb572ee1f5a76e0ae697e8907962b00d04be647601f652b690c6a3c0a0312ec58fae2edaf7a4c3451df1f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e9a080a834b1e5ba4d0ffce1bb8a16d33a37982c3cedac8e58c20b0773a4efbe16bc940a794916eaac9697d6fd34ab8d8e526b99fb5b56f14f4721aaec8ad7c4f705757dcb608653dc48babc5b1e0400ad388e0bfdfc9b8c402193dcafa180b4ed2e191e17585f217f;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h4afab763cc00195c3f0e742b9d34ec9677805883a26f782cc728bb360b46fb81203e84b6ddd2197f3787bc604c601979f3eca0b6ab7c9554c478f0b1a56c332040db7fcc1f5fa70ef7bf599930cac198b9e532474b7eb5ddcb1a80f426b71df98a93d8a73ddba66a2a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1907a6db7e5164a5b7c96a4eb879212b9881940c52f5f4486a727ddfb772d1486c6d932b336726e37113aefb25a94685538f7395dbc71263e5bd87a977b62d38aea43d187f28392de8e61deb993105f5d5d607bee0b729b75fdbb99561e8e700eabfd001b592c2c668b;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1f4d18e28997037f1568a0eccce370ce8fc7c47603567b339204c848f44e30c716761e98e997f2ade6febd079bf9c663d189bd6183c9516d1a1014f38a57329528396e2a89bfc27531559f032a480b3a28db9f0335be64fb234e48d41266578fccf5e67ac21dc874763;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1e1e50d31e808f602254a0627f7fea04a4618ec70254c894b3868dcf216adfd399bf946c70e23ee47a072234ed450c9c56e9eee32e58c1938cd901d3b207581e97add6ad52d7138fca78e75383870e160839cb7dc595187db230263f795d41ec29cbd1fb97f004009d0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h550d1d02d008ecbaef4bcd7484ac0bd560937c26c1d4e13bd8b93946ff921f2f43cfd678b0e5868f6e981e1f1ff9054f1f5feea5ebb556855a33cb128189408d4f339044746110828d955a062f6aebaa40fc7e65c229ca159553acdcf704b0458be4662001e1e639d1;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h10abe73dc67b365031f54999445708a9e778078901cfffab705a8cb8319739d044e1080fd1280714d5e384ae0ac103db4ee9f16da7da94aeb85ef1c8575c371f5ab01eb43c24a4c85aa39fe8c351ef3cfcdb791b44a60dc7c786028b9d9a80fc2bdb9ebedbabadb3d6e;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'hf4e43e96d4d81b2c9f8545949c0c9308bcbcb9382d77203106ed4cbfb4c99899ed58b9f660fd607b39a2a3889a8c378eae7bde29663889f40a7b69077a72cd87ae89138fcd0115dd3686e3fce9576979c7b0fd7993d7c60e0afd1771280b76f1e5225e7e2376096465;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3cd31f4626dc2543f529f695e50821f14257b05cb8dc3525e98c35cb7e06b21de5e00c954d30eef6ba83c69611a113b9c4ec4e19782a4845e2bbffbf9ad8030a09298239cd91b9f4c07093d3b7938fc47a74a0aaa9bf096e384f868e2f1984d52dd0d0d4342458e6e8;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1a54355d4e0b438aa01e579207556f6e8de18e16e9fd35ede915d57ca32cadca0b355140813482574cf47d265aac0c3ef61b49c285b9a6a096a05a44e4347b49df5d7813598aceb9fb24735b7df9597798f2b47fbdadf5f1482a83dc3228c5676750386bba1f3de6a4a;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h3f87de6dd64ff26b3aba5e9bb91bec61860c52daf79a6959c527f10ab2a59612738418da75e82efc1afe64e04eb64bb88beea7bf8233c9fbd709319e50974f5fc1111a3c5907b008146cb71ff34f53885f2b6f4dc667de5ab8a29fd323824f5536894b1219366963f5;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h137ceaa4b540687eb61b2b5fe4e68c526ee9165495e7bdafc3b53a78f495223d099fd5c8a28751cf97e8c5a3c28f74b32432beefd8cc644c09b4333597f35c19e56ff44cc935a3bb50456138c4181b93f67cf674b3fc73c6c90eb9f184a0f8e80031fe4ff86f6068b92;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1417858bf7b9788c19e77ff52c1b2876ea17b5d010eb54b2ab4b188c33a31436c5a1e0335de48f4f7c85ac9f44cf6ef1e0beb4dbd20b14edfc2ae957300d6aee132c1a7eb5a9c3e75d317051d02cb1ed12a3ca1fd188aadb0c4b4951b1a8e9631c7f5feb10a122584b6;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1ada1c7e8740dce725980337e10e0510f0234b2843a6e73f5485a63431101554507c8fd240c8b4c99f68180b11f177e375398ed2b2de22ec308dbed8b777684efeff65e4b979fe66c82aeed45658530f57f78ffa73817fad9652a7901a4414b5f8f2e8aaf8e4674fe64;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h18a70d98b5019c4cb6856feabc3a9e35bb1015740cf2301ca16077da5a1da3a1ccb9008e0944a90dc4e4a1895a92f5c3f0666e63bb632ff34f804f9ff0c2d83ef307a7b63f4599470ddae2ee91ec643f49dc75710ca80baaf56aa05dad6d41fbf4df124059d388553af;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h981444a85a5425a002122a26ddf5400fcc3b9bb72e721b3357adc1f80755a0a22592084aaab476320244690b34495284e5b43259de71be771c8cc3a34726f73395ba4866f5804195b295777ffe1303e48bce725ba72ae7ac7ba5baee4e36c558e40284e20a550bbbed;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h98b567f5d18a86f3ee23b450d16a5cab7f0964c8e74f9616f2142f458e90be3076958129e94c9d7b3916357326f04a5b9baecf6476d3e17e85df0835739d9a371a120db22f5912d8c687d91a256e6f174c111677ed29648e33eca903331400390d0202693930d719d9;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h252785e7b4d708c00d3b2247676e7650feb334203844d659ca16d92e4acc9de98aa8f7f3b1e484315cb666e70ac53bd541120aafa424e31df95b83a1c10f75cc1ef4a7a1f7e8f732078b26e0a85dc3be7e583e8519d12fa1534f190a9c155b18602226ed4f9f2be8aa;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1b857311b0a6760cc18d69c1101323ae081bd8dafce8f13543b9bed40cbf7952282021557b4189ef22c6d5c64b4af7921a1b8f804b9dfd85d45ccfff04422d746761da2480e08552f8a2390898e6f8eefd21b6969e8d9e7bda1e8eda82ffdad21d7d6fdbc1395be4319;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h1008c0c4c6660b1eb04633d8326469cd59aafa3f8e91de4d2f7fd3508bcddeefac479664f2b31e73f11944e66dc670b32c3d554de7437d8ddea248d87c1d7c86a90c2d3297eb9f5ac1d84264866187f59dce19ad76d82d19620ad32cc36a5aa3acc6f02bce0bbe04fd0;
        #1
        {src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 841'h100a6694de6e10817b1131846e74f1137f422a123555c87543988b0dadd8a8b6e2ff79ccde1e61befc2bcc5e51787d5d5073e21b7d3fcbc38840cd151fdf78a8a41060e0d7b98c411646b143d577cfc5f5c2e801277fee4f458c433d331e4fc16b08beabc7e10f9d47b;
        #1
        $finish();
    end
endmodule
