module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    compressor_CLA128_12 compressor_CLA128_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA128_12(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [0:0] comp_out17;
    wire [1:0] comp_out18;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], 1'h0, comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [0:0] dst17,
      output wire [1:0] dst18);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [23:0] stage1_0;
   wire [40:0] stage1_1;
   wire [41:0] stage1_2;
   wire [57:0] stage1_3;
   wire [63:0] stage1_4;
   wire [61:0] stage1_5;
   wire [44:0] stage1_6;
   wire [43:0] stage1_7;
   wire [62:0] stage1_8;
   wire [63:0] stage1_9;
   wire [42:0] stage1_10;
   wire [43:0] stage1_11;
   wire [41:0] stage1_12;
   wire [20:0] stage1_13;
   wire [11:0] stage2_0;
   wire [8:0] stage2_1;
   wire [13:0] stage2_2;
   wire [20:0] stage2_3;
   wire [25:0] stage2_4;
   wire [22:0] stage2_5;
   wire [27:0] stage2_6;
   wire [21:0] stage2_7;
   wire [26:0] stage2_8;
   wire [24:0] stage2_9;
   wire [23:0] stage2_10;
   wire [19:0] stage2_11;
   wire [16:0] stage2_12;
   wire [15:0] stage2_13;
   wire [8:0] stage2_14;
   wire [3:0] stage2_15;
   wire [6:0] stage3_0;
   wire [4:0] stage3_1;
   wire [5:0] stage3_2;
   wire [5:0] stage3_3;
   wire [8:0] stage3_4;
   wire [11:0] stage3_5;
   wire [8:0] stage3_6;
   wire [11:0] stage3_7;
   wire [10:0] stage3_8;
   wire [7:0] stage3_9;
   wire [11:0] stage3_10;
   wire [10:0] stage3_11;
   wire [7:0] stage3_12;
   wire [5:0] stage3_13;
   wire [8:0] stage3_14;
   wire [7:0] stage3_15;
   wire [0:0] stage3_16;
   wire [6:0] stage4_0;
   wire [0:0] stage4_1;
   wire [6:0] stage4_2;
   wire [0:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [5:0] stage4_6;
   wire [2:0] stage4_7;
   wire [5:0] stage4_8;
   wire [4:0] stage4_9;
   wire [2:0] stage4_10;
   wire [3:0] stage4_11;
   wire [5:0] stage4_12;
   wire [2:0] stage4_13;
   wire [2:0] stage4_14;
   wire [4:0] stage4_15;
   wire [1:0] stage4_16;
   wire [0:0] stage4_17;
   wire [0:0] stage4_18;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [1:0] stage5_3;
   wire [1:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [0:0] stage5_17;
   wire [1:0] stage5_18;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49], stage0_0[50]},
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55], stage0_0[56]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc615_5 gpc21 (
      {stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_1[18]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc615_5 gpc22 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_1[19]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[5],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[6],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[7],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[8],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[9],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[10],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[11],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[12],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[13],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[14],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[15],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[16],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[17],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc615_5 gpc41 (
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127]},
      {stage0_3[111]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[18],stage1_4[41],stage1_3[41],stage1_2[41]}
   );
   gpc606_5 gpc42 (
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[1],stage1_5[19],stage1_4[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[2],stage1_5[20],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[3],stage1_5[21],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[4],stage1_5[22],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[5],stage1_5[23],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[6],stage1_5[24],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[7],stage1_5[25],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[8],stage1_5[26],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[9],stage1_5[27],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[10],stage1_5[28],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[11],stage1_5[29],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[12],stage1_5[30],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[13],stage1_5[31],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[14],stage1_5[32],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[15],stage1_5[33],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[16],stage1_5[34],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[17],stage1_5[35],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[18],stage1_5[36],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[19],stage1_5[37],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[20],stage1_5[38],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[20],stage1_7[20],stage1_6[21],stage1_5[39]}
   );
   gpc606_5 gpc63 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[21],stage1_7[21],stage1_6[22],stage1_5[40]}
   );
   gpc606_5 gpc64 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[22],stage1_7[22],stage1_6[23],stage1_5[41]}
   );
   gpc606_5 gpc65 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[23],stage1_7[23],stage1_6[24],stage1_5[42]}
   );
   gpc606_5 gpc66 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[24],stage1_7[24],stage1_6[25],stage1_5[43]}
   );
   gpc606_5 gpc67 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[25],stage1_7[25],stage1_6[26],stage1_5[44]}
   );
   gpc606_5 gpc68 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[26],stage1_7[26],stage1_6[27],stage1_5[45]}
   );
   gpc606_5 gpc69 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[27],stage1_7[27],stage1_6[28],stage1_5[46]}
   );
   gpc606_5 gpc70 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[28],stage1_7[28],stage1_6[29],stage1_5[47]}
   );
   gpc606_5 gpc71 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[29],stage1_7[29],stage1_6[30],stage1_5[48]}
   );
   gpc606_5 gpc72 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[30],stage1_7[30],stage1_6[31],stage1_5[49]}
   );
   gpc606_5 gpc73 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[31],stage1_7[31],stage1_6[32],stage1_5[50]}
   );
   gpc606_5 gpc74 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[32],stage1_7[32],stage1_6[33],stage1_5[51]}
   );
   gpc606_5 gpc75 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[33],stage1_7[33],stage1_6[34],stage1_5[52]}
   );
   gpc606_5 gpc76 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[34],stage1_7[34],stage1_6[35],stage1_5[53]}
   );
   gpc606_5 gpc77 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[35],stage1_7[35],stage1_6[36],stage1_5[54]}
   );
   gpc606_5 gpc78 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[36],stage1_7[36],stage1_6[37],stage1_5[55]}
   );
   gpc606_5 gpc79 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[37],stage1_7[37],stage1_6[38],stage1_5[56]}
   );
   gpc606_5 gpc80 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[38],stage1_7[38],stage1_6[39],stage1_5[57]}
   );
   gpc606_5 gpc81 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[39],stage1_7[39],stage1_6[40],stage1_5[58]}
   );
   gpc606_5 gpc82 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[40],stage1_7[40],stage1_6[41],stage1_5[59]}
   );
   gpc606_5 gpc83 (
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[21],stage1_8[41],stage1_7[41],stage1_6[42]}
   );
   gpc606_5 gpc84 (
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[1],stage1_9[22],stage1_8[42]}
   );
   gpc606_5 gpc85 (
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[2],stage1_9[23],stage1_8[43]}
   );
   gpc606_5 gpc86 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[3],stage1_9[24],stage1_8[44]}
   );
   gpc606_5 gpc87 (
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[4],stage1_9[25],stage1_8[45]}
   );
   gpc606_5 gpc88 (
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[5],stage1_9[26],stage1_8[46]}
   );
   gpc606_5 gpc89 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[6],stage1_9[27],stage1_8[47]}
   );
   gpc606_5 gpc90 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[7],stage1_9[28],stage1_8[48]}
   );
   gpc606_5 gpc91 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[8],stage1_9[29],stage1_8[49]}
   );
   gpc606_5 gpc92 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[9],stage1_9[30],stage1_8[50]}
   );
   gpc606_5 gpc93 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[10],stage1_9[31],stage1_8[51]}
   );
   gpc606_5 gpc94 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[11],stage1_9[32],stage1_8[52]}
   );
   gpc606_5 gpc95 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[12],stage1_9[33],stage1_8[53]}
   );
   gpc606_5 gpc96 (
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[13],stage1_9[34],stage1_8[54]}
   );
   gpc606_5 gpc97 (
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[14],stage1_9[35],stage1_8[55]}
   );
   gpc606_5 gpc98 (
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[15],stage1_9[36],stage1_8[56]}
   );
   gpc606_5 gpc99 (
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[16],stage1_9[37],stage1_8[57]}
   );
   gpc606_5 gpc100 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[17],stage1_9[38],stage1_8[58]}
   );
   gpc615_5 gpc101 (
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112]},
      {stage0_9[0]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[18],stage1_9[39],stage1_8[59]}
   );
   gpc615_5 gpc102 (
      {stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_9[1]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[19],stage1_9[40],stage1_8[60]}
   );
   gpc615_5 gpc103 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122]},
      {stage0_9[2]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[20],stage1_9[41],stage1_8[61]}
   );
   gpc615_5 gpc104 (
      {stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_9[3]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[21],stage1_9[42],stage1_8[62]}
   );
   gpc606_5 gpc105 (
      {stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[21],stage1_11[21],stage1_10[22],stage1_9[43]}
   );
   gpc606_5 gpc106 (
      {stage0_9[10], stage0_9[11], stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[22],stage1_11[22],stage1_10[23],stage1_9[44]}
   );
   gpc606_5 gpc107 (
      {stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[23],stage1_11[23],stage1_10[24],stage1_9[45]}
   );
   gpc606_5 gpc108 (
      {stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[24],stage1_11[24],stage1_10[25],stage1_9[46]}
   );
   gpc606_5 gpc109 (
      {stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[25],stage1_11[25],stage1_10[26],stage1_9[47]}
   );
   gpc606_5 gpc110 (
      {stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[26],stage1_11[26],stage1_10[27],stage1_9[48]}
   );
   gpc606_5 gpc111 (
      {stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[27],stage1_11[27],stage1_10[28],stage1_9[49]}
   );
   gpc606_5 gpc112 (
      {stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[28],stage1_11[28],stage1_10[29],stage1_9[50]}
   );
   gpc606_5 gpc113 (
      {stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[29],stage1_11[29],stage1_10[30],stage1_9[51]}
   );
   gpc606_5 gpc114 (
      {stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[30],stage1_11[30],stage1_10[31],stage1_9[52]}
   );
   gpc606_5 gpc115 (
      {stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[31],stage1_11[31],stage1_10[32],stage1_9[53]}
   );
   gpc606_5 gpc116 (
      {stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[32],stage1_11[32],stage1_10[33],stage1_9[54]}
   );
   gpc606_5 gpc117 (
      {stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[33],stage1_11[33],stage1_10[34],stage1_9[55]}
   );
   gpc606_5 gpc118 (
      {stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[34],stage1_11[34],stage1_10[35],stage1_9[56]}
   );
   gpc606_5 gpc119 (
      {stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[35],stage1_11[35],stage1_10[36],stage1_9[57]}
   );
   gpc606_5 gpc120 (
      {stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[36],stage1_11[36],stage1_10[37],stage1_9[58]}
   );
   gpc606_5 gpc121 (
      {stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[37],stage1_11[37],stage1_10[38],stage1_9[59]}
   );
   gpc606_5 gpc122 (
      {stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[38],stage1_11[38],stage1_10[39],stage1_9[60]}
   );
   gpc606_5 gpc123 (
      {stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[39],stage1_11[39],stage1_10[40],stage1_9[61]}
   );
   gpc615_5 gpc124 (
      {stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122]},
      {stage0_10[126]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[40],stage1_11[40],stage1_10[41],stage1_9[62]}
   );
   gpc615_5 gpc125 (
      {stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127]},
      {stage0_10[127]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[41],stage1_11[41],stage1_10[42],stage1_9[63]}
   );
   gpc1_1 gpc126 (
      {stage0_0[127]},
      {stage1_0[23]}
   );
   gpc1_1 gpc127 (
      {stage0_3[112]},
      {stage1_3[42]}
   );
   gpc1_1 gpc128 (
      {stage0_3[113]},
      {stage1_3[43]}
   );
   gpc1_1 gpc129 (
      {stage0_3[114]},
      {stage1_3[44]}
   );
   gpc1_1 gpc130 (
      {stage0_3[115]},
      {stage1_3[45]}
   );
   gpc1_1 gpc131 (
      {stage0_3[116]},
      {stage1_3[46]}
   );
   gpc1_1 gpc132 (
      {stage0_3[117]},
      {stage1_3[47]}
   );
   gpc1_1 gpc133 (
      {stage0_3[118]},
      {stage1_3[48]}
   );
   gpc1_1 gpc134 (
      {stage0_3[119]},
      {stage1_3[49]}
   );
   gpc1_1 gpc135 (
      {stage0_3[120]},
      {stage1_3[50]}
   );
   gpc1_1 gpc136 (
      {stage0_3[121]},
      {stage1_3[51]}
   );
   gpc1_1 gpc137 (
      {stage0_3[122]},
      {stage1_3[52]}
   );
   gpc1_1 gpc138 (
      {stage0_3[123]},
      {stage1_3[53]}
   );
   gpc1_1 gpc139 (
      {stage0_3[124]},
      {stage1_3[54]}
   );
   gpc1_1 gpc140 (
      {stage0_3[125]},
      {stage1_3[55]}
   );
   gpc1_1 gpc141 (
      {stage0_3[126]},
      {stage1_3[56]}
   );
   gpc1_1 gpc142 (
      {stage0_3[127]},
      {stage1_3[57]}
   );
   gpc1_1 gpc143 (
      {stage0_4[126]},
      {stage1_4[62]}
   );
   gpc1_1 gpc144 (
      {stage0_4[127]},
      {stage1_4[63]}
   );
   gpc1_1 gpc145 (
      {stage0_5[126]},
      {stage1_5[60]}
   );
   gpc1_1 gpc146 (
      {stage0_5[127]},
      {stage1_5[61]}
   );
   gpc1_1 gpc147 (
      {stage0_6[126]},
      {stage1_6[43]}
   );
   gpc1_1 gpc148 (
      {stage0_6[127]},
      {stage1_6[44]}
   );
   gpc1_1 gpc149 (
      {stage0_7[126]},
      {stage1_7[42]}
   );
   gpc1_1 gpc150 (
      {stage0_7[127]},
      {stage1_7[43]}
   );
   gpc1_1 gpc151 (
      {stage0_11[126]},
      {stage1_11[42]}
   );
   gpc1_1 gpc152 (
      {stage0_11[127]},
      {stage1_11[43]}
   );
   gpc2135_5 gpc153 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc154 (
      {stage1_0[5], stage1_0[6], stage1_0[7]},
      {stage1_1[3], stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[1]},
      {stage1_3[2]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc155 (
      {stage1_0[8], stage1_0[9], stage1_0[10]},
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13], stage1_1[14]},
      {stage1_2[2]},
      {stage1_3[3]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc156 (
      {stage1_0[11], stage1_0[12], stage1_0[13]},
      {stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19], stage1_1[20]},
      {stage1_2[3]},
      {stage1_3[4]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc157 (
      {stage1_0[14], stage1_0[15], stage1_0[16]},
      {stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25], stage1_1[26]},
      {stage1_2[4]},
      {stage1_3[5]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc158 (
      {stage1_1[27], stage1_1[28], stage1_1[29], stage1_1[30], stage1_1[31], stage1_1[32]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[0],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc159 (
      {stage1_1[33], stage1_1[34], stage1_1[35], stage1_1[36], stage1_1[37], stage1_1[38]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[1],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc160 (
      {stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[2],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc161 (
      {stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[3],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc615_5 gpc162 (
      {stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage1_3[18]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[4],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc163 (
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26]},
      {stage1_3[19]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[5],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc164 (
      {stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31]},
      {stage1_3[20]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[6],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc165 (
      {stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36]},
      {stage1_3[21]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[7],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc166 (
      {stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_3[22]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[8],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc167 (
      {stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_4[42]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[7],stage2_5[9],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc168 (
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32]},
      {stage1_4[43]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[8],stage2_5[10],stage2_4[15],stage2_3[15]}
   );
   gpc615_5 gpc169 (
      {stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage1_4[44]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[9],stage2_5[11],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc170 (
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42]},
      {stage1_4[45]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[10],stage2_5[12],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc171 (
      {stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage1_4[46]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[11],stage2_5[13],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc172 (
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52]},
      {stage1_4[47]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[12],stage2_5[14],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc173 (
      {stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57]},
      {stage1_4[48]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[13],stage2_5[15],stage2_4[20],stage2_3[20]}
   );
   gpc606_5 gpc174 (
      {stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[7],stage2_6[14],stage2_5[16],stage2_4[21]}
   );
   gpc606_5 gpc175 (
      {stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59], stage1_4[60]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[8],stage2_6[15],stage2_5[17],stage2_4[22]}
   );
   gpc606_5 gpc176 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[2],stage2_7[9],stage2_6[16],stage2_5[18]}
   );
   gpc606_5 gpc177 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[3],stage2_7[10],stage2_6[17],stage2_5[19]}
   );
   gpc606_5 gpc178 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[4],stage2_7[11],stage2_6[18],stage2_5[20]}
   );
   gpc615_5 gpc179 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[18]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[3],stage2_8[5],stage2_7[12],stage2_6[19]}
   );
   gpc615_5 gpc180 (
      {stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21]},
      {stage1_7[19]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[4],stage2_8[6],stage2_7[13],stage2_6[20]}
   );
   gpc615_5 gpc181 (
      {stage1_6[22], stage1_6[23], stage1_6[24], stage1_6[25], stage1_6[26]},
      {stage1_7[20]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[5],stage2_8[7],stage2_7[14],stage2_6[21]}
   );
   gpc615_5 gpc182 (
      {stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30], stage1_6[31]},
      {stage1_7[21]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[6],stage2_8[8],stage2_7[15],stage2_6[22]}
   );
   gpc615_5 gpc183 (
      {stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage1_7[22]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[7],stage2_8[9],stage2_7[16],stage2_6[23]}
   );
   gpc615_5 gpc184 (
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_7[23]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[8],stage2_8[10],stage2_7[17],stage2_6[24]}
   );
   gpc615_5 gpc185 (
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28]},
      {stage1_8[36]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[6],stage2_9[9],stage2_8[11],stage2_7[18]}
   );
   gpc615_5 gpc186 (
      {stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[37]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[7],stage2_9[10],stage2_8[12],stage2_7[19]}
   );
   gpc615_5 gpc187 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38]},
      {stage1_8[38]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[8],stage2_9[11],stage2_8[13],stage2_7[20]}
   );
   gpc615_5 gpc188 (
      {stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42], stage1_7[43]},
      {stage1_8[39]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[9],stage2_9[12],stage2_8[14],stage2_7[21]}
   );
   gpc1163_5 gpc189 (
      {stage1_8[40], stage1_8[41], stage1_8[42]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage1_10[0]},
      {stage1_11[0]},
      {stage2_12[0],stage2_11[4],stage2_10[10],stage2_9[13],stage2_8[15]}
   );
   gpc606_5 gpc190 (
      {stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48]},
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage2_12[1],stage2_11[5],stage2_10[11],stage2_9[14],stage2_8[16]}
   );
   gpc615_5 gpc191 (
      {stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage1_9[30]},
      {stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11], stage1_10[12]},
      {stage2_12[2],stage2_11[6],stage2_10[12],stage2_9[15],stage2_8[17]}
   );
   gpc2135_5 gpc192 (
      {stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_10[13], stage1_10[14], stage1_10[15]},
      {stage1_11[1]},
      {stage1_12[0], stage1_12[1]},
      {stage2_13[0],stage2_12[3],stage2_11[7],stage2_10[13],stage2_9[16]}
   );
   gpc606_5 gpc193 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6], stage1_11[7]},
      {stage2_13[1],stage2_12[4],stage2_11[8],stage2_10[14],stage2_9[17]}
   );
   gpc606_5 gpc194 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12], stage1_11[13]},
      {stage2_13[2],stage2_12[5],stage2_11[9],stage2_10[15],stage2_9[18]}
   );
   gpc606_5 gpc195 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18], stage1_11[19]},
      {stage2_13[3],stage2_12[6],stage2_11[10],stage2_10[16],stage2_9[19]}
   );
   gpc606_5 gpc196 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25]},
      {stage2_13[4],stage2_12[7],stage2_11[11],stage2_10[17],stage2_9[20]}
   );
   gpc606_5 gpc197 (
      {stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21]},
      {stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5], stage1_12[6], stage1_12[7]},
      {stage2_14[0],stage2_13[5],stage2_12[8],stage2_11[12],stage2_10[18]}
   );
   gpc615_5 gpc198 (
      {stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25], stage1_10[26]},
      {stage1_11[26]},
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage2_14[1],stage2_13[6],stage2_12[9],stage2_11[13],stage2_10[19]}
   );
   gpc615_5 gpc199 (
      {stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30], stage1_10[31]},
      {stage1_11[27]},
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage2_14[2],stage2_13[7],stage2_12[10],stage2_11[14],stage2_10[20]}
   );
   gpc615_5 gpc200 (
      {stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35], stage1_10[36]},
      {stage1_11[28]},
      {stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23], stage1_12[24], stage1_12[25]},
      {stage2_14[3],stage2_13[8],stage2_12[11],stage2_11[15],stage2_10[21]}
   );
   gpc615_5 gpc201 (
      {stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_11[29]},
      {stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29], stage1_12[30], stage1_12[31]},
      {stage2_14[4],stage2_13[9],stage2_12[12],stage2_11[16],stage2_10[22]}
   );
   gpc615_5 gpc202 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[32]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[5],stage2_13[10],stage2_12[13],stage2_11[17]}
   );
   gpc615_5 gpc203 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[33]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[6],stage2_13[11],stage2_12[14],stage2_11[18]}
   );
   gpc615_5 gpc204 (
      {stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43], 1'b0},
      {stage1_12[34]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[7],stage2_13[12],stage2_12[15],stage2_11[19]}
   );
   gpc117_4 gpc205 (
      {stage1_12[35], stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_13[18]},
      {1'b0},
      {stage2_15[3],stage2_14[8],stage2_13[13],stage2_12[16]}
   );
   gpc1_1 gpc206 (
      {stage1_0[17]},
      {stage2_0[5]}
   );
   gpc1_1 gpc207 (
      {stage1_0[18]},
      {stage2_0[6]}
   );
   gpc1_1 gpc208 (
      {stage1_0[19]},
      {stage2_0[7]}
   );
   gpc1_1 gpc209 (
      {stage1_0[20]},
      {stage2_0[8]}
   );
   gpc1_1 gpc210 (
      {stage1_0[21]},
      {stage2_0[9]}
   );
   gpc1_1 gpc211 (
      {stage1_0[22]},
      {stage2_0[10]}
   );
   gpc1_1 gpc212 (
      {stage1_0[23]},
      {stage2_0[11]}
   );
   gpc1_1 gpc213 (
      {stage1_1[39]},
      {stage2_1[7]}
   );
   gpc1_1 gpc214 (
      {stage1_1[40]},
      {stage2_1[8]}
   );
   gpc1_1 gpc215 (
      {stage1_4[61]},
      {stage2_4[23]}
   );
   gpc1_1 gpc216 (
      {stage1_4[62]},
      {stage2_4[24]}
   );
   gpc1_1 gpc217 (
      {stage1_4[63]},
      {stage2_4[25]}
   );
   gpc1_1 gpc218 (
      {stage1_5[60]},
      {stage2_5[21]}
   );
   gpc1_1 gpc219 (
      {stage1_5[61]},
      {stage2_5[22]}
   );
   gpc1_1 gpc220 (
      {stage1_6[42]},
      {stage2_6[25]}
   );
   gpc1_1 gpc221 (
      {stage1_6[43]},
      {stage2_6[26]}
   );
   gpc1_1 gpc222 (
      {stage1_6[44]},
      {stage2_6[27]}
   );
   gpc1_1 gpc223 (
      {stage1_8[54]},
      {stage2_8[18]}
   );
   gpc1_1 gpc224 (
      {stage1_8[55]},
      {stage2_8[19]}
   );
   gpc1_1 gpc225 (
      {stage1_8[56]},
      {stage2_8[20]}
   );
   gpc1_1 gpc226 (
      {stage1_8[57]},
      {stage2_8[21]}
   );
   gpc1_1 gpc227 (
      {stage1_8[58]},
      {stage2_8[22]}
   );
   gpc1_1 gpc228 (
      {stage1_8[59]},
      {stage2_8[23]}
   );
   gpc1_1 gpc229 (
      {stage1_8[60]},
      {stage2_8[24]}
   );
   gpc1_1 gpc230 (
      {stage1_8[61]},
      {stage2_8[25]}
   );
   gpc1_1 gpc231 (
      {stage1_8[62]},
      {stage2_8[26]}
   );
   gpc1_1 gpc232 (
      {stage1_9[60]},
      {stage2_9[21]}
   );
   gpc1_1 gpc233 (
      {stage1_9[61]},
      {stage2_9[22]}
   );
   gpc1_1 gpc234 (
      {stage1_9[62]},
      {stage2_9[23]}
   );
   gpc1_1 gpc235 (
      {stage1_9[63]},
      {stage2_9[24]}
   );
   gpc1_1 gpc236 (
      {stage1_10[42]},
      {stage2_10[23]}
   );
   gpc1_1 gpc237 (
      {stage1_13[19]},
      {stage2_13[14]}
   );
   gpc1_1 gpc238 (
      {stage1_13[20]},
      {stage2_13[15]}
   );
   gpc606_5 gpc239 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc240 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc615_5 gpc241 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[6]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc615_5 gpc242 (
      {stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage2_4[6]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[3],stage3_3[3]}
   );
   gpc615_5 gpc243 (
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16]},
      {stage2_4[7]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[3],stage3_4[4],stage3_3[4]}
   );
   gpc615_5 gpc244 (
      {stage2_3[17], stage2_3[18], stage2_3[19], stage2_3[20], 1'b0},
      {stage2_4[8]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[4],stage3_4[5],stage3_3[5]}
   );
   gpc606_5 gpc245 (
      {stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[4],stage3_5[5],stage3_4[6]}
   );
   gpc606_5 gpc246 (
      {stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[5],stage3_5[6],stage3_4[7]}
   );
   gpc615_5 gpc247 (
      {stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_5[18]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[6],stage3_5[7],stage3_4[8]}
   );
   gpc615_5 gpc248 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[3],stage3_7[6],stage3_6[7]}
   );
   gpc615_5 gpc249 (
      {stage2_6[23], stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27]},
      {stage2_7[1]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[4],stage3_7[7],stage3_6[8]}
   );
   gpc615_5 gpc250 (
      {stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5], stage2_7[6]},
      {stage2_8[12]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[2],stage3_8[5],stage3_7[8]}
   );
   gpc615_5 gpc251 (
      {stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage2_8[13]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[3],stage3_9[3],stage3_8[6],stage3_7[9]}
   );
   gpc615_5 gpc252 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16]},
      {stage2_8[14]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[4],stage3_9[4],stage3_8[7],stage3_7[10]}
   );
   gpc615_5 gpc253 (
      {stage2_7[17], stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21]},
      {stage2_8[15]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[5],stage3_9[5],stage3_8[8],stage3_7[11]}
   );
   gpc606_5 gpc254 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[6],stage3_9[6],stage3_8[9]}
   );
   gpc615_5 gpc255 (
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26]},
      {stage2_9[24]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[7],stage3_9[7],stage3_8[10]}
   );
   gpc615_5 gpc256 (
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16]},
      {stage2_11[0]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[0],stage3_12[2],stage3_11[6],stage3_10[8]}
   );
   gpc615_5 gpc257 (
      {stage2_10[17], stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21]},
      {stage2_11[1]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[1],stage3_12[3],stage3_11[7],stage3_10[9]}
   );
   gpc606_5 gpc258 (
      {stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5], stage2_11[6], stage2_11[7]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[2],stage3_13[2],stage3_12[4],stage3_11[8]}
   );
   gpc606_5 gpc259 (
      {stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[3],stage3_13[3],stage3_12[5],stage3_11[9]}
   );
   gpc606_5 gpc260 (
      {stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], 1'b0, 1'b0},
      {stage3_15[2],stage3_14[4],stage3_13[4],stage3_12[6],stage3_11[10]}
   );
   gpc606_5 gpc261 (
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], 1'b0},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[3],stage3_14[5],stage3_13[5],stage3_12[7]}
   );
   gpc1_1 gpc262 (
      {stage2_0[6]},
      {stage3_0[1]}
   );
   gpc1_1 gpc263 (
      {stage2_0[7]},
      {stage3_0[2]}
   );
   gpc1_1 gpc264 (
      {stage2_0[8]},
      {stage3_0[3]}
   );
   gpc1_1 gpc265 (
      {stage2_0[9]},
      {stage3_0[4]}
   );
   gpc1_1 gpc266 (
      {stage2_0[10]},
      {stage3_0[5]}
   );
   gpc1_1 gpc267 (
      {stage2_0[11]},
      {stage3_0[6]}
   );
   gpc1_1 gpc268 (
      {stage2_1[6]},
      {stage3_1[2]}
   );
   gpc1_1 gpc269 (
      {stage2_1[7]},
      {stage3_1[3]}
   );
   gpc1_1 gpc270 (
      {stage2_1[8]},
      {stage3_1[4]}
   );
   gpc1_1 gpc271 (
      {stage2_2[11]},
      {stage3_2[3]}
   );
   gpc1_1 gpc272 (
      {stage2_2[12]},
      {stage3_2[4]}
   );
   gpc1_1 gpc273 (
      {stage2_2[13]},
      {stage3_2[5]}
   );
   gpc1_1 gpc274 (
      {stage2_5[19]},
      {stage3_5[8]}
   );
   gpc1_1 gpc275 (
      {stage2_5[20]},
      {stage3_5[9]}
   );
   gpc1_1 gpc276 (
      {stage2_5[21]},
      {stage3_5[10]}
   );
   gpc1_1 gpc277 (
      {stage2_5[22]},
      {stage3_5[11]}
   );
   gpc1_1 gpc278 (
      {stage2_10[22]},
      {stage3_10[10]}
   );
   gpc1_1 gpc279 (
      {stage2_10[23]},
      {stage3_10[11]}
   );
   gpc1_1 gpc280 (
      {stage2_14[6]},
      {stage3_14[6]}
   );
   gpc1_1 gpc281 (
      {stage2_14[7]},
      {stage3_14[7]}
   );
   gpc1_1 gpc282 (
      {stage2_14[8]},
      {stage3_14[8]}
   );
   gpc1_1 gpc283 (
      {stage2_15[0]},
      {stage3_15[4]}
   );
   gpc1_1 gpc284 (
      {stage2_15[1]},
      {stage3_15[5]}
   );
   gpc1_1 gpc285 (
      {stage2_15[2]},
      {stage3_15[6]}
   );
   gpc1_1 gpc286 (
      {stage2_15[3]},
      {stage3_15[7]}
   );
   gpc606_5 gpc287 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], 1'b0},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc288 (
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1],stage4_4[1]}
   );
   gpc606_5 gpc289 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[1],stage4_5[2]}
   );
   gpc606_5 gpc290 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[2],stage4_6[2],stage4_5[3]}
   );
   gpc615_5 gpc291 (
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4]},
      {stage3_9[0]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[2],stage4_8[3]}
   );
   gpc615_5 gpc292 (
      {stage3_8[5], stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9]},
      {stage3_9[1]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[3],stage4_8[4]}
   );
   gpc606_5 gpc293 (
      {stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[4]}
   );
   gpc615_5 gpc294 (
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc295 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[2],stage4_12[4]}
   );
   gpc1163_5 gpc296 (
      {stage3_14[6], stage3_14[7], stage3_14[8]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage3_16[0]},
      {1'b0},
      {stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[2],stage4_14[2]}
   );
   gpc1_1 gpc297 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc298 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc299 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc300 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc301 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc302 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc303 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc304 (
      {stage3_2[0]},
      {stage4_2[1]}
   );
   gpc1_1 gpc305 (
      {stage3_2[1]},
      {stage4_2[2]}
   );
   gpc1_1 gpc306 (
      {stage3_2[2]},
      {stage4_2[3]}
   );
   gpc1_1 gpc307 (
      {stage3_2[3]},
      {stage4_2[4]}
   );
   gpc1_1 gpc308 (
      {stage3_2[4]},
      {stage4_2[5]}
   );
   gpc1_1 gpc309 (
      {stage3_2[5]},
      {stage4_2[6]}
   );
   gpc1_1 gpc310 (
      {stage3_4[6]},
      {stage4_4[2]}
   );
   gpc1_1 gpc311 (
      {stage3_4[7]},
      {stage4_4[3]}
   );
   gpc1_1 gpc312 (
      {stage3_4[8]},
      {stage4_4[4]}
   );
   gpc1_1 gpc313 (
      {stage3_6[6]},
      {stage4_6[3]}
   );
   gpc1_1 gpc314 (
      {stage3_6[7]},
      {stage4_6[4]}
   );
   gpc1_1 gpc315 (
      {stage3_6[8]},
      {stage4_6[5]}
   );
   gpc1_1 gpc316 (
      {stage3_8[10]},
      {stage4_8[5]}
   );
   gpc1_1 gpc317 (
      {stage3_12[7]},
      {stage4_12[5]}
   );
   gpc1_1 gpc318 (
      {stage3_15[6]},
      {stage4_15[3]}
   );
   gpc1_1 gpc319 (
      {stage3_15[7]},
      {stage4_15[4]}
   );
   gpc606_5 gpc320 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc2135_5 gpc321 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4]},
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[0]},
      {stage4_7[0], stage4_7[1]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[1]}
   );
   gpc615_5 gpc322 (
      {stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[2]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc2135_5 gpc323 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[1],stage5_9[1]}
   );
   gpc1343_5 gpc324 (
      {stage4_11[1], stage4_11[2], stage4_11[3]},
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[1],stage5_11[1]}
   );
   gpc1163_5 gpc325 (
      {stage4_14[1], stage4_14[2], 1'b0},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], 1'b0},
      {stage4_16[0]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[1]}
   );
   gpc1_1 gpc326 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc327 (
      {stage4_1[0]},
      {stage5_1[1]}
   );
   gpc1_1 gpc328 (
      {stage4_2[6]},
      {stage5_2[1]}
   );
   gpc1_1 gpc329 (
      {stage4_3[0]},
      {stage5_3[1]}
   );
   gpc1_1 gpc330 (
      {stage4_5[3]},
      {stage5_5[1]}
   );
   gpc1_1 gpc331 (
      {stage4_16[1]},
      {stage5_16[1]}
   );
   gpc1_1 gpc332 (
      {stage4_18[0]},
      {stage5_18[1]}
   );
endmodule

module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [18:0] srcsum;
    wire [18:0] dstsum;
    wire test;
    compressor_CLA128_12 compressor_CLA128_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h26564ef418f8a67ee261dfc95b235f3eeb6ef82f1225d867d143583165678e7a41c4051f2415d5e3c723d2e8a5184b0969e830e2ae901398052a71a4874ebb3564e7e5bfef1c7b011e9abdd3b8d97aa39ff6967e7b8d62802cf633b4fe32ce0b541e9ade48f200b3781be8386bf3c317824ac739bba223d58a5b0c6bc9040ced7e70ed8f2c0d37bc53b4f13d1d82d12db380b9b5fbb4bdf861d3784ab8fb7089e8c0ca4b68d6806b36f78e73cfffec13c4e4a5e799861809df6e9782997d994;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hdfcd6b39574619f612a8e5dfaabad335a2507c24cc9c3d00326025ec34270ee3775aec3606509242f730696b3a724d27c027ea783815a2bbde9bc8794131cd7607c030cc4fa2aea25614627ec26804e74bd6a82bd0780595b99c593bd59d159b12bd0279c9879f740192f67a9555978e3a59f60c15e4dce62771bcc57441fdfa95d5fa0ff32807f2a8176cb6bfbae200a0a220cf682a0a303c9bdcb67a162249c395bcfa23aa21e1bc38df9b9c6e8b9b0836ff7e88ce0b227a9086f1d261ed2d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h6213bc4f3bd46ec57df7a54340b03ede1ad0af8620cc858e6c7685428630f9f2b8297a174a1cd65e580a0a191ab8ef3e3482fdc1b283ea0ccc14d69dee41c4224e83ca4f97e655c2465c0742f53b80ac14ac9c4768ac2747947b7693f737ef8422fbb589ce00f981c223a85cd06ab30e037ab8a1b4fea00b64b5c971c83b31338710488e1244e262f02355247583e144a13e97d13424fff97692950a4ee7e62430648e14a5ad7a589f04d6a057bf59f82926d020f384e9ee6069e742ef72fb30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h78cc6ada878ce28d9b1de2963cd5a14a11d4d0ba9c590e7fbb3966932acc82bb9f784128fd586e1e85b4d296ff1cef8bcfba13fd558156ea29eb7ada9f5abb82a9f832939c467e778df08b4644938af1eab3938e1a26af58fb2b0ba45d0ab8cc27cb1be74ceb3572165db62c1856da937df4ca59850cade7b5673618c4d827d39eabd70c7d5437920b8ef2479780184b5018f31cf47a4d5787263a89a95a77e2219ae32c1269330ac93ba11b4f2425127064d1cad22717d3ea35bb128c086b27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hbf2d33813635ac3de395da8bf6750c305b33c58e43834cb10f2b857fe293cd00f0d56aa1069981d2a3cbde40eb7bb2d50d90eee9a1b9ae638ea96607f8c207a7132a6641e995663807b9966c180f95951bb0e5dc32eb2f4e23b51d94069033ff401da86bd8f0607a7442265964d75c130dd40f8d44b423e3b44da10f0a509a515015453419036d779f4ed22c4905db57646f20999531c4e247a65ce0ba16549577d07b71c41d6b3a419269b65a51b6ef7fbc2c31c7b4360e656eef78c813c5a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he49b6b08e2e00ebd57f06a92e5c2bf7a56fe1883715bbc24aec50caa9679e3e3430308c83d139a61cbad17297364be9446dac94984d946140a696b32ad020444c264b7f0ed5b7416251fabd459c9589111c8f7f65ecc157d17f5ac3f4fb9a238d7978829506a7430469c94c24f412cd6ef0758bc32c19274f6f84d888d273e89c56ab3ff5a68ce56502870436c2de67c688f6258b357e9007a10e44aa2d8a6100d4f2e51074ecb7e1f06b77275a5fe67ecaf1d33b90a61a3a2ee23f9dbfb3f1f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h91bb56f4150084cf38c78fdba62e2d01b60ea091412e17024067f97dad4c28fbfc902d437b7713334d9f5e674ecdf38f7725f43dfbd1bf99f715db306a4237c38c4132670efaf2ed0dfbaa680b959cb5416e94cd600625e5e5cbd25edd2e446f2da248c84e7454ed2b939aa0211def1fb453ac9bbc16fb19da58dba12dc401780ae0e836e219cd553a547b6831cc929fecb84f196173e92f6cb6027bd04da4445b445909d1db1bdb26230a91f1f91f408542bd43e0af53f38ec7cc792b64b18f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc0145db91eae9c3f3b95ef8be9851bd656797e0ee1e88ef209bef63b06e102ad6a2cf66c970f7ca88dfa8a4baf046cbd075dbd989a6040b524ccf6ea6a6d39c490a7e44190d91d969a559eec751eb0291ddbc6a794072226f7c88b2cd07912fb11be0a3b3a3dbd565ad06bc7acec3ee6519d7e7ff5fdd18ab9acaf8e3454b5ea3a8a45f1bdfa11ff259809d722f84eb6227eccd0deb9c46a0cb93e6943d4055a35c4117acbb309d3f35971cdea61179992b7901fc56b5bed391ab621068ebe96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5776c82ed3fe338e9d31115d45b7a48f5d42308b35134310d75524351602a32db7a0d6e950473e1de50757fb38f3f76d5ef4de8dcf3d44c095256ae5bbd0f4d98a87dfb7bfeb3fa2ee5b8a8b59bc3b5de8d096808d9d110436f92725a7cc86aeb0f235380aa09e8bc52cddc75b57ada086d9fa2e4de6b613cd0535ebfe355bbd23685344aed0546676ecdaab1c3aa2c139cf38c3099b0ee3648a40891b23ff906acbde43839a50fdb9ccd1f6fc133b8a29af355cd3ebe3ae220e8701e766145b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd3535d2b167c86b8d58503517113f1d4a235884a39d4991402a61290ddaf3b5645ef1103e202e04113a29b415090d4390bc16b9f042fe07971b0d96613f2283e6ea83ef900e249c7fded9b5cb8ac3ea41edae266c07265c55f56db5ab0a82a6f7f6edc1d2287491fa67899d8c07987c31b49c2fe5970633f1cc9d831035bdae73e7033ff5b874344da2ebe31fcf121a0d015d62d844fc35342a0d7b4dde72ac7d7d5a802df2d7b0d464e81950298c9a60db1308018aa19121a7e36bf20cdd8e9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb31a522c11b6037a716901c8f3bda73c87ad9288a4b2270b1c34d1feec4e09dc45bf5b0987521b79a63303b96ad7844dcfc8c402a3f587be5e300c566a5d7edb2a55db6ae6c7d27814fb15b3038c9c4474525945061d1ffa64c114e2a3d856875a3e4522992254798507c37b1db1cb8b4409618c2358b109055324735302eb142a18852b618ba8bf2a8f66e3d413f6fec02f4706c1d97ae8725e56337a0a2572309d6af1ca0539822eaa345ce8f52f5ceb817f8b102447ae9d9e07e9661d0e48;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha3d06e9fc82853db4951fdb79f7e8d18b94be15ab1cc7a85909e38b220b7843f2433739fa3fab97bf2a692bc6bc64ed8102359f03e8570e4af4a4a7cbc85f2e846f421ac2ecaad75e71a020c05a43336ac456a762a48620f68730886b45d35b582eea006d730c617ae47cacd557aa3a704e8e21a0203baf9104ea39154024a9d10771cc155b8822f038f173efc7ae364faec480ac64e3577d02a28291562a0d6644cb26f2df18ceb7ba51797afb49740cbf80f6ce486a211ae2b3165645868ef;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hde374b05bf609778da3e8e36fd09dbebcf8666889887a140a2d19de2c2e113bf4df42720b2f97841c5d2ff5a6dfda1867bf206cfa898065efff27cbf32c5727de318bbec69240257c8242f4c686d6bc610bc9dac97f41d4bf7ae94ce34a0df38422169caddd72176f4682401e8c6a755ad15b9f82e49799b532298f22da2d7d5b8faba134cf367bfc49fde7505b0d99281a02dbc208e0a6385944a134a1b47880ef391a03e378de88183c74922333ef94c2b90992b879e7522d7091ead43f0ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8c73c3b566381dbc2a3e1430ea2e4b853889371f53254e1a102449006e82859ff914f961b0a468d40e6bd5fdb49ad5b5e22f7382845d5e170a03cb8ed70536a48cb4d400d8941c8fb0b1d366706fe7a21c4926eb3c29e356d0047543b8ada5e759bfdd23b96f93c5b07fb4434e80b52a50c351b33e4802b0164669ec1740e1fb265916303dc0abbbf710304dd1027e7d224b10ed7d2fd5b0f1ff6d67f6febac85a57bca2df701124f3ad5363dd8c3916a5460b031b51ed0fe571cbed77457ff3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc5511ba4a324ef03fd311664a39828d73aa44009f28fcafbaf80d9ff26e175cabcae59ac22ebb93607753b23daf5b4674dcb17dde13f0b161229d89a991626e95ff07417f5c54c9cbc518e5279ef8f8176ba608aae90367d0c332b53dc942e8bc39eb15588ea958c93c56e48d0c8709f31661702d986a49718afa89db46d0c239de1550a60753e7697d1c927f29a21e63a071ba1fc767d6dfe2321c8843ba8f848deba26d093892dc4e1c8dc83fa7ee42692cec26f241fefcb731fd1b25d994c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd390afc85463f3aa02c89010217d2358e299448de7e6b2bd98da7b2ebdaee2b9ba17583b57218a404d3ca3625f8dbd3293a6f671c6b6fefe8e3cfa6d731a918f0b5e0af4783f3cc3cbb28b574ba4445ec86419b6815e2b58e38a15199602207c4a220def16450c7a62727977b63830da18f2144ce1a6f3d9a40f497eb362858f38d7dfb6ad9b86ee4985ceaa0eeb7a068c2462808d51ea591b00c7be31d3b57277e1f7266c12cd7d7347b39a657d8dcada4ce3e9546b85a3b12a0b29a64c7261;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc93f5b43fbe843072e697877c0c205f8be295332ddb371ee7926b978d8814a1b09597950f8c1991d7ff0cae66a4807f808958618b8571ac99c7154c12890122da83652b71df35555c0921091826871888639a2703471e6c612909c46eff6c93491555d57eea5429f40b837cdb610159e0e1e1296b23d724da83af9108d39b74eeaff4f8ee1a27a068e7fbc84ef4e01a7595e8492c1373624fae00d338643660d635cac73388dfdab8955c60b90d16a73a4be347e371a0bbabba930ce3fb59bc3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hac334ac8dcbe410c3f51025ad83ff35e126b7b3e6c103a7cadc0acfbea4d41b4bd70448f20bc02a0d3629b5034aaaa1bc1084f9aa7dfd6f70ac389fcf5027e8b35bef9ac38be5a8b42c66e625476f7f9868a84050c733d27c1051f4c542a310a00a8110460bccce2fea7d3cb68756b22d43ce3401770ec06140787225e9b89ebc5310c6bbada8bce0f49cfeaf1367164477fc41ba04f9a6f343942ca42a03de6cb55ada17d64de38f5df886b6ec9a77746412c2244e1e0569fb9ae4b50e5a406;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h45aed494d510339f7a654dd7827502f4bf9afe95711597c7ab0201927f1662d36b582e78b1851dcc824ce9180049f9104c28004b144b367af05480ea6ecbebfdbdf623d1cbec201259219892402dcf4da08354ba08f1ba0e3261d7ebd33e09cb1b531447cbffb86b3f29ab36ddf088135e9e39f56501207faf40313f9120d82d168f4b7d21be31a96c95bb36d3767d7c62acb8b1f04a5a8baa77fa6202525207ebc9130011e825154d455a04078cfea2dc8583c9c829e24070c4b42c0d7055fd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc5dc7f97183b2f78a0d444a49ab2d5b5fb9aca8d6994d8439eac6b94bd5c10aa16e5a6aabe0293db0914c0c96e85beab75e279444d8925166870ba35933feb81af8649e08051ffda18609602c7c52b32c2497bd8ed819cee19d053427877005be4146c7d8549f7b5bbed80ec8a88d7ad9807f9c7ceaeb92101e4b83ed0e7f6ec5e76e6bd70abee7da629c4bccc0a51c1579c1b15f73b6bcc6f71df940184505cc695c78690ada6a7a6ae0fcd4ada886a4a9420f02cbd20c59ef4c2e8724762a7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hccb7dcfc7ec91791df177cb17eb9fc6558e16bc75ceeb016cd4d3ef2c41f319b4e7b41593a1aa374eba2f07780035cbf3788bb54b6c2085f45c8e30e069fb5cc9a261e5e295b56395ad6dc1a3eebe64dce57e95dd253b4446c3cf0ff8df1113855584bb29c30aff732c366c0dd113e4c22f1fe76e4e43c242a3fa5b2600f1f94a082c0b5bae06a8a03afae9c5a158b8919ef294e9f1c9dd64c07968ba059a67feeb549c254f4d66604a1bf9f02762bbbeda1654f475da76de8a5648bc76ba310;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h779d6894259e5ec2080ebf520e9af589929ba9f28b1a6dc49b7594aa6908d1e14c8d7b16c8ad881d70e163269f7e71aae9d278674e080e8aee5b2299e68f78b0d180e65592adfbe2d2fcb4c6028ba5424dcd4abcaee444b9823be2da5d4548fffb36a9b6cc3554e46608dc237ffca1fcffbfd167577631c0982919f8abd2f9baccc90b634462b5bfb6abbe75c0e0d77887052c43f25435c5ce57fd3f3ad51286dd5699da060a3b14bda59484d0189eae1d6ecb0718ec8c44eeb9b88b778f4c45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h22437e790292f776e1db8bc3592964b83bc2d12cc9c0c7f9cff9d36d639601978306b18e7df32d5cee771d347f23d0a5518c31d830338a853242019567017c19517d3c49618cb18e3dc17a8e67c087e4da557755e13df85421a2822bab555ff01127f9c461c80370d98547a521e0dfa5e279c033feb20bcf0e75212255ce8e7ea5daa928083f530b9161521b4a6e1d78f623ef48e349163c45ddc7d4378969cf9cb84582d05cff8ab36b098efa8315d6a7ae0c76b283ab9ee7b22584423ff7ea;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf173247dbf54446eb8f73c5bb4701ceffb449de9d4fd0ab70d189cd0c7f3431377573df9cd31d9c26ab58602976011def483be01c9b49c8b45b71942a39f6c3209bf6f040d646054d5b5991c03fd0f48c030d9dbdfd324e5f8b91d6838096a0c046130af4ccadee36e4a76250b4e65f218c38690e36aebb91f4862ad9444f592c238c0221dde46733910d8b38268e696fde8016af4aabd631d2c16a259687b7fcb8104115cba93d15248361ad8b0183776f950c6f44688af27b6f9e8d9540aae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf53b87e2d46a8ebde77ac35b117e55716636c679729ec8ffc7992a07174bd9c262ecd1b146788a11b3780a361f3c25718d7fbab276519c375a26ab372caa7fcaabaae849d5767f3d3e1f17dd0d6ce81cbccd1ce2afda11d9af39b5499567a8910fa990bb86c3d1f53465fd2bcc60f6ee469b93111011cb7288b6efbb2998c255255875d92d43c14389e62d82222b655c8e0089643bee0ee3b297ca1ccd93c72430ecf16be114702d16825d9f8f0ef20db6c4b589be45c12290fa4fe9f12d1b17;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he0f2b2708ec7fc8e9c661f55d55c94acb4e9c10b246462b7b4b4b809fea42992a6981890e8128a2673486ff0e2789dc7b6ddfa49cffd132472d3f3cc454063bbc8c62bd19022c5b2fae5036cdfb7f501ea4ba5967b790797cefd94962453d5ba2601925e9186100f04de5917f52ff1ddcd7f2b1aefd7778318f791f4299634286d3b801b2ffac1ed6ea2c445ea8beb646fcfbcd5e7397b4ee0b2fcac5c22bfac345f976fa1c65eef533f20e10bfe1c3b5a46542633d0a8f6f70279466f80164b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h4336b7999493efd725201cd2451306434a4d2eb98186bbbd88d8c9be29b7f9185ecdc30f7b597ef6c051d2d776916fbee859e3acc978b066ee4317dab13d73f15935b243874e56ee0b81a5ff252770d06d752597f6f27b365c70fcc036bd771e25d7481d7af4bc546fc9533a1493e90d092c21b0f307a2393e2d00d5eec09b61bc81f634e66e0722517ab2342a36836eb7489ceafcc84e7536f8126911a1403760d32d6b3743666f12cb80bd8db19ff4ff619a68236fb4f35c1c5fb374c1dcc8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h838d90147738f026b1e2ecba1272178126af3b67ea683fb2b28804ab6b37d97f581ada303eafc4360818ab10ef0d2f183d5290d2a05ce695645f7bf5c2c39ccd72876211eef1da12fafdba7bbc1f02d4241d4b3fd15f857b00f61429d876c17a3d37c64b81bc0d295a130e2dc1ec44e256589961884c4d5a22b5784cdc54eacb836d80d5b1c710bd11a0a24fb2ee20b492c972049cc6d3d0204e0704cc20bde64b31d037b6c47ab39b1d8fe75120d3f3c92b06b5f41a752ce8dc15dc4ea51134;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h93923e558cffa1c6c8198f4085ff5ea5db72d62962c5ebbfb161464f5a6e6d880304e370674ee083e18ae017ebabbd232a14b480d6609f8ba360a7d90592bab963eace021a38669d7f36793c980e3696bfc9356a016526e194f55553dd7ffed145eecd2e3e18bb07d7c816c576209f2e39920b3c4d48ed85e61c50a3dca923693272e50cb1d6027d9d0dbff96e099ae273e2b301667e809c721d2306f227f2b8bea69c0d24ef02028f9a803cb6ad8ac30297ebb0e4eee5972498b5e35c015d27;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5f897337aa3a74b706b85136d752836b9b6f59e929325c321a474db0bfb9401394155080b52ffd7ba8040840b7889692d486e3e0570e7e5b1d69cd0f030e9257923ea4a427c145d154728bfd4552206540f17d3d12b7541168d0bf40059ac6f8c4145040f066a758a3cd3c4bc6e3b133d1e3fe85ac91e11e89763e5d4666e031cf2d187578537e9d4f03cebadff63f9de082b0ce3718505f4a4265ebbc6014995a50d09ef43ba29806ea555f328a66ac0ccd4d87277acfb6fd9a7ecebc221609;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he0c652a0229fb3a1babdb74e251effd44dc695e5e125e9c76956b10b865a1fc52e2eb6a85e5b2fd1623a78d3e9f01f57beeceabded8265f1599430373c577aeef16505713d91432d0c735792d112a754461c208451fec3dd5bd172ae9398159403957540e2537c2bbd67d29d77e1b78eb19f5f4c5a7040b8cd36f6b4faad4aa892c4c7caa432be2a42398d7d4fd4688bd09e6371549e4098055a1787b369c7b30782b27c7d3bef007ffc02dafbf497e30d9a6a0e62fb9e6d75bfb7207dc46bdf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h78b55450e0d2c1b9d77819611f653919f054e82a469082793dd74a6bd2411ce3af3bb9d2866be4f98adf1dfb122110d4a22a9a726a1f6776b35a8163c64cf44ba32c271686fc8037bc9457070aebc5df8031ca851ae5605a791260d700b3d1c3e80e00d400510d6c7a7cae300c2ea66529180e87f7779e2c0c4752e24ee78dfd8eb3ab36255a6f304b5f9805b584210724e84dddfb42a08472df5eddcaa4b12d4c247c067451b1a3f7c61ca79ee91b8db6f27a6a2201c1d1c2d2385c1ba5dd6b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h9b6e7d8b4a51b3fccaa65fbbcf3cfd42d55643cc654d4254268e3426a75896da82b1b58ee6f597c973a980eab1d7ab2aaf75523a902d00c0437c22e1bc6c7aa0560450824a8316e3dd3c2acf5f3ca4827b5d4ceefb7264de18d215707469a772b8e8a1d5cea34a45819c9cc45cc22a501c8c02d3b4d614774ce945d7d0f414d8b81a3de1fa9f12cc8d0dc4a20e3a2d2d7d20a751119a3a32ff2502aee93e35bc658d724c3242a89193ab9a32fa595f3c7f81a129e4b1c4244a40e98c683579ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h9db61f442255a4b4ab19e9e98c7729e73a5608b9571793afd8987d56620c9dc504ba016c01c34a3e8624560ffe03f42f44c12372b097242784fcc86e8891e424003dd17cdd48e56c3d729869b30aef7fdeecbe6ac0485dcbba49e888a13289ac0973d236a37b11b89a1fb9d84d77902a4f5f647de2272e3f880c52d62bc3ca42643c56b0faac13df7c39db90139441e269abb481de7d4555022eb244c6965962a2bc745781ebb9693918dd3d2c6733d08f292b2b6c5f348f272b1917e774c692;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hdbf804c2b93de72b5bc88cff625e6b0b6bd72105856f720d5cd0dbb61915fd530f5a440c57ccceb4d1a354a7ec14a74b5d18ab815647f82e6e6932a85a2b2aa7fa077aca6f5aba85a102e585770d84454e5fbe0856d58a8b2e35ba4a2e663dc7ac612275454c13d27844de276bfa2cdfd4422fb58c2e660b8b868881bb0f5cd6175e54eff9d6460b1d5338fbe4123e82bf9ce7c032c3dbac39b171a8ba9fe8d80b835089208a6c1ece1af15468b690bcc95a89935739b9cf4d6c6a684a4f38cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h6d873d5044face1e5ab54a33c17696d38b669b8b69285320daf4049c0fbd868d80bf0ceb860352ef6b9cb1763d6536173a2b25560a4bd5ea3f429cc330c84b93ca5a447a165ca963e401adc5d1e54329cdc559b287960b41c18382e55e3d237f3156a95a1edc3fd0beb422a42728d1b1477657f63532fb4c5f9ae4346a8d7f7eb4f49f72076b532e6558b3f70e9363d6bbbf3f9192ba46b8d7092192e58b6765677eb60b8a121e0137705476b3a15efc7c8f9ca45bc510fa63cd169365d6dfa6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hbfb23dc684c40e22336413b8efc5ce3fe71b66fdfb571f755da729d20ac3cfefb802f970034beb4667a47f35b3360af80e359acbf4fb3383f8c0351bc8ff485070a8ef7155d85eb1e4d323b02f41ef5db18451f03e6a8da78603b60733b7bf8319413432e5cc3322162b8b157000983b855b566017070b400e45435b611622d47e1a4c9de96867e027855fa89b1ac0a069ce4c5d1b78ef36d3d71c7262c5fea2e9d2c1771a6d8385ec9149af30c9bc30080d3921e031eded707513cbd9eb0ec0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h12b05f038201d44978e99570cb0722529f0d44a94d4208614dbf093a38aa67d330f6951c5ae1df944f49c99f3c546df9115822dc5592e8ef0a587ecfa92c1065de2b1aea2d69ab9c7e8e4bd59579b03418849c034c3a9e32923a292f81060bbd02d71c1092b5a5ee4dcaa2e29e2c028d7e2578ef3e5ca0ad1ca86f79d4854efabfb98d1bd2060524cacedbf0746dbf193121b2699e85fa1ea6a477a48896c7cd3892e54804f1ffd9b0f9214f56fae0647643e31af17345f5794c098b7ede58a4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf39d8e490f33be540b3410d028e05391dc4e2461b41864a264f796b296ed1520e7d90790df5f0350cf83818bef33aeb15ca70f1d80edda46fa98a0d3293f39a98005fd4d646de75057ab5d0047f3eb169c6994900cb1c3ff3f256d7ba0b5b89dc6fd420221d0ee121c9ce8b30fe6e48840816b1c61d4897c360af9b2e051cacc4cb5b35edeff68788050921c705a28266f27b00ff576bf96a03802879e91aff2b6d31194f5bec5f505c09c62af4e68c94017ca3d00e806de346c13a159a11c0a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h50412b7b1b16e72c26038020ccc11b7600d26f9cf17a325949733ab159c70d6517f4f4d5423f0c790839b3f19433c51b46e26df293138637c3708e98d6a5b719bb3b4c3aee4d39050839f890c2164d222ab7c2344b674e992f60983d77f1467036f4a5ec047a726a2d308124c408d0ce89f918034df9ed08f8ce060dcfae3aaef95e89e3b7e406aed0598db9e384e7c67bbce0260d19c1f55dbc32b77357d8246e5f35969c3030b5cfd368f7b09a3eb8b56c3712cb97bcca8ae4f49667bb3ef4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hed6bde3a79cacae3a068b8f8e4c44dc47fbef2a7a4e7a7bd69ea6790b6c01cfa4c9a484c3b3c813e92811c4d702671917e8da22b0020b9483232417188cb1ef3e4ac2326181987a24e87ded461afeccd9aa1953835a2eb852f86447bf365a9de4b4ba363298ebe6272b597356555a309fb638da5274ecce689d0fa02a1bd970414c428c036ef5b4ab7d8ce0585c2081b061429c537d714c1c65a69fb981c6109a0fb05d66cf11429840ec03479b567aed51896f3352d45a96ea5d3c972c98cc0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hebc283e2fc893ca114ca42a4269c8710b63d37fd63df8ad435dfb851134b985e613a5a658a053c57c2b9ed53609019a12677425273eaa128fb4bb7673497adbef189151f00010e828ac8ba98336f6c5e17834237b8315da078745ffcccacbe537bcc2bbccf565188760ced5e9b0f2fa637197644072f593805db2df6caa8d68d80956e87533feba7b61121712226593932e6e34844069917ee5b0420745a00e0640503ea943eb03f760066170ddd5687545e7dfc270ef9cd5c5ab1c7d4ebedcf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h4ae530d58af88c51e79f7f07d92121b0426e4814e214e61eefd3419af5072535ce31032586a2b9ed83e1d4d088db1c133e97912dada82a9d05a844348db2799de84fa9ada14c006d23f617c3f758fc6797160f6ad738ad9f13d65b64e28ffe6702c131c05ea1e919bbfd19be691a71b969644aa1838517ea3ad24b5e2d72f2311f177c72e405613edc63ae60bd39ea56e1cd14f9e9852b18c9718ad519bbb5b66f97f9db20b6c0c946ceb7b008a3a8e5a747b644ee246976a1f43ad97c16bfc9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h29e22540a3cbe70fc99b18d579b53e0c85438a9b2be263018c2ff0037b77a7db2204ffabb9e9efd67c0e2cac6274ac6aa7e3cc234042218b29b269b823d084fb64ffbca217bde32f908d63a6b4a870f8bb60b52344186754a0dea33e52867468dbeb9e37c9ca1c24083c489e7ddf8b18e6c4217bac48198d1a28da409b611e3e1ddf91e1b54d4d238ad4b54d385f58d39cd25dff0cc030efbc902b56c65ac5c886d3be1970e50581221f9f055138c14114dd91d8d826a728a195bf77056f1a9c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h3abe63db0ceed78f6a542ff8fbc1c90ee1dff8f51037c3e15fa2651291d459d1feb7d01dda48cf23757c209601f4ad3a8396c1bf3ec6c95dfacb9daf8a869d0725f4be6a3d3b12e11d3b1ece9e22dbe819965ac6cff9f5253471c37578885f1a413280cd69d85b782a9fb6a449e6cf4eb23aeaa84a526521a774782a88ddbe38338e6e420ea98e48d82615b0ae293b63600785b27b4a8b771cfc146e24a422dedece4eae19dab44704345396a76f76f7db8903de64bae1179adcb69f0d40c753;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h15f35b681da9dcc19ea6d28db1867d399c90a33daac4739a5c0913d7fe95b90b0e473a4d50ddf38581933daf8bfc37c8a50e45b438a470c23e7a77aa2626708de15ae82709061927931ae63d4085a9bd3d354d60ff87e0dc72196d3f84d71ef491037fe0137acfeebf96f0a2dce139df0cf890e55db30c603326f34fcfb50b62fb72df5f701197000f12ceec5282307f3b88d7baaba43a495149f48f7b4b398434856aab69261da706523c2172cdabcc34f090679282f1b2e468855cfa804d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf81e6ff424223e7223f4bcd7b2e545b9f6b347af3f160128691ff9d8e0ce62da79db1c59609ea736cfd1dce9181ce13194f81089fcd5ea224e373f6d993559269917ef98e58c2753bdfe281273f99d37a2a616685513905db89f67013d183af014902a7b9b9b6882a7684d6545239459f1a531540952e13b0fb594f6a41b95b59d1df8c9ffdedf01862b7143aaa4825633c5e8b5922ee9099249df28c1c6335eee0666c5cd98a5c6e4bb4337931c5d6be45c2630f19099d69312a60abf87fa46;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf64e0d990dce10e62a750da98a6f03f018a4c1d624e8ead9e8dbabd55cbe5bec9d392db80dce49618a7735c5a8bef7ac394c149e2ca9ec361d2ee3e56bb487edd54a363025b0529a5942b1fbace1f8d4de8157a8c72adab80bd2e4f94971ce8ad3c9014688cabf3b3c50a6605d1dac8614c18ce03bc34dd5173b7d9217174617a0ded6a9a9fcb8a5f09e355ea7f12923df02e75cfd05237646a53db407ab710f36642da5f586db884281366c5b578994d35bd8c513362522b39ab5c22285c0ed;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h782ee5613bbf11168cd6d304a0f5c1cf20d82490dfc79d165946b21d57ab9d8a3cbe60dba4b2b851aaba18aea17fe6dc91b3317675c347496efc1290acdc8e958f3ad2e31dd13da4947c6c5f4fb963ce535c7af35c52209dc51a140903a86dd08ecb289bc037b5e7e8d7caae98ff2036a4d228dc65a6cbcfd95f053bb78528786e494c14b930347818bcd5e9bd723253fc260f22b87cbd5a6836220edacdbd0363dde135f1a854125032b2b87f6f4c1bb7fe9b55e89dc1fdfb81f7a4ef66aea2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h977b1add59d7905cec2dcbb1e2f809431a6c356ad07d66f54a542d93cf0556141dac35194b673eccf83ebce674731d9d1be90689d3ba92e21ce250cdf9cb7a1b1a2cd5ead54fd952eb9fcceed2b27e32ca2a66e325617e66349382354d3056c568491320c0f9dac34b4a709b72fcaea46910284eb4719bb82fc04dac740be507bb22b0ef117f27001216c7c4698d9500248b4401887016a14703c90a533130a8e4286bcc17ff9e2786cd7b7278204c6aa0099dfaee20fa7044b551910b1bd525;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he68e0e5fa86bd930355c815332f27b25a25f9536191673fba4151f8d5aef8120b17599c85e775bce05148a993ee1f68da9a4501ffb0accf12dfdea6ff34d70106c45969bfb7e2120843001be619dbd8f80ef23f5321b79d84c17db529a32fe0e3b8b0cdd20b87e9c7a3cddcbe03062e5e238f337fdb982b096324178f026b00c09c6a4599e5ac46dada2aaa3c36434c5f2d9f71ef35d79e1658f0be3cd16ca680466355245e62e6d0b4be65847d0ad46a920ea2af568233fcce28c7be2f8ef4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h599fb6744a7da9c428dc2d8d875aeec799e26639678394151a25d71cd7cf9e528a7d8715f93e8986de7e88847340ef85ff2a86fddf4a855f4d05a408d79690a0be2e964f40c66a2d424a5990f0885fc2d50ad59d7188133a27945e462cc740b7044d602719918e40cd35a2fc16bc64e7a818c80dd0b97e66f37b3496bbba2c229fbaddecdb6e54413987506db0abc0683b7675f428a0dc60a1ad2803de03bb024327301bd2a57d58af6845c87f59e9bf5e0a332fa6139b4064da32acd76f6ffd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hc94d787042a3151a69bcbba6930aadd1ac38ac9e6bf5e746851f993725b43b1b45fe47a4dc5b20f13be0e5143a4aeba29d28b15ed16b4a437b6b61d2fb078c9889c7638406a7ff936a67c7d9623d67c5676f9463a915e2d4cbce65d2e3a86638b9695bd75bbc20dede9270dbaa8ec8e8dc98c9057e89fff8f660c247020fc3dbeb292e8714457d2bf09cd4fb554b24dd400b404f6179f4a23dd73493dd696f826fc64ecec9b04f0d3c59e2942d6370e1e036b85e20fb21b06f1c0cfa6579e36e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8a84e131b596c898504d10ea539b9e6be66c9bb0f508fa569416e8a0ceefa889eb53bbd4c033f759defd9c2ff1a944eb913c952a84b979afd57fc3d74656cac56ee38aca0da8433c171c2d545a405da2c770e634b13e461bf1670019c7e215144791caa58a6c54e8785fd10018fc6246f691f7972042868189a93cd54699e2021357ba997fee878c7ac31c5dab8dca2cf8155cfa0624f546487079abe24bfbea349966629b1932a66615257b95d7d935a6db0c84b728c1fa49acae4c98108823;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he77fe5f4c8e9c2949b66a6f8e55047a092ab82256ea622c73029d2a895bfa38c9b86697b94bc9e8f7d1e7fb1cee540c14bd77505f24bb4be430953c6916fa21fbf4bda3d275899713d3f53c6777d8d9c08803d3156cc1cf3731367880414de2bc929a67bf27d9adf14f40aa1f49d1a54c33bb44ac0a032e3e9e3d5e7f22207891597d90092c2ae98f6812b67a0e634641a83fd1629672d5cbd5ce7b50ac4ce3f333a1bf4eebcfb82167ebc285f2b6a1b5598af3cb7789bab2f08f09261dac60;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h2e501e08d8c03d9c3255889508ab22298b1d0b3baacdabdc46ff8f6d5667c8a270558e9f9e8e7ca5715a427958610128b32f24e41b4821ac02c38d52432033c1a2c79782deafdb9eb21f4b5229d5c9f69f2ecf0094b347d68dfb922c937a36b32f07edd346c0f8729808e5354faa0c16b4431753c1944373f825ae11112764d3f58349c5ecdd6076a2c81a1abaa910722ad3ae66f76130ff329bb6aaf3346415ac4420fe88ecc6ddbe5e39bb17d9d0409fb6174561eed3595d81ead771b5a44;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8a1a2ede1fffdea4c64c621593be8db7c4ddaa33c9586c4d1d6d40da953fea482c2090b48597a70075e4fc50456356c72c9e386913a099aaaf269cd1ae5f853b0122a4863017d9a580d060c9351023d46977f91042e280c9de694c5d92dd8dc8819c8d95edf6f9462ceffa28e50c0a0e2ba3bd79cb300f2bb1e75039482224ff0486566c602f27f43fcc20d6fc9a0ed3064f8602cdb65fd273dea7ce455c0f3f779607f62618d03d84d9efa362932d30ed3756bd12d774ac7212364f4750a2d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h51bb087fcecd9209ef39414286a4f305ec8c9fc21d13ff4e9fe27f006470b0b0b6c931a154743e0fc7a94495ca46f3c27e06f58b25dde40912936bd1ef3863001e26c5108a40d6ffa1fdfb7e242f100fcff72cfb35d6fb02a0825c2035f6882184a09962310f000ce63eeb9cf26aa5472e9cbbd31499ff0281fcde8a0a79b8678e7192fda931752b51358c18a6c4b86adafee3fe055c149ab68f4ed981feabee12ba5c483a7675977c3b44b9697e1f0f776266a91f2cb055a81a65ad0c113bf5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h796ec2a39ba93c10abcb5637325b01406bbc54106dd56b51abfdc867b7067fbeaa1b55351ea5963ccb38ce3a08b82bf446ce3d5f8b213a109ead6196b2921906254fdaaaf7c0bd8c15beaabca9fbcfa9783f4c59d6127ae58b03430b681c782c004bc04863d047cd5529c95b78fbf481c19902b722503282bc0577284d4a1f4bde13c2f5c3ae9fda75b176f29d425255a170a45b441ac067f55abca1b0579bc512995d16528d512d59d7d7fa1a77b132ca5b70465f3a4e204a93ae654a801966;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb1f116c5c3952b87b80b0fcafb4b20cd369f71771361c416186c2c546c27e338ad53c4a076e6a60ae209c137a9d557775d11d3c89d03bc60398fa6a0992301b880f3fec9b3716f0dc1d80a82b2e8c31d6a507a79137954648c672b8bf2433daf06c1696d8dcf61202fe1e1778cc70df0de68b5a67ef2ed9cacdbb4d106677eeb467cb646ad180f1e0dc0d690dcae0592117038d947fc5f61e910af53ebd70c400dfb7ea27f25c49b1834a6f7414bb9554dbdce05a1515ff0b742a2f91fc84d91;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha4473a27902bb57084e25e04c62fe1bf8914c2fee4e7eb964ce2d6304440a4e0cf4c81eb9d8510ca2b39fa01008a92aee2ed7124e0ebeb40fdc954b2cbb9097e9b8f1ba663227137d285ca78555b7e10baf2684b4629bc6942416170b70374a18801bc3edc3913d86499cc901d33cf2ce4c3279d86cb5e08eb5f216a3592b6f270a71591548481e16b94c1be9c14c7e446bf12820baa3793f26df1199cb7554d767aed6f6fed262874b2e70f43ce3665e780e2dc98b7a0cc6db9c2d08a44afeb;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'he54cfcca26512019765ac5bf0df6dc13fdda11abc71fbf3ba17b8841b9e0db2bfe3cc2dd81c1127714faaf56d7de5cdea70c0bf797aa26e7f98099454d1cb3d0475d10c118256e35d62090a5d5100934fdccb96d61ca94bd942a3e3c09fe31f8d20ab29b787f2529ff23b4c0e754d109bd0708f1032510bbf1cc51ef51a83919b3daaf0b7ae442027bf7def0055f74487f873e12c9bbfccfa4dde681d6687d02a95c1c9ea66645ceea6d3318347f112ebb0da5048b298deedb99ca117bcf8057;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd6c31c449a35c95189258dd297dbaff22fd6c6a6d4f180c32888f0d7f73c36647cd2210029fc87f493e8cf0e64da1bf08afb0cafd8d6bdff93d1f93d968b2e50cad25606537a368e8d598992d60570a804c5cdc5b51dc6efdb7f7c3330085391df70041d0795bd8fcdd78d37012ecd39e3a84e0e8eef378ba4192cec8b5b27f347e631deb5be7e54949bbe6ba8c22eaba57fe371b931dedba876b5d85953a4dce17e92f13182dba45aed6f0b6dde917b600af7b108e05f219538af58261ec776;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf421d677c716be6e8f63692ed336cc1ace172c64d019001631f6776b5d7a8f5452504342d59c35394947850b990ebb4d6b0a85b118d809802b9043e964996eec56bc31913203a42f7ee9d76648ef0116bc256cc6e12cc82a38b7b413a5174f061625a954e280ff0088864b3614419f870395584758b151000bbb9de38939f75f4b43e03a611ea81c5fd8005253cafc56d6f9955a52a26db41236288808a911acc2c7e6c3bb2430c7e2c34c02344d036b9823af1bc4e2610b76b6f428f506aa30;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb43edabf042c2cbe2fc234cb5b99b2f0d67179f90c7ce0a49716876c023c9b210c3dedef4af013663c256b69f4a0ebc34278bc168da27c0fa1921e495d41d8e58daa6f6398b92631e48c45a863a2baf52efdeaaaf72d6b49aa7a34d0b11984e011857824698ac9a3dbd0094fe6214afe2008660ce4a1c235ca2dd2115357ef56cd6650ffc023bf50be744de40071c7336645976747c2047d84cfec6688687fc65b537f700b1490d1cf150a9f3cdb422dcfb5806d01f3a66fe18d8e48c14f3e55;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h9fb7b3b6a0c1007237e8e20f87d82ae36806b47407108835f5eacb8ff33cbf64d410ecc89e55ec1563d3829c268b051be45875aaca5ec1363ff495814fb6d4df74599ba4b417f3f8730955d93e2cf8827143f2b0f58a644f5ddd1974b0fa8df9f5a185a3d633f39988ba975b59ecef14efcd8e1733fd4ec9ccdba7ac14b651b99a4a69c088a2b1f7534f952323e814becc677a17519e54214b5cbeb0d3d5f5e769b19d1365f697557b5f07461213adc8e1421d7815a8eb0dff5a97c97c421814;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hb3778c9c723acda2a6116365548bbf293dce67b48e276da772721f1f2662b083170d1f4162d2e4788e62e4fbc74113e320e8314257201e306eb017f76cbf1159fef8adfeac25226c176fa494adf28d1b20a387ebb58a3d2a3cba6f4fc465540019f86f5e53bd988cce36c497a4058260718941c2a2f9a857668de3dc98916a651e46c75cec9254250384eadcaf05c5953038fed25626c4434680cb8376705a1aa6db0b0876a562444446f8f6cd68d5a19c672c34d5736ef7b49dd575716a8d05;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h19ac3acfa3135a09d67c15f5e6aceb53bc23927c1959fe2904068b6eecefc28dfbcfc92a92d1561c72254991e9c4a2bf2e5fb8e6b64d8ae5437e6fa4884d8a74696028f17d43a6d186a1c309ff1f3f1c0aa5416a6d84efa1e14a05ca11271d6a62fa47980d1ed0fab41d5913aedd875f971bc435bfabcc34b648fbdac50489b62aff8603abcd471f6caf713f6e0161da41ada65f4b3580d6ec97ede669d01d75c566bb09b188b70dea91820fa6090bd1261c99ff55248e44b0b97266553ceaf5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hbd571d37f976b5e218b4f5fb14d89d30fb91981f1e2443db61b2ccddd0a6f47bee6676471d7717f4b874b00017c1330ce7fde819dde8aaa20022b76e8f0fdc0bf4c8f0b2b9f9a1b6d369dc1c78f403a1cab62a9547ec3c1629132464b1b27688e12f27195c7f29bb90191cc5bd4384a4d08abee3bc61da69c904911fe1a777bee93f9e5602c823a3cf4a5e925cde92b2a209a169582f35f289bbdb58717437d2b14b7043df46bf6f076b3f07d72ff5ca58b263c77afadf9a222855b27c38f211;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'heb5efd1b82526dff6d9194b28ac278b25264ac16b20987997c61e72f623e7760f05c8ca45aa4eaf17bf3929b6a3cc49978873c911b7ecd114ab3ef3bcc3decd97d73b407dc317ef91e3efc0b14b92595fdb8aa77d6c77f155dc5b81faaedd4c1806277c4d07bfd4b9db3b6b4a9ffb8fb05d7eac99d7746ead3d2995c31eb7b6d7c5651452bd8bd0cc9920efe0ac726e4cc229896fafa80257daac04091bbc3529143d669d1d1c2276f9893fb257289b0e1fe63579fe160c22f39d3eeab2f5901;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd69ebab7bf7ca11c745f847edb7cdc61273070dc0175937927b852443205e0cd5615febce14871117128999145f7e7f386db23b8444f931d1122d315649ee32bd0fe254e19e09692a72bc8a7296bc37d2c6f4bafce27bcd1bcbae4bae83195f4cd161dcd200a6a8476d3c097817b3c111b933a7f7f5b67fb46f4e2fb92961341423d60eaa1e5fa67c0e3923cef38cdfdcb5baea03bad9d20d5ab280bd7abdaeb70510eb5bc1c7300270519a678ed5d04dfc9b5e46ea03e1f05c3d18e293847e7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h6858c59653c83246d4dbc05d482420bf5a62da3847256a002032904aa45596b7cefc77fc9b22803a1a4afb92ac5ccbb05a11592e692a15c2a65945082a1b560703cc598358dac91bdcaa36637daab2b06ff738e95bc16b53093b9cb683e16fdb2ea1832cfc24b30ed208a992800aa0dbabb47e3909da00067d777ca6ca65441aa4cb81b7521351c70390747a1cebf4d7697caea6ae9e7e84e01bc76c9ad37e4c721558ef51177c1e34ab5d1b49fcf5f0fcdd6812046b89f110a2d365b695152c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hdf9f9582b848047462adca99b0815456af817352a6d2787be5de41bcbccc0c5fe54c70d390a862dea49e5e5d922082eb0476e8404daa5ad59a33e583a6c8c34a70b162a3016638d992ab8bb95784e7c1482c3b91902f522bb80cb236e759f62537fa1a04dca08630a63b01b0f7b59b744bccab576edeb18b1dfb391e15a0063f0ec7a5e562cd4798988a88934661a1e3e4ae0b0c71e633f7dd621c9fecbc3b56944b12597857b4604151ca6c0c4d55d78d8f98873aa41c7aa74e12ea6e7e3fa2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7751ae3e83bab04b0a7a6129132e4f9b6fca2458b674d1ee74aeb528af75d8f6868f7cc068db9099c319a70de9257c1e7e2437e3af67e8d4143eb4db9347c6b49e0c449be107036cc6f9837b69cc682a844aaf8933ca48e5621bcfefd4f42c6a9ac3506c05edbce1babfd14a1f0a34a193ac41763fb73966bab29696c4edbd2f7cf6008a62c26a82d0856dabb5e8e74017267cfeebfc6880d4f5d1a04f6d64ebc4ff304db3d6671f8d263af3503512b20a015194d520d3c623afa05f3c6b7c1c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf5d0034c56c42b05ce17faf27c06af647284532869aef13835eed7639fefe792298483e78c1b33f6183142b719432a978563fdd556461e94fe727b99fcd77f12c2cae85e81dfd94bb4a09acddffc154624b6fd0b626dbbab405abab6fef9f1cd4c6a01ec2f0ec3551c7941a565cdc626d3bb2741162f77bb01d6c3c5b5deccee88394ca2d2beb3677651f906f18d7e732fd72355bdf9b8557baf6c18c18edb53f1281a9eff46e2bb2c5963b1448fc223e7f81f2fa74a637afb3f1cd2accc9f0c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf4f5c2f26bfad7f5502f2cfd257b685c577bbdd7b9d3e929022870730a666b3017a4174bab58082e11ae04694a244470219398c98414e52c53e2bd431f77234b7ddb205054405bfbb04f959eee96181ef927299521f7b2b5ceff67e6b143c6e7b45936c7c8a6eb79fdd7fb9c4df644018f01bac53b82d005264f48f8a5b43c30e7a109eed5dbabe8b4386edd947814d23c344399f7d4c1ac371553a6c1343ca1b6fb1083bf00bcbfbadcc033eacde812ac7925f59e19adf8a4c4daadceac248b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h76ad89cdc214cd5c8ca633f98a39b4601cd50010088d903642b4076b0fe1201a25b60513a847ce1775b91cb16536be453e7095d14f3c0e566fb3ef9e383178d25ddc71ed0d5e1ff9eef55f090a2fb06e31799ce6590b8b8c92035f0d4ce1ade8904e189cd14a230c4db2ff79c0a64f57f59c6d9fa108091a904b4f169b88707d0e66a9f4a1a89b3455d2bfe6144c3ba27fa78a316102683aff44bf0d9e2ececc13cbe95f6203519405ed934b77900c481065e063392232160ac7d2a235c091d9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf936428d56f574e0a868a07b7ac87f2660450b0c1b1043206b426eb5c6700fa2fd4bbd21c7e6e04e624e0c6275940abb62b6e746d7f82f1e1fba635d24f3471d4a97a7c31fd2a39b340cbb4ddb3e4f0db389b8dc8b775da137fa65bc17ba1db1ab6ff03de14b76f7672ee1ef2e7729bd16c416e0b796824220e0b0b3eb8039978a73404faa0a6ca8e43014b49c5a010d97a0ae06838915cbb4b80651aaeaba1435956773d7c80a0751f1383fd5dad09c075e595d73b42d5eb2aefaafe4acaea6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h50135fd013e81050592626e630324a84b18d83e3ad1a0865596795dd14953bff99f7272ac2c6a2753f4c4820542f4d269c8cc86d6761c9f5e3daa5ddd993a765309739dec3eca038d37d690cc83968b5e48a75159aa1d6ffaef655c5c97d39951eecec679f2e0dc0516bdf045c4ab52cd6bbcd0f842ebf809689c083d90c06bcce0087506d95329f3f3873650d604a78847dde2fc624be10a1e3b1ca72c0c97c0bac25492689572d11ba68310d9541b054ff54027fa78b9f1395dffbfaa8009f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h19d01263d3b2618570319fdb8e2fe4574b8debdbe5ed8f23aec52e5819228a1a3ee006bd53f4158aca6837d8beb298d1a29aaad4e95532f7bbb6df549248ce8339fdf7917558784fbb7b448468e13b54eb8b93a8e8a447650b56ff484d9172d71c8a7aa48364dc801966150e0db1d1ac7bebd9f090b1c451a4ebbc8d522fdf0088aedf3a4368151cf947a9d5e4dc709a9264e0b632e1586672aff38d918fe5ce22beaf3d98f48f4f2855e6fb6406786054ea0b10014cb24d90ecba37191187a8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7fff36d58c6737e940f50881eb53b6bfec92ffae7464b584451e859e5c619e3007d215f3f0da56642b47835056ea38eba6c467d6ad73ba612381f73c96fbd08ac7d80f7fea847462f891b8b63739393688cc65c4401f6612e49ebe7170837f02f0aad2575cfd00714e402531b6d11510b29b6b1e8ac7ac4537157db4dfcf08b88cadefeb1d456aea289d17a1a2117f3c55d0a2ab994b6c28c6cd972a46d4565fc941fb3117c00d0488a4c31140f9f5490f96b89aaeaa6ff65bd396c3b3411421;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h30c25a9d9498eaac9d1ed5d92f5581a299b04ea2cca5a2611321af84ff3f1a5d1a35753e17175311ec343e0f26c3f44640afb6ccf341623350526058ccdee1877b9647757141dc7a92bf6ebf6e6056a983c67a2d4c1bb845ff8a77c7a2b01b11784e3ed311aac845a6a6c37016746d7fa39daaca90a88de2e1b2051a595df4571a8fcf98f3a792525ad2d5ba52a3de9471e69af1f9a7d8d54953b3433bea9b409a604ed80d5cd4977330dbf239dc80857deacbbeea554dc97fb89dd821588c88;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h40d47eced0c7a319d34efccfe50fa06c0bb0978b21081343762d888f191c0576e62cd1c06de950ea5b1726bd7f7c581b954aff1bc92e713a53943a3b63a62c632f0b4ed545f858c5f467353e7b2b9cd480d51cb5d5d2c58bc8af0239e2fcbd5e8a01b6d8734fa2c70692d4b59e6fd2d42e789a0256a48f3327e2918c1d29a9c2162567d399548e7cfd692a74837a563011621ca6364fc1f0fdcea12c226d936f7a72b6b7067ac14b941966b9b23898bb75aff3bf76818fa3cb02ecfb9c6a9668;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha93ebf65c4f225a8d6183b020963e8014d4e8c458a210e704024ceaa92792c107c974be6c8d295780c747abfb7f6a10ab6bc5df86d61ae2e9b114e738dbca761699b6a1c438e8f85e5f5be656be4be5383bbd77152b5b6a7792e571e0d12a992bfc3e8f3c77d89f3fb02600b84b113e3bfa5bed649f7753e356a45082e5e01f462688348e6cbf7c1f86696492f77d8899da07d8cf7008d7b57df9a187203edac630c70e0553f21c712e885fd9587565ff42b2801b52cc6c9d7f3bcd00c282618;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h4aa4c7646b04ef8d23ec81dda6d182c5c40f9ae84fe4f0b3776cb9dd0a6ed02420c797fe32b2bd608fe2a0213fdea2cb3f838b940de4975c0ef975238f4b84bb4af168268835ffa0c1cd6f3b866149ddf166d5def759f9b1b7db1396b2e3fb287f9ca90fbd36c5947c1633b621ffd98ba0365ad8539369bc49735a4b19c820893d5626d6c9024cd0345f350843d4c0ad355d91c491b8ad17a46ea15b45d9f0bf40d90a9d844f89a971b027cb6e78a1dfd9d57b17d6192035e51240ab71c402cd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h48c8a7dc6349582e920f965799d1c6be41ee491967833c75af09f52b4bf03a73d3211cb9f729000771a5dc927842970441e3014cf1786c2320e74b0fe27f713d701b7cc3f785f283a208f1b9d00d0f339a644e477a332c4e78967e298bfa419dec60046c24888f45658602445b789c182697cac14f9229a9fbed228fdb07f858405cc4e0bd5b6f08ca897c6ea652788d608a3339ca7090ae403bf9299597e05fc8edb2066da3175f5051a1159a050259cb61a8506684e951e3fb1243511866a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h5fa0bf982d4cadb9a0204dfb6c4505dbd76f22cf3ac99a035af15ca7963b5488348cc782a813c842341f1bd19196dbdcddb139399e37aaf5ed99ff2ffd3d31de8e7592a4020aa9038d781ca7e0271bf9e9cdf8cab031e97fe2c32e90a9096003100f7ac64c303414c742110f8fda252cd7ed588093e1b46dd7b4d1057811c755edf20a991de1829561bed8042ee1a501f59179cf1a961e7603037a061890a96279630934c7491722b75e3718176d2a49128c8392d8962c6f40c56ad23600281d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd17300328864d0fc4b71d5f1e1a202321ede8c9a8440f43a2df06e36980892de03c86e40a4e513ed8e87bc35cca4e555f0f606449c522368365cb3e7a363144ad7c97b3ffb32d64bab456ba7a2bba0b0d5ac7e3c7d6f00eebbcc69e74bc15a6b1135c41ffbc3403e5b2b05d04afb0d38eee537a16e14e742026a5bd3eee178b09d7bd1334ef5a768261e765837e83c158f0be8db1cc0f46be359558f541af339762e9064bf2ed0407f3d99215ed568cf96080b2f930566720cf4f06e1f06e250;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'ha9985439a110bd6d403cafcd784ad486cbc125420729eef3e766d1626bbc59a97c3d5780d452e399d086f04d428cdad60324085c0d9dd092596e0d4087870e75307ec8f0a66450bdfcd1c4f3f698af2327786befad4691e874f679db846cad1e692457cad27816013062daca3139da376bcb67149e57b67d547c66bd1d01261da6c595fff60142dc663eb70e415b31765fcec6bea528ccc2b521a9bfd50202432f776fb59d730f9c88656f2717862f5569b8145c85ebd8a3ec3e09f22db2c9d5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd6bca7560fd68ff88b085b0e6b7e4d972c24c7a8fa0d288c1dcec0792b2576ff115442a23b6d1464a7b40b39cfc9ea90be9c0ec4d97c10998d4ed8328ec264b9cebfde178e0fe5604cf35c5904ced0da69cb0e02aa8508c63f0ca7912c545017ffde4893036778d27a7ee88d7088e3b07b779fea2bc17f5e4d92cd6590fa058f253c6c10fb30bef67d60821bbdf3f39c6829c4c238d0658f57c31cd69dcbda9ddc456cb89d816ee4366400d1d41639d6cf2736868730c29aa76385420f866513;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h4d8b2ca9acd065f1d0fa7a6bd2d500ed7ccdbf09f8222114aa6ff7c4adb11f3928bd719ae547939f594e23b2f379d1de9b787dfa3ed61f8fb19db62a9404343c0c8d6860603a39aa5899f0ee46ba4a292c0950b302e54276c4a255f1cf253f29694821e524a37494fdbf694b8adc2d76688d01a53483cd5ac020b0492653452a682ce13730554fcd6a7d23811b71bc976821646b61f380e46cfc4df54a279f546d54d7d5f024c6a11324cb1fa6357de0df8752c9200ac1d5f89b1de3862634c1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h116b0381042b180e29dcd571cc2e5f55464c42f388adafc74e44c990a04f99537928e8fb79b791cf7ce28f9bf9d8d57324b6c606d6d5c2281b04c8f87b9f49c81266b44b8ba890d1ef9552ad2c28829aec0d7dd01136e7addbccd769856b84fb541e0f11543458a92c200a0ab9bd28bbaaf4bbd50ac81d4015c221f4981ecb800e0147bc01e5fce34eaf8af20c8b9f92ff6094048babbe05e71ce8e8e4efce8abccef431aca673a8cfe861bb82d0bbbf0c7748f17d57c7cd7caf22fe2f7683d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hcf2fbe1fc2fd33aae11af88204e2f1af2dc06f402042e425cb68ff89209840f7ecde34cbd6951eef1b57d2d2c48d78655662ec8fa98719a0d575becbf66a15969d00dc288b75390bfdce64ec4a6e6d0b41fada9a24750ac5ca97cba1f89fcbaa7008a467e2a17f5ac700476fa0217e5b7265a8a4477a7f8df49e9dd27c4574fe7bbc83ac4e79e4c458a24555a5f2e2d7e71fc90a79350c1b9f314168a6500d68cf9a4cb94247b57ab8787815a6645c1debcad3ff09833cbefa1002bc7a2dc937;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hfaacdef58d4f7e8946ee2aac087a44fcb64d1f2bd4dce196fe37d24b82711aac7393d30ff1c339a25ccde71ea9527c2b519de270cc706bfd950a131930537950a6aeccc9aac5ac930ce7fcdf6d65002decee423c978c9ff7edd2cbf3b3b414435b6a27ad224fa303e097ffaab3486efa055625bb39804ff6afe73a6e4784f9a269f54245ab853a0fe4f2c429d929066a9749e51b6e21df81e689e0e7b1d2435a1165ad4f84b88c36bf5195d752dbe0ae0c0d14b85e9d189b00468547e75bea49;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hf65ccc967875b7f8e9ada813ebc2563bf99e4129076a953654f86af5390248c2ef8495b00b5e4695c01d693530152345ce350ec42e3383604ac3e097ddcffd88c59d5a7bff64f3f416f7e53f39918cbc47b1b677c6a92dd745b632c38b8a1041fcbe9e189f2ecef1940a07f0d6640e81191c2ae080a439e65ecf7666e9fcb870923f469554da0a1b8fd68e7f1285e7864207723a86b21a37c67ac405cbf810d89f3199bfba4c8907ac8f230f778fe0b379764e0eeab70cde6ef545723f402fc5;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hd0001fc62169137e1c991379b8b1627353cd7e8913e10f5b8d82ab1f1213daebf199f7cb4e092b43c8840b154b3df44e52c8fda4f7b661be1f497bff9271546c9a15fb9177b5e7af5a2cc9b8efb43bd532db4eb1f45aca7cf11d3e103e79df95c30c93caa9a0df83bbd8c1db33bf7f6bb454ba851987c063121a69f6464b3cd2bc9af89844bf88d39297df3274f686d0b3d3ba00313bb7d8bdce6993b3ef71c3acb6c330dbb2a0e50d320da780f706752298c6a1b64c896d103ce0b67d4dbcd2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'hcda3a8e60660768d6c4d97025ae06816b0d946c11ff7b8803fe43a233c46acb204b06643a242f0df58dbc96d50cf0e435975b815aede88b157133e549274a3fea4300ad4741f34a60c5bc8d90e4c52d2a0e1f9d6834162b2108388fe40b19e7e08dda5b1d15a78d18038099a7cad056c735d343dd83b4f37a392356d0b70c2cf3725d81dd800f222ba3e0ebe031de84b2f78bd0f03978612905ce16d70c27bf0d9e844b502c88f7e4539c66cd76fe1befa24ba7e29d5c16447a1642a4009e80;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h7842e8999f6a0f8d191e819d28d3462445fe665b8b9c72133a52ec3949e07596e4d51168c69bba6aaaf4c3aec940c4f8910bbde8e78e245f615b82dddad28d743d1dc3b045afe39a66663b32826805961e879129d2d90c88e64caf75cc7cd9d51e2cea6537ee23e8897b1f64e18d79d259ce227cfd249f3861994fe627bb1090147acce8f85fe04751a923f27ab2eae9edc05a78b3dbc26544a7625482eaf1e24888625f790ba3ce257b4275ab52336ed9cf4780f0899f2ffe886c9a0b553c4c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h216c813ee738460401de48950d5020b5f7e3ea28943dd59731ee22069d6556c06e74bb8a70ece5be22e10159c374e2ba4fec877371df73d4d10886e47a68585c6ed204e4eb3b900f3b48d463c2ad57c4ec598230de85db8dbbb9e638cb7861afb731c4a9bf69ee9e5f6e5246172484cc9d3b5c9eba3b011f60deefcee96f3dbd9bfdace916971530429ff8272f2db5efa09ae32c56b3f63f41ef6c5128d435565fd185152323b39eb9998f165224ba676ffc0789450c3dbda84b065ddb4dd5a1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1536'h8364fa80544281ea380134bcd4d30b2915458108086a8876de478ab782f9fd899a81ccd0ce99bd350196819c963c9e1eb0e151755c4b4a630e2d7d564f2922b4fb6d4e781c65f95d89eb78a01c86445d040828adb3ef78156e429672f77334195c35582d3b3576f128b431df571208bafa13a25dfbc02e8dfe30be594b0f82fcaf0a560d2aee3dc6d62f9b006c82c279eac898a6b6783deac93653bca56a933cf2623e5a104892bb417405a53536e93c17049758ba044d3608cc63457e5b0a12;
        #1
        $finish();
    end
endmodule
