module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    compressor_CLA256_12 compressor_CLA256_12(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
    end
endmodule
module compressor_CLA256_12(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19);

    wire [1:0] comp_out0;
    wire [0:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [0:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], 1'h0, comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], 1'h0, comp_out0[1]}),
        .dst({dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      output wire [1:0] dst0,
      output wire [0:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [0:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [47:0] stage1_0;
   wire [89:0] stage1_1;
   wire [84:0] stage1_2;
   wire [96:0] stage1_3;
   wire [126:0] stage1_4;
   wire [128:0] stage1_5;
   wire [88:0] stage1_6;
   wire [90:0] stage1_7;
   wire [154:0] stage1_8;
   wire [119:0] stage1_9;
   wire [121:0] stage1_10;
   wire [82:0] stage1_11;
   wire [71:0] stage1_12;
   wire [41:0] stage1_13;
   wire [18:0] stage2_0;
   wire [24:0] stage2_1;
   wire [25:0] stage2_2;
   wire [41:0] stage2_3;
   wire [49:0] stage2_4;
   wire [41:0] stage2_5;
   wire [53:0] stage2_6;
   wire [47:0] stage2_7;
   wire [70:0] stage2_8;
   wire [42:0] stage2_9;
   wire [49:0] stage2_10;
   wire [46:0] stage2_11;
   wire [35:0] stage2_12;
   wire [35:0] stage2_13;
   wire [15:0] stage2_14;
   wire [4:0] stage2_15;
   wire [18:0] stage3_0;
   wire [4:0] stage3_1;
   wire [12:0] stage3_2;
   wire [10:0] stage3_3;
   wire [18:0] stage3_4;
   wire [17:0] stage3_5;
   wire [22:0] stage3_6;
   wire [20:0] stage3_7;
   wire [23:0] stage3_8;
   wire [27:0] stage3_9;
   wire [19:0] stage3_10;
   wire [21:0] stage3_11;
   wire [18:0] stage3_12;
   wire [12:0] stage3_13;
   wire [11:0] stage3_14;
   wire [12:0] stage3_15;
   wire [2:0] stage3_16;
   wire [13:0] stage4_0;
   wire [5:0] stage4_1;
   wire [3:0] stage4_2;
   wire [3:0] stage4_3;
   wire [6:0] stage4_4;
   wire [6:0] stage4_5;
   wire [12:0] stage4_6;
   wire [6:0] stage4_7;
   wire [11:0] stage4_8;
   wire [10:0] stage4_9;
   wire [8:0] stage4_10;
   wire [11:0] stage4_11;
   wire [8:0] stage4_12;
   wire [8:0] stage4_13;
   wire [4:0] stage4_14;
   wire [11:0] stage4_15;
   wire [3:0] stage4_16;
   wire [1:0] stage4_17;
   wire [5:0] stage5_0;
   wire [1:0] stage5_1;
   wire [3:0] stage5_2;
   wire [1:0] stage5_3;
   wire [4:0] stage5_4;
   wire [1:0] stage5_5;
   wire [4:0] stage5_6;
   wire [2:0] stage5_7;
   wire [3:0] stage5_8;
   wire [5:0] stage5_9;
   wire [4:0] stage5_10;
   wire [2:0] stage5_11;
   wire [3:0] stage5_12;
   wire [5:0] stage5_13;
   wire [5:0] stage5_14;
   wire [1:0] stage5_15;
   wire [5:0] stage5_16;
   wire [3:0] stage5_17;
   wire [1:0] stage6_0;
   wire [0:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [0:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [0:0] stage6_19;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[2]},
      {stage0_3[4]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[13], stage0_0[14], stage0_0[15]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[3]},
      {stage0_3[5]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[16], stage0_0[17], stage0_0[18]},
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[4]},
      {stage0_3[6]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[19], stage0_0[20], stage0_0[21]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[5]},
      {stage0_3[7]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[6]},
      {stage0_3[8]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29], stage0_0[30]},
      {stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35], stage0_0[36]},
      {stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60]},
      {stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66]},
      {stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72]},
      {stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78]},
      {stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84]},
      {stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96]},
      {stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102]},
      {stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[103], stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108]},
      {stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[109], stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114]},
      {stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[115], stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120]},
      {stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[121], stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126]},
      {stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[127], stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132]},
      {stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[133], stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138]},
      {stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[139], stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144]},
      {stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[145], stage0_0[146], stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150]},
      {stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[151], stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156]},
      {stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[157], stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162]},
      {stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[163], stage0_0[164], stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168]},
      {stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[169], stage0_0[170], stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174]},
      {stage0_2[151], stage0_2[152], stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[175], stage0_0[176], stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180]},
      {stage0_2[157], stage0_2[158], stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[181], stage0_0[182], stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186]},
      {stage0_2[163], stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[187], stage0_0[188], stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192]},
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198]},
      {stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204]},
      {stage0_2[181], stage0_2[182], stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210]},
      {stage0_2[187], stage0_2[188], stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214], stage0_0[215], stage0_0[216]},
      {stage0_2[193], stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220], stage0_0[221], stage0_0[222]},
      {stage0_2[199], stage0_2[200], stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226], stage0_0[227], stage0_0[228]},
      {stage0_2[205], stage0_2[206], stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232], stage0_0[233], stage0_0[234]},
      {stage0_2[211], stage0_2[212], stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238], stage0_0[239], stage0_0[240]},
      {stage0_2[217], stage0_2[218], stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244], stage0_0[245], stage0_0[246]},
      {stage0_2[223], stage0_2[224], stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250], stage0_0[251], stage0_0[252]},
      {stage0_2[229], stage0_2[230], stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[0],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[1],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[2],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[3],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38]},
      {stage1_5[4],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44]},
      {stage1_5[5],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50]},
      {stage1_5[6],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage1_5[7],stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62]},
      {stage1_5[8],stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68]},
      {stage1_5[9],stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74]},
      {stage1_5[10],stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80]},
      {stage1_5[11],stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage1_5[12],stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92]},
      {stage1_5[13],stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98]},
      {stage1_5[14],stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104]},
      {stage1_5[15],stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110]},
      {stage1_5[16],stage1_4[61],stage1_3[61],stage1_2[61],stage1_1[61]}
   );
   gpc606_5 gpc62 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage1_5[17],stage1_4[62],stage1_3[62],stage1_2[62],stage1_1[62]}
   );
   gpc606_5 gpc63 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122]},
      {stage1_5[18],stage1_4[63],stage1_3[63],stage1_2[63],stage1_1[63]}
   );
   gpc606_5 gpc64 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126], stage0_3[127], stage0_3[128]},
      {stage1_5[19],stage1_4[64],stage1_3[64],stage1_2[64],stage1_1[64]}
   );
   gpc606_5 gpc65 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132], stage0_3[133], stage0_3[134]},
      {stage1_5[20],stage1_4[65],stage1_3[65],stage1_2[65],stage1_1[65]}
   );
   gpc606_5 gpc66 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139], stage0_3[140]},
      {stage1_5[21],stage1_4[66],stage1_3[66],stage1_2[66],stage1_1[66]}
   );
   gpc606_5 gpc67 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144], stage0_3[145], stage0_3[146]},
      {stage1_5[22],stage1_4[67],stage1_3[67],stage1_2[67],stage1_1[67]}
   );
   gpc606_5 gpc68 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150], stage0_3[151], stage0_3[152]},
      {stage1_5[23],stage1_4[68],stage1_3[68],stage1_2[68],stage1_1[68]}
   );
   gpc606_5 gpc69 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158]},
      {stage1_5[24],stage1_4[69],stage1_3[69],stage1_2[69],stage1_1[69]}
   );
   gpc606_5 gpc70 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage1_5[25],stage1_4[70],stage1_3[70],stage1_2[70],stage1_1[70]}
   );
   gpc606_5 gpc71 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169], stage0_3[170]},
      {stage1_5[26],stage1_4[71],stage1_3[71],stage1_2[71],stage1_1[71]}
   );
   gpc606_5 gpc72 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174], stage0_3[175], stage0_3[176]},
      {stage1_5[27],stage1_4[72],stage1_3[72],stage1_2[72],stage1_1[72]}
   );
   gpc606_5 gpc73 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180], stage0_3[181], stage0_3[182]},
      {stage1_5[28],stage1_4[73],stage1_3[73],stage1_2[73],stage1_1[73]}
   );
   gpc606_5 gpc74 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188]},
      {stage1_5[29],stage1_4[74],stage1_3[74],stage1_2[74],stage1_1[74]}
   );
   gpc606_5 gpc75 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage1_5[30],stage1_4[75],stage1_3[75],stage1_2[75],stage1_1[75]}
   );
   gpc606_5 gpc76 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199], stage0_3[200]},
      {stage1_5[31],stage1_4[76],stage1_3[76],stage1_2[76],stage1_1[76]}
   );
   gpc606_5 gpc77 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204], stage0_3[205], stage0_3[206]},
      {stage1_5[32],stage1_4[77],stage1_3[77],stage1_2[77],stage1_1[77]}
   );
   gpc606_5 gpc78 (
      {stage0_1[234], stage0_1[235], stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239]},
      {stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210], stage0_3[211], stage0_3[212]},
      {stage1_5[33],stage1_4[78],stage1_3[78],stage1_2[78],stage1_1[78]}
   );
   gpc606_5 gpc79 (
      {stage0_1[240], stage0_1[241], stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245]},
      {stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218]},
      {stage1_5[34],stage1_4[79],stage1_3[79],stage1_2[79],stage1_1[79]}
   );
   gpc615_5 gpc80 (
      {stage0_2[235], stage0_2[236], stage0_2[237], stage0_2[238], stage0_2[239]},
      {stage0_3[219]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[35],stage1_4[80],stage1_3[80],stage1_2[80]}
   );
   gpc615_5 gpc81 (
      {stage0_2[240], stage0_2[241], stage0_2[242], stage0_2[243], stage0_2[244]},
      {stage0_3[220]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[36],stage1_4[81],stage1_3[81],stage1_2[81]}
   );
   gpc615_5 gpc82 (
      {stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248], stage0_2[249]},
      {stage0_3[221]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[37],stage1_4[82],stage1_3[82],stage1_2[82]}
   );
   gpc615_5 gpc83 (
      {stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage0_3[222]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[38],stage1_4[83],stage1_3[83],stage1_2[83]}
   );
   gpc615_5 gpc84 (
      {stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226], stage0_3[227]},
      {stage0_4[24]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[4],stage1_5[39],stage1_4[84],stage1_3[84]}
   );
   gpc615_5 gpc85 (
      {stage0_3[228], stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232]},
      {stage0_4[25]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[5],stage1_5[40],stage1_4[85],stage1_3[85]}
   );
   gpc615_5 gpc86 (
      {stage0_3[233], stage0_3[234], stage0_3[235], stage0_3[236], stage0_3[237]},
      {stage0_4[26]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[6],stage1_5[41],stage1_4[86],stage1_3[86]}
   );
   gpc615_5 gpc87 (
      {stage0_3[238], stage0_3[239], stage0_3[240], stage0_3[241], stage0_3[242]},
      {stage0_4[27]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[7],stage1_5[42],stage1_4[87],stage1_3[87]}
   );
   gpc615_5 gpc88 (
      {stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246], stage0_3[247]},
      {stage0_4[28]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[8],stage1_5[43],stage1_4[88],stage1_3[88]}
   );
   gpc606_5 gpc89 (
      {stage0_4[29], stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[5],stage1_6[9],stage1_5[44],stage1_4[89]}
   );
   gpc606_5 gpc90 (
      {stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[6],stage1_6[10],stage1_5[45],stage1_4[90]}
   );
   gpc606_5 gpc91 (
      {stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[7],stage1_6[11],stage1_5[46],stage1_4[91]}
   );
   gpc606_5 gpc92 (
      {stage0_4[47], stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[8],stage1_6[12],stage1_5[47],stage1_4[92]}
   );
   gpc606_5 gpc93 (
      {stage0_4[53], stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[9],stage1_6[13],stage1_5[48],stage1_4[93]}
   );
   gpc606_5 gpc94 (
      {stage0_4[59], stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[10],stage1_6[14],stage1_5[49],stage1_4[94]}
   );
   gpc606_5 gpc95 (
      {stage0_4[65], stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[11],stage1_6[15],stage1_5[50],stage1_4[95]}
   );
   gpc606_5 gpc96 (
      {stage0_4[71], stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[12],stage1_6[16],stage1_5[51],stage1_4[96]}
   );
   gpc606_5 gpc97 (
      {stage0_4[77], stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[13],stage1_6[17],stage1_5[52],stage1_4[97]}
   );
   gpc606_5 gpc98 (
      {stage0_4[83], stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[14],stage1_6[18],stage1_5[53],stage1_4[98]}
   );
   gpc606_5 gpc99 (
      {stage0_4[89], stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[15],stage1_6[19],stage1_5[54],stage1_4[99]}
   );
   gpc606_5 gpc100 (
      {stage0_4[95], stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[16],stage1_6[20],stage1_5[55],stage1_4[100]}
   );
   gpc606_5 gpc101 (
      {stage0_4[101], stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[17],stage1_6[21],stage1_5[56],stage1_4[101]}
   );
   gpc606_5 gpc102 (
      {stage0_4[107], stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[18],stage1_6[22],stage1_5[57],stage1_4[102]}
   );
   gpc606_5 gpc103 (
      {stage0_4[113], stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[19],stage1_6[23],stage1_5[58],stage1_4[103]}
   );
   gpc606_5 gpc104 (
      {stage0_4[119], stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[20],stage1_6[24],stage1_5[59],stage1_4[104]}
   );
   gpc606_5 gpc105 (
      {stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[21],stage1_6[25],stage1_5[60],stage1_4[105]}
   );
   gpc606_5 gpc106 (
      {stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[22],stage1_6[26],stage1_5[61],stage1_4[106]}
   );
   gpc606_5 gpc107 (
      {stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[23],stage1_6[27],stage1_5[62],stage1_4[107]}
   );
   gpc606_5 gpc108 (
      {stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[24],stage1_6[28],stage1_5[63],stage1_4[108]}
   );
   gpc606_5 gpc109 (
      {stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[25],stage1_6[29],stage1_5[64],stage1_4[109]}
   );
   gpc606_5 gpc110 (
      {stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[26],stage1_6[30],stage1_5[65],stage1_4[110]}
   );
   gpc606_5 gpc111 (
      {stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[27],stage1_6[31],stage1_5[66],stage1_4[111]}
   );
   gpc606_5 gpc112 (
      {stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[28],stage1_6[32],stage1_5[67],stage1_4[112]}
   );
   gpc606_5 gpc113 (
      {stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177], stage0_4[178]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[29],stage1_6[33],stage1_5[68],stage1_4[113]}
   );
   gpc606_5 gpc114 (
      {stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183], stage0_4[184]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[30],stage1_6[34],stage1_5[69],stage1_4[114]}
   );
   gpc606_5 gpc115 (
      {stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189], stage0_4[190]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[31],stage1_6[35],stage1_5[70],stage1_4[115]}
   );
   gpc606_5 gpc116 (
      {stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195], stage0_4[196]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[32],stage1_6[36],stage1_5[71],stage1_4[116]}
   );
   gpc606_5 gpc117 (
      {stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201], stage0_4[202]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[33],stage1_6[37],stage1_5[72],stage1_4[117]}
   );
   gpc606_5 gpc118 (
      {stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207], stage0_4[208]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[34],stage1_6[38],stage1_5[73],stage1_4[118]}
   );
   gpc606_5 gpc119 (
      {stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213], stage0_4[214]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[35],stage1_6[39],stage1_5[74],stage1_4[119]}
   );
   gpc606_5 gpc120 (
      {stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219], stage0_4[220]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[36],stage1_6[40],stage1_5[75],stage1_4[120]}
   );
   gpc606_5 gpc121 (
      {stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225], stage0_4[226]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[37],stage1_6[41],stage1_5[76],stage1_4[121]}
   );
   gpc606_5 gpc122 (
      {stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231], stage0_4[232]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[38],stage1_6[42],stage1_5[77],stage1_4[122]}
   );
   gpc606_5 gpc123 (
      {stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237], stage0_4[238]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[39],stage1_6[43],stage1_5[78],stage1_4[123]}
   );
   gpc606_5 gpc124 (
      {stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243], stage0_4[244]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[40],stage1_6[44],stage1_5[79],stage1_4[124]}
   );
   gpc606_5 gpc125 (
      {stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249], stage0_4[250]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[41],stage1_6[45],stage1_5[80],stage1_4[125]}
   );
   gpc615_5 gpc126 (
      {stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255]},
      {stage0_5[30]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[42],stage1_6[46],stage1_5[81],stage1_4[126]}
   );
   gpc606_5 gpc127 (
      {stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[38],stage1_7[43],stage1_6[47],stage1_5[82]}
   );
   gpc606_5 gpc128 (
      {stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[39],stage1_7[44],stage1_6[48],stage1_5[83]}
   );
   gpc606_5 gpc129 (
      {stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[40],stage1_7[45],stage1_6[49],stage1_5[84]}
   );
   gpc606_5 gpc130 (
      {stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[41],stage1_7[46],stage1_6[50],stage1_5[85]}
   );
   gpc606_5 gpc131 (
      {stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[42],stage1_7[47],stage1_6[51],stage1_5[86]}
   );
   gpc606_5 gpc132 (
      {stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[43],stage1_7[48],stage1_6[52],stage1_5[87]}
   );
   gpc606_5 gpc133 (
      {stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[44],stage1_7[49],stage1_6[53],stage1_5[88]}
   );
   gpc606_5 gpc134 (
      {stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[45],stage1_7[50],stage1_6[54],stage1_5[89]}
   );
   gpc606_5 gpc135 (
      {stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[46],stage1_7[51],stage1_6[55],stage1_5[90]}
   );
   gpc606_5 gpc136 (
      {stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[47],stage1_7[52],stage1_6[56],stage1_5[91]}
   );
   gpc606_5 gpc137 (
      {stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[48],stage1_7[53],stage1_6[57],stage1_5[92]}
   );
   gpc606_5 gpc138 (
      {stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[49],stage1_7[54],stage1_6[58],stage1_5[93]}
   );
   gpc606_5 gpc139 (
      {stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[50],stage1_7[55],stage1_6[59],stage1_5[94]}
   );
   gpc606_5 gpc140 (
      {stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[51],stage1_7[56],stage1_6[60],stage1_5[95]}
   );
   gpc606_5 gpc141 (
      {stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119], stage0_5[120]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[52],stage1_7[57],stage1_6[61],stage1_5[96]}
   );
   gpc606_5 gpc142 (
      {stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125], stage0_5[126]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[53],stage1_7[58],stage1_6[62],stage1_5[97]}
   );
   gpc606_5 gpc143 (
      {stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131], stage0_5[132]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[54],stage1_7[59],stage1_6[63],stage1_5[98]}
   );
   gpc606_5 gpc144 (
      {stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137], stage0_5[138]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[55],stage1_7[60],stage1_6[64],stage1_5[99]}
   );
   gpc606_5 gpc145 (
      {stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143], stage0_5[144]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[56],stage1_7[61],stage1_6[65],stage1_5[100]}
   );
   gpc606_5 gpc146 (
      {stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149], stage0_5[150]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[57],stage1_7[62],stage1_6[66],stage1_5[101]}
   );
   gpc606_5 gpc147 (
      {stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155], stage0_5[156]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[58],stage1_7[63],stage1_6[67],stage1_5[102]}
   );
   gpc606_5 gpc148 (
      {stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161], stage0_5[162]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[59],stage1_7[64],stage1_6[68],stage1_5[103]}
   );
   gpc606_5 gpc149 (
      {stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167], stage0_5[168]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[60],stage1_7[65],stage1_6[69],stage1_5[104]}
   );
   gpc606_5 gpc150 (
      {stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173], stage0_5[174]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[61],stage1_7[66],stage1_6[70],stage1_5[105]}
   );
   gpc606_5 gpc151 (
      {stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179], stage0_5[180]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[62],stage1_7[67],stage1_6[71],stage1_5[106]}
   );
   gpc606_5 gpc152 (
      {stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[63],stage1_7[68],stage1_6[72],stage1_5[107]}
   );
   gpc606_5 gpc153 (
      {stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[64],stage1_7[69],stage1_6[73],stage1_5[108]}
   );
   gpc606_5 gpc154 (
      {stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[65],stage1_7[70],stage1_6[74],stage1_5[109]}
   );
   gpc606_5 gpc155 (
      {stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[66],stage1_7[71],stage1_6[75],stage1_5[110]}
   );
   gpc606_5 gpc156 (
      {stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[67],stage1_7[72],stage1_6[76],stage1_5[111]}
   );
   gpc606_5 gpc157 (
      {stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[68],stage1_7[73],stage1_6[77],stage1_5[112]}
   );
   gpc606_5 gpc158 (
      {stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[69],stage1_7[74],stage1_6[78],stage1_5[113]}
   );
   gpc606_5 gpc159 (
      {stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[70],stage1_7[75],stage1_6[79],stage1_5[114]}
   );
   gpc606_5 gpc160 (
      {stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[71],stage1_7[76],stage1_6[80],stage1_5[115]}
   );
   gpc615_5 gpc161 (
      {stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_6[228]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[72],stage1_7[77],stage1_6[81],stage1_5[116]}
   );
   gpc615_5 gpc162 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244]},
      {stage0_6[229]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[73],stage1_7[78],stage1_6[82],stage1_5[117]}
   );
   gpc615_5 gpc163 (
      {stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233], stage0_6[234]},
      {stage0_7[216]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[36],stage1_8[74],stage1_7[79],stage1_6[83]}
   );
   gpc615_5 gpc164 (
      {stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage0_7[217]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[37],stage1_8[75],stage1_7[80],stage1_6[84]}
   );
   gpc615_5 gpc165 (
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244]},
      {stage0_7[218]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[38],stage1_8[76],stage1_7[81],stage1_6[85]}
   );
   gpc615_5 gpc166 (
      {stage0_6[245], stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249]},
      {stage0_7[219]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[39],stage1_8[77],stage1_7[82],stage1_6[86]}
   );
   gpc615_5 gpc167 (
      {stage0_6[250], stage0_6[251], stage0_6[252], stage0_6[253], stage0_6[254]},
      {stage0_7[220]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[40],stage1_8[78],stage1_7[83],stage1_6[87]}
   );
   gpc615_5 gpc168 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[30]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[5],stage1_9[41],stage1_8[79],stage1_7[84]}
   );
   gpc615_5 gpc169 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[31]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[6],stage1_9[42],stage1_8[80],stage1_7[85]}
   );
   gpc615_5 gpc170 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[32]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[7],stage1_9[43],stage1_8[81],stage1_7[86]}
   );
   gpc615_5 gpc171 (
      {stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239], stage0_7[240]},
      {stage0_8[33]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[8],stage1_9[44],stage1_8[82],stage1_7[87]}
   );
   gpc615_5 gpc172 (
      {stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage0_8[34]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[9],stage1_9[45],stage1_8[83],stage1_7[88]}
   );
   gpc615_5 gpc173 (
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250]},
      {stage0_8[35]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[10],stage1_9[46],stage1_8[84],stage1_7[89]}
   );
   gpc615_5 gpc174 (
      {stage0_7[251], stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255]},
      {stage0_8[36]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[11],stage1_9[47],stage1_8[85],stage1_7[90]}
   );
   gpc606_5 gpc175 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[7],stage1_10[12],stage1_9[48],stage1_8[86]}
   );
   gpc606_5 gpc176 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[8],stage1_10[13],stage1_9[49],stage1_8[87]}
   );
   gpc606_5 gpc177 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[9],stage1_10[14],stage1_9[50],stage1_8[88]}
   );
   gpc606_5 gpc178 (
      {stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[10],stage1_10[15],stage1_9[51],stage1_8[89]}
   );
   gpc606_5 gpc179 (
      {stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[11],stage1_10[16],stage1_9[52],stage1_8[90]}
   );
   gpc606_5 gpc180 (
      {stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[12],stage1_10[17],stage1_9[53],stage1_8[91]}
   );
   gpc606_5 gpc181 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[13],stage1_10[18],stage1_9[54],stage1_8[92]}
   );
   gpc606_5 gpc182 (
      {stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[14],stage1_10[19],stage1_9[55],stage1_8[93]}
   );
   gpc606_5 gpc183 (
      {stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[15],stage1_10[20],stage1_9[56],stage1_8[94]}
   );
   gpc606_5 gpc184 (
      {stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[16],stage1_10[21],stage1_9[57],stage1_8[95]}
   );
   gpc606_5 gpc185 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[17],stage1_10[22],stage1_9[58],stage1_8[96]}
   );
   gpc606_5 gpc186 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[18],stage1_10[23],stage1_9[59],stage1_8[97]}
   );
   gpc606_5 gpc187 (
      {stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[19],stage1_10[24],stage1_9[60],stage1_8[98]}
   );
   gpc606_5 gpc188 (
      {stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[20],stage1_10[25],stage1_9[61],stage1_8[99]}
   );
   gpc606_5 gpc189 (
      {stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[21],stage1_10[26],stage1_9[62],stage1_8[100]}
   );
   gpc606_5 gpc190 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[22],stage1_10[27],stage1_9[63],stage1_8[101]}
   );
   gpc606_5 gpc191 (
      {stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[23],stage1_10[28],stage1_9[64],stage1_8[102]}
   );
   gpc606_5 gpc192 (
      {stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[24],stage1_10[29],stage1_9[65],stage1_8[103]}
   );
   gpc606_5 gpc193 (
      {stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[25],stage1_10[30],stage1_9[66],stage1_8[104]}
   );
   gpc606_5 gpc194 (
      {stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[26],stage1_10[31],stage1_9[67],stage1_8[105]}
   );
   gpc606_5 gpc195 (
      {stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[27],stage1_10[32],stage1_9[68],stage1_8[106]}
   );
   gpc606_5 gpc196 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167], stage0_8[168]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[28],stage1_10[33],stage1_9[69],stage1_8[107]}
   );
   gpc606_5 gpc197 (
      {stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173], stage0_8[174]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[29],stage1_10[34],stage1_9[70],stage1_8[108]}
   );
   gpc606_5 gpc198 (
      {stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179], stage0_8[180]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[30],stage1_10[35],stage1_9[71],stage1_8[109]}
   );
   gpc606_5 gpc199 (
      {stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[31],stage1_10[36],stage1_9[72],stage1_8[110]}
   );
   gpc606_5 gpc200 (
      {stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[32],stage1_10[37],stage1_9[73],stage1_8[111]}
   );
   gpc606_5 gpc201 (
      {stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197], stage0_8[198]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[33],stage1_10[38],stage1_9[74],stage1_8[112]}
   );
   gpc606_5 gpc202 (
      {stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203], stage0_8[204]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[34],stage1_10[39],stage1_9[75],stage1_8[113]}
   );
   gpc606_5 gpc203 (
      {stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209], stage0_8[210]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[35],stage1_10[40],stage1_9[76],stage1_8[114]}
   );
   gpc606_5 gpc204 (
      {stage0_8[211], stage0_8[212], stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[36],stage1_10[41],stage1_9[77],stage1_8[115]}
   );
   gpc606_5 gpc205 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[30],stage1_11[37],stage1_10[42],stage1_9[78]}
   );
   gpc606_5 gpc206 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[31],stage1_11[38],stage1_10[43],stage1_9[79]}
   );
   gpc606_5 gpc207 (
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[32],stage1_11[39],stage1_10[44],stage1_9[80]}
   );
   gpc606_5 gpc208 (
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[33],stage1_11[40],stage1_10[45],stage1_9[81]}
   );
   gpc615_5 gpc209 (
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70]},
      {stage0_10[180]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[34],stage1_11[41],stage1_10[46],stage1_9[82]}
   );
   gpc615_5 gpc210 (
      {stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75]},
      {stage0_10[181]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[35],stage1_11[42],stage1_10[47],stage1_9[83]}
   );
   gpc615_5 gpc211 (
      {stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80]},
      {stage0_10[182]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[36],stage1_11[43],stage1_10[48],stage1_9[84]}
   );
   gpc615_5 gpc212 (
      {stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85]},
      {stage0_10[183]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[37],stage1_11[44],stage1_10[49],stage1_9[85]}
   );
   gpc615_5 gpc213 (
      {stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90]},
      {stage0_10[184]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[38],stage1_11[45],stage1_10[50],stage1_9[86]}
   );
   gpc615_5 gpc214 (
      {stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage0_10[185]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[39],stage1_11[46],stage1_10[51],stage1_9[87]}
   );
   gpc615_5 gpc215 (
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100]},
      {stage0_10[186]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[40],stage1_11[47],stage1_10[52],stage1_9[88]}
   );
   gpc615_5 gpc216 (
      {stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105]},
      {stage0_10[187]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[41],stage1_11[48],stage1_10[53],stage1_9[89]}
   );
   gpc615_5 gpc217 (
      {stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110]},
      {stage0_10[188]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[42],stage1_11[49],stage1_10[54],stage1_9[90]}
   );
   gpc615_5 gpc218 (
      {stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115]},
      {stage0_10[189]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[43],stage1_11[50],stage1_10[55],stage1_9[91]}
   );
   gpc615_5 gpc219 (
      {stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120]},
      {stage0_10[190]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[44],stage1_11[51],stage1_10[56],stage1_9[92]}
   );
   gpc615_5 gpc220 (
      {stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage0_10[191]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[45],stage1_11[52],stage1_10[57],stage1_9[93]}
   );
   gpc615_5 gpc221 (
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130]},
      {stage0_10[192]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[46],stage1_11[53],stage1_10[58],stage1_9[94]}
   );
   gpc615_5 gpc222 (
      {stage0_9[131], stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135]},
      {stage0_10[193]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[47],stage1_11[54],stage1_10[59],stage1_9[95]}
   );
   gpc615_5 gpc223 (
      {stage0_9[136], stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140]},
      {stage0_10[194]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[48],stage1_11[55],stage1_10[60],stage1_9[96]}
   );
   gpc615_5 gpc224 (
      {stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145]},
      {stage0_10[195]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[49],stage1_11[56],stage1_10[61],stage1_9[97]}
   );
   gpc615_5 gpc225 (
      {stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150]},
      {stage0_10[196]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[50],stage1_11[57],stage1_10[62],stage1_9[98]}
   );
   gpc615_5 gpc226 (
      {stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_10[197]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[51],stage1_11[58],stage1_10[63],stage1_9[99]}
   );
   gpc615_5 gpc227 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_10[198]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[52],stage1_11[59],stage1_10[64],stage1_9[100]}
   );
   gpc615_5 gpc228 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165]},
      {stage0_10[199]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[53],stage1_11[60],stage1_10[65],stage1_9[101]}
   );
   gpc615_5 gpc229 (
      {stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_10[200]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[54],stage1_11[61],stage1_10[66],stage1_9[102]}
   );
   gpc615_5 gpc230 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175]},
      {stage0_10[201]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[55],stage1_11[62],stage1_10[67],stage1_9[103]}
   );
   gpc615_5 gpc231 (
      {stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_10[202]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[56],stage1_11[63],stage1_10[68],stage1_9[104]}
   );
   gpc615_5 gpc232 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_10[203]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[57],stage1_11[64],stage1_10[69],stage1_9[105]}
   );
   gpc615_5 gpc233 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190]},
      {stage0_10[204]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[58],stage1_11[65],stage1_10[70],stage1_9[106]}
   );
   gpc615_5 gpc234 (
      {stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_10[205]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[59],stage1_11[66],stage1_10[71],stage1_9[107]}
   );
   gpc615_5 gpc235 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_10[206]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[60],stage1_11[67],stage1_10[72],stage1_9[108]}
   );
   gpc615_5 gpc236 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205]},
      {stage0_10[207]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[61],stage1_11[68],stage1_10[73],stage1_9[109]}
   );
   gpc615_5 gpc237 (
      {stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_10[208]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[62],stage1_11[69],stage1_10[74],stage1_9[110]}
   );
   gpc615_5 gpc238 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_10[209]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[63],stage1_11[70],stage1_10[75],stage1_9[111]}
   );
   gpc615_5 gpc239 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220]},
      {stage0_10[210]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[64],stage1_11[71],stage1_10[76],stage1_9[112]}
   );
   gpc615_5 gpc240 (
      {stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_10[211]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[65],stage1_11[72],stage1_10[77],stage1_9[113]}
   );
   gpc615_5 gpc241 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_10[212]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[66],stage1_11[73],stage1_10[78],stage1_9[114]}
   );
   gpc615_5 gpc242 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235]},
      {stage0_10[213]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[67],stage1_11[74],stage1_10[79],stage1_9[115]}
   );
   gpc615_5 gpc243 (
      {stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_10[214]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[68],stage1_11[75],stage1_10[80],stage1_9[116]}
   );
   gpc615_5 gpc244 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_10[215]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[69],stage1_11[76],stage1_10[81],stage1_9[117]}
   );
   gpc615_5 gpc245 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250]},
      {stage0_10[216]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[70],stage1_11[77],stage1_10[82],stage1_9[118]}
   );
   gpc615_5 gpc246 (
      {stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_10[217]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[71],stage1_11[78],stage1_10[83],stage1_9[119]}
   );
   gpc1_1 gpc247 (
      {stage0_0[253]},
      {stage1_0[45]}
   );
   gpc1_1 gpc248 (
      {stage0_0[254]},
      {stage1_0[46]}
   );
   gpc1_1 gpc249 (
      {stage0_0[255]},
      {stage1_0[47]}
   );
   gpc1_1 gpc250 (
      {stage0_1[246]},
      {stage1_1[80]}
   );
   gpc1_1 gpc251 (
      {stage0_1[247]},
      {stage1_1[81]}
   );
   gpc1_1 gpc252 (
      {stage0_1[248]},
      {stage1_1[82]}
   );
   gpc1_1 gpc253 (
      {stage0_1[249]},
      {stage1_1[83]}
   );
   gpc1_1 gpc254 (
      {stage0_1[250]},
      {stage1_1[84]}
   );
   gpc1_1 gpc255 (
      {stage0_1[251]},
      {stage1_1[85]}
   );
   gpc1_1 gpc256 (
      {stage0_1[252]},
      {stage1_1[86]}
   );
   gpc1_1 gpc257 (
      {stage0_1[253]},
      {stage1_1[87]}
   );
   gpc1_1 gpc258 (
      {stage0_1[254]},
      {stage1_1[88]}
   );
   gpc1_1 gpc259 (
      {stage0_1[255]},
      {stage1_1[89]}
   );
   gpc1_1 gpc260 (
      {stage0_2[255]},
      {stage1_2[84]}
   );
   gpc1_1 gpc261 (
      {stage0_3[248]},
      {stage1_3[89]}
   );
   gpc1_1 gpc262 (
      {stage0_3[249]},
      {stage1_3[90]}
   );
   gpc1_1 gpc263 (
      {stage0_3[250]},
      {stage1_3[91]}
   );
   gpc1_1 gpc264 (
      {stage0_3[251]},
      {stage1_3[92]}
   );
   gpc1_1 gpc265 (
      {stage0_3[252]},
      {stage1_3[93]}
   );
   gpc1_1 gpc266 (
      {stage0_3[253]},
      {stage1_3[94]}
   );
   gpc1_1 gpc267 (
      {stage0_3[254]},
      {stage1_3[95]}
   );
   gpc1_1 gpc268 (
      {stage0_3[255]},
      {stage1_3[96]}
   );
   gpc1_1 gpc269 (
      {stage0_5[245]},
      {stage1_5[118]}
   );
   gpc1_1 gpc270 (
      {stage0_5[246]},
      {stage1_5[119]}
   );
   gpc1_1 gpc271 (
      {stage0_5[247]},
      {stage1_5[120]}
   );
   gpc1_1 gpc272 (
      {stage0_5[248]},
      {stage1_5[121]}
   );
   gpc1_1 gpc273 (
      {stage0_5[249]},
      {stage1_5[122]}
   );
   gpc1_1 gpc274 (
      {stage0_5[250]},
      {stage1_5[123]}
   );
   gpc1_1 gpc275 (
      {stage0_5[251]},
      {stage1_5[124]}
   );
   gpc1_1 gpc276 (
      {stage0_5[252]},
      {stage1_5[125]}
   );
   gpc1_1 gpc277 (
      {stage0_5[253]},
      {stage1_5[126]}
   );
   gpc1_1 gpc278 (
      {stage0_5[254]},
      {stage1_5[127]}
   );
   gpc1_1 gpc279 (
      {stage0_5[255]},
      {stage1_5[128]}
   );
   gpc1_1 gpc280 (
      {stage0_6[255]},
      {stage1_6[88]}
   );
   gpc1_1 gpc281 (
      {stage0_8[217]},
      {stage1_8[116]}
   );
   gpc1_1 gpc282 (
      {stage0_8[218]},
      {stage1_8[117]}
   );
   gpc1_1 gpc283 (
      {stage0_8[219]},
      {stage1_8[118]}
   );
   gpc1_1 gpc284 (
      {stage0_8[220]},
      {stage1_8[119]}
   );
   gpc1_1 gpc285 (
      {stage0_8[221]},
      {stage1_8[120]}
   );
   gpc1_1 gpc286 (
      {stage0_8[222]},
      {stage1_8[121]}
   );
   gpc1_1 gpc287 (
      {stage0_8[223]},
      {stage1_8[122]}
   );
   gpc1_1 gpc288 (
      {stage0_8[224]},
      {stage1_8[123]}
   );
   gpc1_1 gpc289 (
      {stage0_8[225]},
      {stage1_8[124]}
   );
   gpc1_1 gpc290 (
      {stage0_8[226]},
      {stage1_8[125]}
   );
   gpc1_1 gpc291 (
      {stage0_8[227]},
      {stage1_8[126]}
   );
   gpc1_1 gpc292 (
      {stage0_8[228]},
      {stage1_8[127]}
   );
   gpc1_1 gpc293 (
      {stage0_8[229]},
      {stage1_8[128]}
   );
   gpc1_1 gpc294 (
      {stage0_8[230]},
      {stage1_8[129]}
   );
   gpc1_1 gpc295 (
      {stage0_8[231]},
      {stage1_8[130]}
   );
   gpc1_1 gpc296 (
      {stage0_8[232]},
      {stage1_8[131]}
   );
   gpc1_1 gpc297 (
      {stage0_8[233]},
      {stage1_8[132]}
   );
   gpc1_1 gpc298 (
      {stage0_8[234]},
      {stage1_8[133]}
   );
   gpc1_1 gpc299 (
      {stage0_8[235]},
      {stage1_8[134]}
   );
   gpc1_1 gpc300 (
      {stage0_8[236]},
      {stage1_8[135]}
   );
   gpc1_1 gpc301 (
      {stage0_8[237]},
      {stage1_8[136]}
   );
   gpc1_1 gpc302 (
      {stage0_8[238]},
      {stage1_8[137]}
   );
   gpc1_1 gpc303 (
      {stage0_8[239]},
      {stage1_8[138]}
   );
   gpc1_1 gpc304 (
      {stage0_8[240]},
      {stage1_8[139]}
   );
   gpc1_1 gpc305 (
      {stage0_8[241]},
      {stage1_8[140]}
   );
   gpc1_1 gpc306 (
      {stage0_8[242]},
      {stage1_8[141]}
   );
   gpc1_1 gpc307 (
      {stage0_8[243]},
      {stage1_8[142]}
   );
   gpc1_1 gpc308 (
      {stage0_8[244]},
      {stage1_8[143]}
   );
   gpc1_1 gpc309 (
      {stage0_8[245]},
      {stage1_8[144]}
   );
   gpc1_1 gpc310 (
      {stage0_8[246]},
      {stage1_8[145]}
   );
   gpc1_1 gpc311 (
      {stage0_8[247]},
      {stage1_8[146]}
   );
   gpc1_1 gpc312 (
      {stage0_8[248]},
      {stage1_8[147]}
   );
   gpc1_1 gpc313 (
      {stage0_8[249]},
      {stage1_8[148]}
   );
   gpc1_1 gpc314 (
      {stage0_8[250]},
      {stage1_8[149]}
   );
   gpc1_1 gpc315 (
      {stage0_8[251]},
      {stage1_8[150]}
   );
   gpc1_1 gpc316 (
      {stage0_8[252]},
      {stage1_8[151]}
   );
   gpc1_1 gpc317 (
      {stage0_8[253]},
      {stage1_8[152]}
   );
   gpc1_1 gpc318 (
      {stage0_8[254]},
      {stage1_8[153]}
   );
   gpc1_1 gpc319 (
      {stage0_8[255]},
      {stage1_8[154]}
   );
   gpc1_1 gpc320 (
      {stage0_10[218]},
      {stage1_10[84]}
   );
   gpc1_1 gpc321 (
      {stage0_10[219]},
      {stage1_10[85]}
   );
   gpc1_1 gpc322 (
      {stage0_10[220]},
      {stage1_10[86]}
   );
   gpc1_1 gpc323 (
      {stage0_10[221]},
      {stage1_10[87]}
   );
   gpc1_1 gpc324 (
      {stage0_10[222]},
      {stage1_10[88]}
   );
   gpc1_1 gpc325 (
      {stage0_10[223]},
      {stage1_10[89]}
   );
   gpc1_1 gpc326 (
      {stage0_10[224]},
      {stage1_10[90]}
   );
   gpc1_1 gpc327 (
      {stage0_10[225]},
      {stage1_10[91]}
   );
   gpc1_1 gpc328 (
      {stage0_10[226]},
      {stage1_10[92]}
   );
   gpc1_1 gpc329 (
      {stage0_10[227]},
      {stage1_10[93]}
   );
   gpc1_1 gpc330 (
      {stage0_10[228]},
      {stage1_10[94]}
   );
   gpc1_1 gpc331 (
      {stage0_10[229]},
      {stage1_10[95]}
   );
   gpc1_1 gpc332 (
      {stage0_10[230]},
      {stage1_10[96]}
   );
   gpc1_1 gpc333 (
      {stage0_10[231]},
      {stage1_10[97]}
   );
   gpc1_1 gpc334 (
      {stage0_10[232]},
      {stage1_10[98]}
   );
   gpc1_1 gpc335 (
      {stage0_10[233]},
      {stage1_10[99]}
   );
   gpc1_1 gpc336 (
      {stage0_10[234]},
      {stage1_10[100]}
   );
   gpc1_1 gpc337 (
      {stage0_10[235]},
      {stage1_10[101]}
   );
   gpc1_1 gpc338 (
      {stage0_10[236]},
      {stage1_10[102]}
   );
   gpc1_1 gpc339 (
      {stage0_10[237]},
      {stage1_10[103]}
   );
   gpc1_1 gpc340 (
      {stage0_10[238]},
      {stage1_10[104]}
   );
   gpc1_1 gpc341 (
      {stage0_10[239]},
      {stage1_10[105]}
   );
   gpc1_1 gpc342 (
      {stage0_10[240]},
      {stage1_10[106]}
   );
   gpc1_1 gpc343 (
      {stage0_10[241]},
      {stage1_10[107]}
   );
   gpc1_1 gpc344 (
      {stage0_10[242]},
      {stage1_10[108]}
   );
   gpc1_1 gpc345 (
      {stage0_10[243]},
      {stage1_10[109]}
   );
   gpc1_1 gpc346 (
      {stage0_10[244]},
      {stage1_10[110]}
   );
   gpc1_1 gpc347 (
      {stage0_10[245]},
      {stage1_10[111]}
   );
   gpc1_1 gpc348 (
      {stage0_10[246]},
      {stage1_10[112]}
   );
   gpc1_1 gpc349 (
      {stage0_10[247]},
      {stage1_10[113]}
   );
   gpc1_1 gpc350 (
      {stage0_10[248]},
      {stage1_10[114]}
   );
   gpc1_1 gpc351 (
      {stage0_10[249]},
      {stage1_10[115]}
   );
   gpc1_1 gpc352 (
      {stage0_10[250]},
      {stage1_10[116]}
   );
   gpc1_1 gpc353 (
      {stage0_10[251]},
      {stage1_10[117]}
   );
   gpc1_1 gpc354 (
      {stage0_10[252]},
      {stage1_10[118]}
   );
   gpc1_1 gpc355 (
      {stage0_10[253]},
      {stage1_10[119]}
   );
   gpc1_1 gpc356 (
      {stage0_10[254]},
      {stage1_10[120]}
   );
   gpc1_1 gpc357 (
      {stage0_10[255]},
      {stage1_10[121]}
   );
   gpc1_1 gpc358 (
      {stage0_11[252]},
      {stage1_11[79]}
   );
   gpc1_1 gpc359 (
      {stage0_11[253]},
      {stage1_11[80]}
   );
   gpc1_1 gpc360 (
      {stage0_11[254]},
      {stage1_11[81]}
   );
   gpc1_1 gpc361 (
      {stage0_11[255]},
      {stage1_11[82]}
   );
   gpc1163_5 gpc362 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc363 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc364 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc365 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc366 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc367 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc368 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc369 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc370 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc371 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc372 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc373 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc374 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc7_3 gpc375 (
      {stage1_1[72], stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77], stage1_1[78]},
      {stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc376 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[0],stage2_4[13],stage2_3[14],stage2_2[14]}
   );
   gpc606_5 gpc377 (
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[1],stage2_4[14],stage2_3[15],stage2_2[15]}
   );
   gpc606_5 gpc378 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[2],stage2_4[15],stage2_3[16],stage2_2[16]}
   );
   gpc606_5 gpc379 (
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[3],stage2_4[16],stage2_3[17],stage2_2[17]}
   );
   gpc606_5 gpc380 (
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[4],stage2_4[17],stage2_3[18],stage2_2[18]}
   );
   gpc606_5 gpc381 (
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[5],stage2_4[18],stage2_3[19],stage2_2[19]}
   );
   gpc606_5 gpc382 (
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[6],stage2_4[19],stage2_3[20],stage2_2[20]}
   );
   gpc606_5 gpc383 (
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[7],stage2_4[20],stage2_3[21],stage2_2[21]}
   );
   gpc606_5 gpc384 (
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[8],stage2_4[21],stage2_3[22],stage2_2[22]}
   );
   gpc606_5 gpc385 (
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[9],stage2_4[22],stage2_3[23],stage2_2[23]}
   );
   gpc606_5 gpc386 (
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82], stage1_2[83]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[10],stage2_4[23],stage2_3[24],stage2_2[24]}
   );
   gpc615_5 gpc387 (
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16]},
      {stage1_4[66]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[11],stage2_5[11],stage2_4[24],stage2_3[25]}
   );
   gpc615_5 gpc388 (
      {stage1_3[17], stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[67]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[12],stage2_5[12],stage2_4[25],stage2_3[26]}
   );
   gpc615_5 gpc389 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26]},
      {stage1_4[68]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[13],stage2_5[13],stage2_4[26],stage2_3[27]}
   );
   gpc615_5 gpc390 (
      {stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage1_4[69]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[14],stage2_5[14],stage2_4[27],stage2_3[28]}
   );
   gpc615_5 gpc391 (
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36]},
      {stage1_4[70]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[15],stage2_5[15],stage2_4[28],stage2_3[29]}
   );
   gpc615_5 gpc392 (
      {stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage1_4[71]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[16],stage2_5[16],stage2_4[29],stage2_3[30]}
   );
   gpc615_5 gpc393 (
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46]},
      {stage1_4[72]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[17],stage2_5[17],stage2_4[30],stage2_3[31]}
   );
   gpc615_5 gpc394 (
      {stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51]},
      {stage1_4[73]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[18],stage2_5[18],stage2_4[31],stage2_3[32]}
   );
   gpc615_5 gpc395 (
      {stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55], stage1_3[56]},
      {stage1_4[74]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[19],stage2_5[19],stage2_4[32],stage2_3[33]}
   );
   gpc615_5 gpc396 (
      {stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage1_4[75]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[20],stage2_5[20],stage2_4[33],stage2_3[34]}
   );
   gpc615_5 gpc397 (
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66]},
      {stage1_4[76]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[21],stage2_5[21],stage2_4[34],stage2_3[35]}
   );
   gpc615_5 gpc398 (
      {stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage1_4[77]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[22],stage2_5[22],stage2_4[35],stage2_3[36]}
   );
   gpc615_5 gpc399 (
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76]},
      {stage1_4[78]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[23],stage2_5[23],stage2_4[36],stage2_3[37]}
   );
   gpc615_5 gpc400 (
      {stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81]},
      {stage1_4[79]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[24],stage2_5[24],stage2_4[37],stage2_3[38]}
   );
   gpc615_5 gpc401 (
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86]},
      {stage1_4[80]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[25],stage2_5[25],stage2_4[38],stage2_3[39]}
   );
   gpc615_5 gpc402 (
      {stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91]},
      {stage1_4[81]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[26],stage2_5[26],stage2_4[39],stage2_3[40]}
   );
   gpc615_5 gpc403 (
      {stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95], stage1_3[96]},
      {stage1_4[82]},
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage2_7[16],stage2_6[27],stage2_5[27],stage2_4[40],stage2_3[41]}
   );
   gpc606_5 gpc404 (
      {stage1_4[83], stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[17],stage2_6[28],stage2_5[28],stage2_4[41]}
   );
   gpc606_5 gpc405 (
      {stage1_4[89], stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[18],stage2_6[29],stage2_5[29],stage2_4[42]}
   );
   gpc606_5 gpc406 (
      {stage1_4[95], stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[19],stage2_6[30],stage2_5[30],stage2_4[43]}
   );
   gpc606_5 gpc407 (
      {stage1_4[101], stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[20],stage2_6[31],stage2_5[31],stage2_4[44]}
   );
   gpc606_5 gpc408 (
      {stage1_4[107], stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[21],stage2_6[32],stage2_5[32],stage2_4[45]}
   );
   gpc606_5 gpc409 (
      {stage1_4[113], stage1_4[114], stage1_4[115], stage1_4[116], stage1_4[117], stage1_4[118]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[22],stage2_6[33],stage2_5[33],stage2_4[46]}
   );
   gpc606_5 gpc410 (
      {stage1_4[119], stage1_4[120], stage1_4[121], stage1_4[122], stage1_4[123], stage1_4[124]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[23],stage2_6[34],stage2_5[34],stage2_4[47]}
   );
   gpc606_5 gpc411 (
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[7],stage2_7[24],stage2_6[35],stage2_5[35]}
   );
   gpc606_5 gpc412 (
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[8],stage2_7[25],stage2_6[36],stage2_5[36]}
   );
   gpc606_5 gpc413 (
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[9],stage2_7[26],stage2_6[37],stage2_5[37]}
   );
   gpc606_5 gpc414 (
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[10],stage2_7[27],stage2_6[38],stage2_5[38]}
   );
   gpc615_5 gpc415 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46]},
      {stage1_7[24]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[4],stage2_8[11],stage2_7[28],stage2_6[39]}
   );
   gpc615_5 gpc416 (
      {stage1_6[47], stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51]},
      {stage1_7[25]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[5],stage2_8[12],stage2_7[29],stage2_6[40]}
   );
   gpc615_5 gpc417 (
      {stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55], stage1_6[56]},
      {stage1_7[26]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[6],stage2_8[13],stage2_7[30],stage2_6[41]}
   );
   gpc615_5 gpc418 (
      {stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60], stage1_6[61]},
      {stage1_7[27]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[7],stage2_8[14],stage2_7[31],stage2_6[42]}
   );
   gpc615_5 gpc419 (
      {stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65], stage1_6[66]},
      {stage1_7[28]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[8],stage2_8[15],stage2_7[32],stage2_6[43]}
   );
   gpc615_5 gpc420 (
      {stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage1_7[29]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[9],stage2_8[16],stage2_7[33],stage2_6[44]}
   );
   gpc615_5 gpc421 (
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76]},
      {stage1_7[30]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[10],stage2_8[17],stage2_7[34],stage2_6[45]}
   );
   gpc615_5 gpc422 (
      {stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81]},
      {stage1_7[31]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[11],stage2_8[18],stage2_7[35],stage2_6[46]}
   );
   gpc615_5 gpc423 (
      {stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36]},
      {stage1_8[48]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[8],stage2_9[12],stage2_8[19],stage2_7[36]}
   );
   gpc615_5 gpc424 (
      {stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage1_8[49]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[9],stage2_9[13],stage2_8[20],stage2_7[37]}
   );
   gpc615_5 gpc425 (
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46]},
      {stage1_8[50]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[10],stage2_9[14],stage2_8[21],stage2_7[38]}
   );
   gpc615_5 gpc426 (
      {stage1_7[47], stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51]},
      {stage1_8[51]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[11],stage2_9[15],stage2_8[22],stage2_7[39]}
   );
   gpc615_5 gpc427 (
      {stage1_7[52], stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56]},
      {stage1_8[52]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[12],stage2_9[16],stage2_8[23],stage2_7[40]}
   );
   gpc615_5 gpc428 (
      {stage1_7[57], stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61]},
      {stage1_8[53]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[13],stage2_9[17],stage2_8[24],stage2_7[41]}
   );
   gpc615_5 gpc429 (
      {stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66]},
      {stage1_8[54]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[14],stage2_9[18],stage2_8[25],stage2_7[42]}
   );
   gpc615_5 gpc430 (
      {stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage1_8[55]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[15],stage2_9[19],stage2_8[26],stage2_7[43]}
   );
   gpc615_5 gpc431 (
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76]},
      {stage1_8[56]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[16],stage2_9[20],stage2_8[27],stage2_7[44]}
   );
   gpc615_5 gpc432 (
      {stage1_7[77], stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81]},
      {stage1_8[57]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[17],stage2_9[21],stage2_8[28],stage2_7[45]}
   );
   gpc615_5 gpc433 (
      {stage1_7[82], stage1_7[83], stage1_7[84], stage1_7[85], stage1_7[86]},
      {stage1_8[58]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[18],stage2_9[22],stage2_8[29],stage2_7[46]}
   );
   gpc615_5 gpc434 (
      {stage1_7[87], stage1_7[88], stage1_7[89], stage1_7[90], 1'b0},
      {stage1_8[59]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[19],stage2_9[23],stage2_8[30],stage2_7[47]}
   );
   gpc606_5 gpc435 (
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[12],stage2_10[20],stage2_9[24],stage2_8[31]}
   );
   gpc606_5 gpc436 (
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[13],stage2_10[21],stage2_9[25],stage2_8[32]}
   );
   gpc606_5 gpc437 (
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[14],stage2_10[22],stage2_9[26],stage2_8[33]}
   );
   gpc606_5 gpc438 (
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[15],stage2_10[23],stage2_9[27],stage2_8[34]}
   );
   gpc606_5 gpc439 (
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[16],stage2_10[24],stage2_9[28],stage2_8[35]}
   );
   gpc606_5 gpc440 (
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[17],stage2_10[25],stage2_9[29],stage2_8[36]}
   );
   gpc606_5 gpc441 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[18],stage2_10[26],stage2_9[30],stage2_8[37]}
   );
   gpc606_5 gpc442 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[19],stage2_10[27],stage2_9[31],stage2_8[38]}
   );
   gpc606_5 gpc443 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[20],stage2_10[28],stage2_9[32],stage2_8[39]}
   );
   gpc606_5 gpc444 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[21],stage2_10[29],stage2_9[33],stage2_8[40]}
   );
   gpc606_5 gpc445 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[22],stage2_10[30],stage2_9[34],stage2_8[41]}
   );
   gpc606_5 gpc446 (
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[11],stage2_11[23],stage2_10[31],stage2_9[35]}
   );
   gpc606_5 gpc447 (
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[12],stage2_11[24],stage2_10[32],stage2_9[36]}
   );
   gpc606_5 gpc448 (
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[13],stage2_11[25],stage2_10[33],stage2_9[37]}
   );
   gpc606_5 gpc449 (
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[14],stage2_11[26],stage2_10[34],stage2_9[38]}
   );
   gpc606_5 gpc450 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[15],stage2_11[27],stage2_10[35],stage2_9[39]}
   );
   gpc606_5 gpc451 (
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[16],stage2_11[28],stage2_10[36],stage2_9[40]}
   );
   gpc606_5 gpc452 (
      {stage1_9[108], stage1_9[109], stage1_9[110], stage1_9[111], stage1_9[112], stage1_9[113]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[17],stage2_11[29],stage2_10[37],stage2_9[41]}
   );
   gpc606_5 gpc453 (
      {stage1_9[114], stage1_9[115], stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[18],stage2_11[30],stage2_10[38],stage2_9[42]}
   );
   gpc606_5 gpc454 (
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[8],stage2_12[19],stage2_11[31],stage2_10[39]}
   );
   gpc615_5 gpc455 (
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76]},
      {stage1_11[48]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[9],stage2_12[20],stage2_11[32],stage2_10[40]}
   );
   gpc615_5 gpc456 (
      {stage1_10[77], stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81]},
      {stage1_11[49]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[10],stage2_12[21],stage2_11[33],stage2_10[41]}
   );
   gpc615_5 gpc457 (
      {stage1_10[82], stage1_10[83], stage1_10[84], stage1_10[85], stage1_10[86]},
      {stage1_11[50]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[11],stage2_12[22],stage2_11[34],stage2_10[42]}
   );
   gpc615_5 gpc458 (
      {stage1_10[87], stage1_10[88], stage1_10[89], stage1_10[90], stage1_10[91]},
      {stage1_11[51]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[12],stage2_12[23],stage2_11[35],stage2_10[43]}
   );
   gpc615_5 gpc459 (
      {stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95], stage1_10[96]},
      {stage1_11[52]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[13],stage2_12[24],stage2_11[36],stage2_10[44]}
   );
   gpc615_5 gpc460 (
      {stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage1_11[53]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[14],stage2_12[25],stage2_11[37],stage2_10[45]}
   );
   gpc615_5 gpc461 (
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_11[54]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[15],stage2_12[26],stage2_11[38],stage2_10[46]}
   );
   gpc615_5 gpc462 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111]},
      {stage1_11[55]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[16],stage2_12[27],stage2_11[39],stage2_10[47]}
   );
   gpc615_5 gpc463 (
      {stage1_10[112], stage1_10[113], stage1_10[114], stage1_10[115], stage1_10[116]},
      {stage1_11[56]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[17],stage2_12[28],stage2_11[40],stage2_10[48]}
   );
   gpc615_5 gpc464 (
      {stage1_10[117], stage1_10[118], stage1_10[119], stage1_10[120], stage1_10[121]},
      {stage1_11[57]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[18],stage2_12[29],stage2_11[41],stage2_10[49]}
   );
   gpc615_5 gpc465 (
      {stage1_11[58], stage1_11[59], stage1_11[60], stage1_11[61], stage1_11[62]},
      {stage1_12[66]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[11],stage2_13[19],stage2_12[30],stage2_11[42]}
   );
   gpc615_5 gpc466 (
      {stage1_11[63], stage1_11[64], stage1_11[65], stage1_11[66], stage1_11[67]},
      {stage1_12[67]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[12],stage2_13[20],stage2_12[31],stage2_11[43]}
   );
   gpc615_5 gpc467 (
      {stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71], stage1_11[72]},
      {stage1_12[68]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[13],stage2_13[21],stage2_12[32],stage2_11[44]}
   );
   gpc615_5 gpc468 (
      {stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage1_12[69]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[14],stage2_13[22],stage2_12[33],stage2_11[45]}
   );
   gpc615_5 gpc469 (
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82]},
      {stage1_12[70]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[15],stage2_13[23],stage2_12[34],stage2_11[46]}
   );
   gpc1_1 gpc470 (
      {stage1_0[42]},
      {stage2_0[13]}
   );
   gpc1_1 gpc471 (
      {stage1_0[43]},
      {stage2_0[14]}
   );
   gpc1_1 gpc472 (
      {stage1_0[44]},
      {stage2_0[15]}
   );
   gpc1_1 gpc473 (
      {stage1_0[45]},
      {stage2_0[16]}
   );
   gpc1_1 gpc474 (
      {stage1_0[46]},
      {stage2_0[17]}
   );
   gpc1_1 gpc475 (
      {stage1_0[47]},
      {stage2_0[18]}
   );
   gpc1_1 gpc476 (
      {stage1_1[79]},
      {stage2_1[14]}
   );
   gpc1_1 gpc477 (
      {stage1_1[80]},
      {stage2_1[15]}
   );
   gpc1_1 gpc478 (
      {stage1_1[81]},
      {stage2_1[16]}
   );
   gpc1_1 gpc479 (
      {stage1_1[82]},
      {stage2_1[17]}
   );
   gpc1_1 gpc480 (
      {stage1_1[83]},
      {stage2_1[18]}
   );
   gpc1_1 gpc481 (
      {stage1_1[84]},
      {stage2_1[19]}
   );
   gpc1_1 gpc482 (
      {stage1_1[85]},
      {stage2_1[20]}
   );
   gpc1_1 gpc483 (
      {stage1_1[86]},
      {stage2_1[21]}
   );
   gpc1_1 gpc484 (
      {stage1_1[87]},
      {stage2_1[22]}
   );
   gpc1_1 gpc485 (
      {stage1_1[88]},
      {stage2_1[23]}
   );
   gpc1_1 gpc486 (
      {stage1_1[89]},
      {stage2_1[24]}
   );
   gpc1_1 gpc487 (
      {stage1_2[84]},
      {stage2_2[25]}
   );
   gpc1_1 gpc488 (
      {stage1_4[125]},
      {stage2_4[48]}
   );
   gpc1_1 gpc489 (
      {stage1_4[126]},
      {stage2_4[49]}
   );
   gpc1_1 gpc490 (
      {stage1_5[126]},
      {stage2_5[39]}
   );
   gpc1_1 gpc491 (
      {stage1_5[127]},
      {stage2_5[40]}
   );
   gpc1_1 gpc492 (
      {stage1_5[128]},
      {stage2_5[41]}
   );
   gpc1_1 gpc493 (
      {stage1_6[82]},
      {stage2_6[47]}
   );
   gpc1_1 gpc494 (
      {stage1_6[83]},
      {stage2_6[48]}
   );
   gpc1_1 gpc495 (
      {stage1_6[84]},
      {stage2_6[49]}
   );
   gpc1_1 gpc496 (
      {stage1_6[85]},
      {stage2_6[50]}
   );
   gpc1_1 gpc497 (
      {stage1_6[86]},
      {stage2_6[51]}
   );
   gpc1_1 gpc498 (
      {stage1_6[87]},
      {stage2_6[52]}
   );
   gpc1_1 gpc499 (
      {stage1_6[88]},
      {stage2_6[53]}
   );
   gpc1_1 gpc500 (
      {stage1_8[126]},
      {stage2_8[42]}
   );
   gpc1_1 gpc501 (
      {stage1_8[127]},
      {stage2_8[43]}
   );
   gpc1_1 gpc502 (
      {stage1_8[128]},
      {stage2_8[44]}
   );
   gpc1_1 gpc503 (
      {stage1_8[129]},
      {stage2_8[45]}
   );
   gpc1_1 gpc504 (
      {stage1_8[130]},
      {stage2_8[46]}
   );
   gpc1_1 gpc505 (
      {stage1_8[131]},
      {stage2_8[47]}
   );
   gpc1_1 gpc506 (
      {stage1_8[132]},
      {stage2_8[48]}
   );
   gpc1_1 gpc507 (
      {stage1_8[133]},
      {stage2_8[49]}
   );
   gpc1_1 gpc508 (
      {stage1_8[134]},
      {stage2_8[50]}
   );
   gpc1_1 gpc509 (
      {stage1_8[135]},
      {stage2_8[51]}
   );
   gpc1_1 gpc510 (
      {stage1_8[136]},
      {stage2_8[52]}
   );
   gpc1_1 gpc511 (
      {stage1_8[137]},
      {stage2_8[53]}
   );
   gpc1_1 gpc512 (
      {stage1_8[138]},
      {stage2_8[54]}
   );
   gpc1_1 gpc513 (
      {stage1_8[139]},
      {stage2_8[55]}
   );
   gpc1_1 gpc514 (
      {stage1_8[140]},
      {stage2_8[56]}
   );
   gpc1_1 gpc515 (
      {stage1_8[141]},
      {stage2_8[57]}
   );
   gpc1_1 gpc516 (
      {stage1_8[142]},
      {stage2_8[58]}
   );
   gpc1_1 gpc517 (
      {stage1_8[143]},
      {stage2_8[59]}
   );
   gpc1_1 gpc518 (
      {stage1_8[144]},
      {stage2_8[60]}
   );
   gpc1_1 gpc519 (
      {stage1_8[145]},
      {stage2_8[61]}
   );
   gpc1_1 gpc520 (
      {stage1_8[146]},
      {stage2_8[62]}
   );
   gpc1_1 gpc521 (
      {stage1_8[147]},
      {stage2_8[63]}
   );
   gpc1_1 gpc522 (
      {stage1_8[148]},
      {stage2_8[64]}
   );
   gpc1_1 gpc523 (
      {stage1_8[149]},
      {stage2_8[65]}
   );
   gpc1_1 gpc524 (
      {stage1_8[150]},
      {stage2_8[66]}
   );
   gpc1_1 gpc525 (
      {stage1_8[151]},
      {stage2_8[67]}
   );
   gpc1_1 gpc526 (
      {stage1_8[152]},
      {stage2_8[68]}
   );
   gpc1_1 gpc527 (
      {stage1_8[153]},
      {stage2_8[69]}
   );
   gpc1_1 gpc528 (
      {stage1_8[154]},
      {stage2_8[70]}
   );
   gpc1_1 gpc529 (
      {stage1_12[71]},
      {stage2_12[35]}
   );
   gpc1_1 gpc530 (
      {stage1_13[30]},
      {stage2_13[24]}
   );
   gpc1_1 gpc531 (
      {stage1_13[31]},
      {stage2_13[25]}
   );
   gpc1_1 gpc532 (
      {stage1_13[32]},
      {stage2_13[26]}
   );
   gpc1_1 gpc533 (
      {stage1_13[33]},
      {stage2_13[27]}
   );
   gpc1_1 gpc534 (
      {stage1_13[34]},
      {stage2_13[28]}
   );
   gpc1_1 gpc535 (
      {stage1_13[35]},
      {stage2_13[29]}
   );
   gpc1_1 gpc536 (
      {stage1_13[36]},
      {stage2_13[30]}
   );
   gpc1_1 gpc537 (
      {stage1_13[37]},
      {stage2_13[31]}
   );
   gpc1_1 gpc538 (
      {stage1_13[38]},
      {stage2_13[32]}
   );
   gpc1_1 gpc539 (
      {stage1_13[39]},
      {stage2_13[33]}
   );
   gpc1_1 gpc540 (
      {stage1_13[40]},
      {stage2_13[34]}
   );
   gpc1_1 gpc541 (
      {stage1_13[41]},
      {stage2_13[35]}
   );
   gpc606_5 gpc542 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc543 (
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc606_5 gpc544 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[2],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc545 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[3],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc546 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[4],stage3_4[4],stage3_3[4],stage3_2[4]}
   );
   gpc615_5 gpc547 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10]},
      {stage2_3[24]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[5],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc615_5 gpc548 (
      {stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15]},
      {stage2_3[25]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[6],stage3_4[6],stage3_3[6],stage3_2[6]}
   );
   gpc615_5 gpc549 (
      {stage2_2[16], stage2_2[17], stage2_2[18], stage2_2[19], stage2_2[20]},
      {stage2_3[26]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[7],stage3_4[7],stage3_3[7],stage3_2[7]}
   );
   gpc615_5 gpc550 (
      {stage2_3[27], stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31]},
      {stage2_4[24]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[4],stage3_5[8],stage3_4[8],stage3_3[8]}
   );
   gpc615_5 gpc551 (
      {stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35], stage2_3[36]},
      {stage2_4[25]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[5],stage3_5[9],stage3_4[9],stage3_3[9]}
   );
   gpc615_5 gpc552 (
      {stage2_3[37], stage2_3[38], stage2_3[39], stage2_3[40], stage2_3[41]},
      {stage2_4[26]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[6],stage3_5[10],stage3_4[10],stage3_3[10]}
   );
   gpc606_5 gpc553 (
      {stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31], stage2_4[32]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[3],stage3_6[7],stage3_5[11],stage3_4[11]}
   );
   gpc606_5 gpc554 (
      {stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37], stage2_4[38]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[4],stage3_6[8],stage3_5[12],stage3_4[12]}
   );
   gpc606_5 gpc555 (
      {stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42], stage2_4[43], stage2_4[44]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[5],stage3_6[9],stage3_5[13],stage3_4[13]}
   );
   gpc606_5 gpc556 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[3],stage3_7[6],stage3_6[10],stage3_5[14]}
   );
   gpc606_5 gpc557 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[4],stage3_7[7],stage3_6[11],stage3_5[15]}
   );
   gpc606_5 gpc558 (
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[5],stage3_7[8],stage3_6[12],stage3_5[16]}
   );
   gpc606_5 gpc559 (
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage3_9[3],stage3_8[6],stage3_7[9],stage3_6[13],stage3_5[17]}
   );
   gpc606_5 gpc560 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[4],stage3_8[7],stage3_7[10],stage3_6[14]}
   );
   gpc606_5 gpc561 (
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[5],stage3_8[8],stage3_7[11],stage3_6[15]}
   );
   gpc606_5 gpc562 (
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[6],stage3_8[9],stage3_7[12],stage3_6[16]}
   );
   gpc615_5 gpc563 (
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40]},
      {stage2_7[24]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[7],stage3_8[10],stage3_7[13],stage3_6[17]}
   );
   gpc615_5 gpc564 (
      {stage2_6[41], stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45]},
      {stage2_7[25]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[8],stage3_8[11],stage3_7[14],stage3_6[18]}
   );
   gpc615_5 gpc565 (
      {stage2_6[46], stage2_6[47], stage2_6[48], stage2_6[49], stage2_6[50]},
      {stage2_7[26]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[9],stage3_8[12],stage3_7[15],stage3_6[19]}
   );
   gpc615_5 gpc566 (
      {stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage2_8[36]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[6],stage3_9[10],stage3_8[13],stage3_7[16]}
   );
   gpc615_5 gpc567 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[37]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[7],stage3_9[11],stage3_8[14],stage3_7[17]}
   );
   gpc615_5 gpc568 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[38]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[8],stage3_9[12],stage3_8[15],stage3_7[18]}
   );
   gpc615_5 gpc569 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[39]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[9],stage3_9[13],stage3_8[16],stage3_7[19]}
   );
   gpc615_5 gpc570 (
      {stage2_8[40], stage2_8[41], stage2_8[42], stage2_8[43], stage2_8[44]},
      {stage2_9[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[10],stage3_9[14],stage3_8[17]}
   );
   gpc615_5 gpc571 (
      {stage2_8[45], stage2_8[46], stage2_8[47], stage2_8[48], stage2_8[49]},
      {stage2_9[25]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[11],stage3_9[15],stage3_8[18]}
   );
   gpc615_5 gpc572 (
      {stage2_8[50], stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54]},
      {stage2_9[26]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[12],stage3_9[16],stage3_8[19]}
   );
   gpc615_5 gpc573 (
      {stage2_8[55], stage2_8[56], stage2_8[57], stage2_8[58], stage2_8[59]},
      {stage2_9[27]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[7],stage3_10[13],stage3_9[17],stage3_8[20]}
   );
   gpc615_5 gpc574 (
      {stage2_8[60], stage2_8[61], stage2_8[62], stage2_8[63], stage2_8[64]},
      {stage2_9[28]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[8],stage3_10[14],stage3_9[18],stage3_8[21]}
   );
   gpc615_5 gpc575 (
      {stage2_8[65], stage2_8[66], stage2_8[67], stage2_8[68], stage2_8[69]},
      {stage2_9[29]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[9],stage3_10[15],stage3_9[19],stage3_8[22]}
   );
   gpc606_5 gpc576 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[6],stage3_11[10],stage3_10[16],stage3_9[20]}
   );
   gpc615_5 gpc577 (
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40]},
      {stage2_11[6]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[7],stage3_11[11],stage3_10[17]}
   );
   gpc615_5 gpc578 (
      {stage2_10[41], stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45]},
      {stage2_11[7]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[2],stage3_12[8],stage3_11[12],stage3_10[18]}
   );
   gpc615_5 gpc579 (
      {stage2_10[46], stage2_10[47], stage2_10[48], stage2_10[49], 1'b0},
      {stage2_11[8]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[3],stage3_12[9],stage3_11[13],stage3_10[19]}
   );
   gpc606_5 gpc580 (
      {stage2_11[9], stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[4],stage3_12[10],stage3_11[14]}
   );
   gpc606_5 gpc581 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[5],stage3_12[11],stage3_11[15]}
   );
   gpc606_5 gpc582 (
      {stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[6],stage3_12[12],stage3_11[16]}
   );
   gpc606_5 gpc583 (
      {stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[6],stage3_13[7],stage3_12[13],stage3_11[17]}
   );
   gpc606_5 gpc584 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[7],stage3_13[8],stage3_12[14],stage3_11[18]}
   );
   gpc606_5 gpc585 (
      {stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[8],stage3_13[9],stage3_12[15],stage3_11[19]}
   );
   gpc1406_5 gpc586 (
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[6],stage3_14[9],stage3_13[10],stage3_12[16]}
   );
   gpc606_5 gpc587 (
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage2_14[4], stage2_14[5], stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9]},
      {stage3_16[1],stage3_15[7],stage3_14[10],stage3_13[11],stage3_12[17]}
   );
   gpc606_5 gpc588 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[10], stage2_14[11], stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15]},
      {stage3_16[2],stage3_15[8],stage3_14[11],stage3_13[12],stage3_12[18]}
   );
   gpc1_1 gpc589 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc590 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc591 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc592 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc593 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc594 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc595 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc596 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc597 (
      {stage2_0[8]},
      {stage3_0[8]}
   );
   gpc1_1 gpc598 (
      {stage2_0[9]},
      {stage3_0[9]}
   );
   gpc1_1 gpc599 (
      {stage2_0[10]},
      {stage3_0[10]}
   );
   gpc1_1 gpc600 (
      {stage2_0[11]},
      {stage3_0[11]}
   );
   gpc1_1 gpc601 (
      {stage2_0[12]},
      {stage3_0[12]}
   );
   gpc1_1 gpc602 (
      {stage2_0[13]},
      {stage3_0[13]}
   );
   gpc1_1 gpc603 (
      {stage2_0[14]},
      {stage3_0[14]}
   );
   gpc1_1 gpc604 (
      {stage2_0[15]},
      {stage3_0[15]}
   );
   gpc1_1 gpc605 (
      {stage2_0[16]},
      {stage3_0[16]}
   );
   gpc1_1 gpc606 (
      {stage2_0[17]},
      {stage3_0[17]}
   );
   gpc1_1 gpc607 (
      {stage2_0[18]},
      {stage3_0[18]}
   );
   gpc1_1 gpc608 (
      {stage2_1[24]},
      {stage3_1[4]}
   );
   gpc1_1 gpc609 (
      {stage2_2[21]},
      {stage3_2[8]}
   );
   gpc1_1 gpc610 (
      {stage2_2[22]},
      {stage3_2[9]}
   );
   gpc1_1 gpc611 (
      {stage2_2[23]},
      {stage3_2[10]}
   );
   gpc1_1 gpc612 (
      {stage2_2[24]},
      {stage3_2[11]}
   );
   gpc1_1 gpc613 (
      {stage2_2[25]},
      {stage3_2[12]}
   );
   gpc1_1 gpc614 (
      {stage2_4[45]},
      {stage3_4[14]}
   );
   gpc1_1 gpc615 (
      {stage2_4[46]},
      {stage3_4[15]}
   );
   gpc1_1 gpc616 (
      {stage2_4[47]},
      {stage3_4[16]}
   );
   gpc1_1 gpc617 (
      {stage2_4[48]},
      {stage3_4[17]}
   );
   gpc1_1 gpc618 (
      {stage2_4[49]},
      {stage3_4[18]}
   );
   gpc1_1 gpc619 (
      {stage2_6[51]},
      {stage3_6[20]}
   );
   gpc1_1 gpc620 (
      {stage2_6[52]},
      {stage3_6[21]}
   );
   gpc1_1 gpc621 (
      {stage2_6[53]},
      {stage3_6[22]}
   );
   gpc1_1 gpc622 (
      {stage2_7[47]},
      {stage3_7[20]}
   );
   gpc1_1 gpc623 (
      {stage2_8[70]},
      {stage3_8[23]}
   );
   gpc1_1 gpc624 (
      {stage2_9[36]},
      {stage3_9[21]}
   );
   gpc1_1 gpc625 (
      {stage2_9[37]},
      {stage3_9[22]}
   );
   gpc1_1 gpc626 (
      {stage2_9[38]},
      {stage3_9[23]}
   );
   gpc1_1 gpc627 (
      {stage2_9[39]},
      {stage3_9[24]}
   );
   gpc1_1 gpc628 (
      {stage2_9[40]},
      {stage3_9[25]}
   );
   gpc1_1 gpc629 (
      {stage2_9[41]},
      {stage3_9[26]}
   );
   gpc1_1 gpc630 (
      {stage2_9[42]},
      {stage3_9[27]}
   );
   gpc1_1 gpc631 (
      {stage2_11[45]},
      {stage3_11[20]}
   );
   gpc1_1 gpc632 (
      {stage2_11[46]},
      {stage3_11[21]}
   );
   gpc1_1 gpc633 (
      {stage2_15[1]},
      {stage3_15[9]}
   );
   gpc1_1 gpc634 (
      {stage2_15[2]},
      {stage3_15[10]}
   );
   gpc1_1 gpc635 (
      {stage2_15[3]},
      {stage3_15[11]}
   );
   gpc1_1 gpc636 (
      {stage2_15[4]},
      {stage3_15[12]}
   );
   gpc606_5 gpc637 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc615_5 gpc638 (
      {stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9], stage3_2[10]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc2135_5 gpc639 (
      {stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage3_4[6], stage3_4[7], stage3_4[8]},
      {stage3_5[0]},
      {stage3_6[0], stage3_6[1]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[2],stage4_3[2]}
   );
   gpc2135_5 gpc640 (
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10]},
      {stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_5[1]},
      {stage3_6[2], stage3_6[3]},
      {stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[3],stage4_3[3]}
   );
   gpc615_5 gpc641 (
      {stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15], stage3_4[16]},
      {stage3_5[2]},
      {stage3_6[4], stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage4_8[0],stage4_7[2],stage4_6[3],stage4_5[3],stage4_4[4]}
   );
   gpc615_5 gpc642 (
      {stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6], stage3_5[7]},
      {stage3_6[10]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[4],stage4_5[4]}
   );
   gpc615_5 gpc643 (
      {stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11], stage3_5[12]},
      {stage3_6[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[4],stage4_6[5],stage4_5[5]}
   );
   gpc615_5 gpc644 (
      {stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_6[12]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[3],stage4_7[5],stage4_6[6],stage4_5[6]}
   );
   gpc2135_5 gpc645 (
      {stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage3_7[18], stage3_7[19], stage3_7[20]},
      {stage3_8[0]},
      {stage3_9[0], stage3_9[1]},
      {stage4_10[0],stage4_9[3],stage4_8[4],stage4_7[6],stage4_6[7]}
   );
   gpc135_4 gpc646 (
      {stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[1],stage4_9[4],stage4_8[5]}
   );
   gpc135_4 gpc647 (
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10]},
      {stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_10[1]},
      {stage4_11[1],stage4_10[2],stage4_9[5],stage4_8[6]}
   );
   gpc615_5 gpc648 (
      {stage3_8[11], stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15]},
      {stage3_9[8]},
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage4_12[0],stage4_11[2],stage4_10[3],stage4_9[6],stage4_8[7]}
   );
   gpc615_5 gpc649 (
      {stage3_8[16], stage3_8[17], stage3_8[18], stage3_8[19], stage3_8[20]},
      {stage3_9[9]},
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11], stage3_10[12], stage3_10[13]},
      {stage4_12[1],stage4_11[3],stage4_10[4],stage4_9[7],stage4_8[8]}
   );
   gpc606_5 gpc650 (
      {stage3_9[10], stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[4],stage4_10[5],stage4_9[8]}
   );
   gpc606_5 gpc651 (
      {stage3_9[16], stage3_9[17], stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[3],stage4_11[5],stage4_10[6],stage4_9[9]}
   );
   gpc606_5 gpc652 (
      {stage3_9[22], stage3_9[23], stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[4],stage4_11[6],stage4_10[7],stage4_9[10]}
   );
   gpc606_5 gpc653 (
      {stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18], stage3_10[19]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[3],stage4_12[5],stage4_11[7],stage4_10[8]}
   );
   gpc606_5 gpc654 (
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[4],stage4_12[6]}
   );
   gpc606_5 gpc655 (
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[1],stage4_14[2],stage4_13[5],stage4_12[7]}
   );
   gpc1406_5 gpc656 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[2],stage4_15[2],stage4_14[3],stage4_13[6]}
   );
   gpc2116_5 gpc657 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {1'b0},
      {stage3_15[4]},
      {stage3_16[1], stage3_16[2]},
      {stage4_17[1],stage4_16[3],stage4_15[3],stage4_14[4],stage4_13[7]}
   );
   gpc1_1 gpc658 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc659 (
      {stage3_0[7]},
      {stage4_0[2]}
   );
   gpc1_1 gpc660 (
      {stage3_0[8]},
      {stage4_0[3]}
   );
   gpc1_1 gpc661 (
      {stage3_0[9]},
      {stage4_0[4]}
   );
   gpc1_1 gpc662 (
      {stage3_0[10]},
      {stage4_0[5]}
   );
   gpc1_1 gpc663 (
      {stage3_0[11]},
      {stage4_0[6]}
   );
   gpc1_1 gpc664 (
      {stage3_0[12]},
      {stage4_0[7]}
   );
   gpc1_1 gpc665 (
      {stage3_0[13]},
      {stage4_0[8]}
   );
   gpc1_1 gpc666 (
      {stage3_0[14]},
      {stage4_0[9]}
   );
   gpc1_1 gpc667 (
      {stage3_0[15]},
      {stage4_0[10]}
   );
   gpc1_1 gpc668 (
      {stage3_0[16]},
      {stage4_0[11]}
   );
   gpc1_1 gpc669 (
      {stage3_0[17]},
      {stage4_0[12]}
   );
   gpc1_1 gpc670 (
      {stage3_0[18]},
      {stage4_0[13]}
   );
   gpc1_1 gpc671 (
      {stage3_1[0]},
      {stage4_1[1]}
   );
   gpc1_1 gpc672 (
      {stage3_1[1]},
      {stage4_1[2]}
   );
   gpc1_1 gpc673 (
      {stage3_1[2]},
      {stage4_1[3]}
   );
   gpc1_1 gpc674 (
      {stage3_1[3]},
      {stage4_1[4]}
   );
   gpc1_1 gpc675 (
      {stage3_1[4]},
      {stage4_1[5]}
   );
   gpc1_1 gpc676 (
      {stage3_2[11]},
      {stage4_2[2]}
   );
   gpc1_1 gpc677 (
      {stage3_2[12]},
      {stage4_2[3]}
   );
   gpc1_1 gpc678 (
      {stage3_4[17]},
      {stage4_4[5]}
   );
   gpc1_1 gpc679 (
      {stage3_4[18]},
      {stage4_4[6]}
   );
   gpc1_1 gpc680 (
      {stage3_6[18]},
      {stage4_6[8]}
   );
   gpc1_1 gpc681 (
      {stage3_6[19]},
      {stage4_6[9]}
   );
   gpc1_1 gpc682 (
      {stage3_6[20]},
      {stage4_6[10]}
   );
   gpc1_1 gpc683 (
      {stage3_6[21]},
      {stage4_6[11]}
   );
   gpc1_1 gpc684 (
      {stage3_6[22]},
      {stage4_6[12]}
   );
   gpc1_1 gpc685 (
      {stage3_8[21]},
      {stage4_8[9]}
   );
   gpc1_1 gpc686 (
      {stage3_8[22]},
      {stage4_8[10]}
   );
   gpc1_1 gpc687 (
      {stage3_8[23]},
      {stage4_8[11]}
   );
   gpc1_1 gpc688 (
      {stage3_11[18]},
      {stage4_11[8]}
   );
   gpc1_1 gpc689 (
      {stage3_11[19]},
      {stage4_11[9]}
   );
   gpc1_1 gpc690 (
      {stage3_11[20]},
      {stage4_11[10]}
   );
   gpc1_1 gpc691 (
      {stage3_11[21]},
      {stage4_11[11]}
   );
   gpc1_1 gpc692 (
      {stage3_12[18]},
      {stage4_12[8]}
   );
   gpc1_1 gpc693 (
      {stage3_13[12]},
      {stage4_13[8]}
   );
   gpc1_1 gpc694 (
      {stage3_15[5]},
      {stage4_15[4]}
   );
   gpc1_1 gpc695 (
      {stage3_15[6]},
      {stage4_15[5]}
   );
   gpc1_1 gpc696 (
      {stage3_15[7]},
      {stage4_15[6]}
   );
   gpc1_1 gpc697 (
      {stage3_15[8]},
      {stage4_15[7]}
   );
   gpc1_1 gpc698 (
      {stage3_15[9]},
      {stage4_15[8]}
   );
   gpc1_1 gpc699 (
      {stage3_15[10]},
      {stage4_15[9]}
   );
   gpc1_1 gpc700 (
      {stage3_15[11]},
      {stage4_15[10]}
   );
   gpc1_1 gpc701 (
      {stage3_15[12]},
      {stage4_15[11]}
   );
   gpc2135_5 gpc702 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc2135_5 gpc703 (
      {stage4_0[5], stage4_0[6], stage4_0[7], stage4_0[8], stage4_0[9]},
      {stage4_1[3], stage4_1[4], stage4_1[5]},
      {stage4_2[1]},
      {stage4_3[2], stage4_3[3]},
      {stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1],stage5_0[1]}
   );
   gpc615_5 gpc704 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4]},
      {stage4_5[0]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[2]}
   );
   gpc606_5 gpc705 (
      {stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[1],stage5_5[1]}
   );
   gpc615_5 gpc706 (
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10]},
      {stage4_7[6]},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[1],stage5_8[2],stage5_7[2],stage5_6[2]}
   );
   gpc7_3 gpc707 (
      {stage4_8[6], stage4_8[7], stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], 1'b0},
      {stage5_10[1],stage5_9[2],stage5_8[3]}
   );
   gpc1343_5 gpc708 (
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[3]}
   );
   gpc1343_5 gpc709 (
      {stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage4_12[1]},
      {stage5_13[1],stage5_12[1],stage5_11[1],stage5_10[3],stage5_9[4]}
   );
   gpc615_5 gpc710 (
      {stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10]},
      {stage4_10[8]},
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage5_13[2],stage5_12[2],stage5_11[2],stage5_10[4],stage5_9[5]}
   );
   gpc7_3 gpc711 (
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7], stage4_12[8]},
      {stage5_14[0],stage5_13[3],stage5_12[3]}
   );
   gpc615_5 gpc712 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4]},
      {stage4_14[0]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[1],stage5_13[4]}
   );
   gpc615_5 gpc713 (
      {stage4_13[5], stage4_13[6], stage4_13[7], stage4_13[8], 1'b0},
      {stage4_14[1]},
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage5_17[1],stage5_16[1],stage5_15[1],stage5_14[2],stage5_13[5]}
   );
   gpc1_1 gpc714 (
      {stage4_0[10]},
      {stage5_0[2]}
   );
   gpc1_1 gpc715 (
      {stage4_0[11]},
      {stage5_0[3]}
   );
   gpc1_1 gpc716 (
      {stage4_0[12]},
      {stage5_0[4]}
   );
   gpc1_1 gpc717 (
      {stage4_0[13]},
      {stage5_0[5]}
   );
   gpc1_1 gpc718 (
      {stage4_2[2]},
      {stage5_2[2]}
   );
   gpc1_1 gpc719 (
      {stage4_2[3]},
      {stage5_2[3]}
   );
   gpc1_1 gpc720 (
      {stage4_4[5]},
      {stage5_4[3]}
   );
   gpc1_1 gpc721 (
      {stage4_4[6]},
      {stage5_4[4]}
   );
   gpc1_1 gpc722 (
      {stage4_6[11]},
      {stage5_6[3]}
   );
   gpc1_1 gpc723 (
      {stage4_6[12]},
      {stage5_6[4]}
   );
   gpc1_1 gpc724 (
      {stage4_14[2]},
      {stage5_14[3]}
   );
   gpc1_1 gpc725 (
      {stage4_14[3]},
      {stage5_14[4]}
   );
   gpc1_1 gpc726 (
      {stage4_14[4]},
      {stage5_14[5]}
   );
   gpc1_1 gpc727 (
      {stage4_16[0]},
      {stage5_16[2]}
   );
   gpc1_1 gpc728 (
      {stage4_16[1]},
      {stage5_16[3]}
   );
   gpc1_1 gpc729 (
      {stage4_16[2]},
      {stage5_16[4]}
   );
   gpc1_1 gpc730 (
      {stage4_16[3]},
      {stage5_16[5]}
   );
   gpc1_1 gpc731 (
      {stage4_17[0]},
      {stage5_17[2]}
   );
   gpc1_1 gpc732 (
      {stage4_17[1]},
      {stage5_17[3]}
   );
   gpc1325_5 gpc733 (
      {stage5_0[0], stage5_0[1], stage5_0[2], stage5_0[3], stage5_0[4]},
      {stage5_1[0], stage5_1[1]},
      {stage5_2[0], stage5_2[1], stage5_2[2]},
      {stage5_3[0]},
      {stage6_4[0],stage6_3[0],stage6_2[0],stage6_1[0],stage6_0[0]}
   );
   gpc615_5 gpc734 (
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4]},
      {stage5_5[0]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], 1'b0},
      {stage6_8[0],stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[1]}
   );
   gpc1343_5 gpc735 (
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0], stage5_9[1], stage5_9[2]},
      {stage5_10[0]},
      {stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[1],stage6_7[1]}
   );
   gpc1343_5 gpc736 (
      {stage5_9[3], stage5_9[4], stage5_9[5]},
      {stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4]},
      {stage5_11[0], stage5_11[1], stage5_11[2]},
      {stage5_12[0]},
      {stage6_13[0],stage6_12[0],stage6_11[1],stage6_10[1],stage6_9[1]}
   );
   gpc1163_5 gpc737 (
      {stage5_12[1], stage5_12[2], stage5_12[3]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[0]},
      {stage5_15[0]},
      {stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[1],stage6_12[1]}
   );
   gpc615_5 gpc738 (
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[1]},
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage6_18[0],stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[1]}
   );
   gpc117_4 gpc739 (
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], 1'b0, 1'b0, 1'b0},
      {1'b0},
      {1'b0},
      {stage6_19[0],stage6_18[1],stage6_17[1]}
   );
   gpc1_1 gpc740 (
      {stage5_0[5]},
      {stage6_0[1]}
   );
   gpc1_1 gpc741 (
      {stage5_2[3]},
      {stage6_2[1]}
   );
   gpc1_1 gpc742 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc743 (
      {stage5_5[1]},
      {stage6_5[1]}
   );
endmodule

module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor_CLA256_12 compressor_CLA256_12(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h1b395358a517dc210d3587c4a6076e79e310f217b7f6691db9211f42133dcfbaf3f71bc3c2e9662b6896576e2559f5b8b1f815f76de39f04f75b4748083a5013f19204f35a0e51b86e4f1434a772203990a340e91815c3983aa6730c6107ed548e2aa0d7220a3c7d58eb8c28579fa7df569f5b6a5f9a560457c3c1106c98ff5e76c3ea05ffeae269f7b8674cd51a41649544bd4c0bea7f9c9397d579b591882ce3abdbd379b2054ecbd310db315712fb1b6bbf2614a2d9eee1b6684f2a37d8952f962442bdabb6449a25fb1f09709dfeeea1770f661e240e47272759ea178fef4d147f00d7860e83e6d9173c97d080b425ba2aa5ec0741698afcf32302231910e617fbddf31de0c92f7980fa3b3015f39a4e03272be93527a1fde7d44dc910e95ef125614ee9cde33c50dc2e484308def5ef3bbe7f619ca92af9f6a80321193fa319969c954b04b6847f3f89b055485934f2dc4e3843a0d359b3b3201e8c9b0d8e6813b11d3472230aad42dbc0d5f1cd693a1d05fac2e59e4e782abd4e0696c3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h898a81e5573acb6d95ac044582b08e652a5b07111c792acff54e15c73ea2aefe73373395e45efca8411e215ab0c20de93654613c12ca9ff117f53ab65c1815f94075ecdcaf5b097a68315dba3aa7fd217edeba83da1e852f0b240556bb59bc789f4947ce105b3c1a63ce8432c781faf2a8f8239d2e0d92b63a41642ab04629622f51b7c95f963d4aa9b608e04c94882936d7ffa9e8a80c17d0a997d0484e524dd605438426143b175de6d92ffd60213482687915e57de1cbba59e4415848dde981cae0290cec052c65839d673fbaaf449c5cff937c728fb2e43df5f84e8920fd18a9d85e4b9f29b8a19f93d5e9044d36614271cc1c17fc1cab9c6bb7d083423c606d66a02e5bbb166648a55eb3a144bb4d898094db6ff48992d24c0e2d011a7d2d5a0b56da3f5723987ba5ed226644ef8260c86b5fa4f79fc65c54b7981b808a3df455d0881f4ebc86e1d85bb593187d7e4f1e0fc256987634ef63d9a99be299a644c1b935aede1268c76393ad019e0331242d48c7e478d8a7f8831ed1ef0cde;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hb1f7bba0111a0b711f30b29a4270a465ef2356ae6367854dae1068664ea0fd0447092cb96409a455d6c03d6a68a387ac62fb44074291b59d533fdd8d6efa9ca34dbdcf7df1b3a3c9ec3c4e21bfc9f796622c9ea2ae7cbc4cb5a236e678b88fb17165acbfd1288a685923b6d75749bbfb1768cc0b00ce1889fb334426b9120b6a445f388070339850cb9fa5ca60bed0408baed493360217619b2d3ff651887b98bb3cdd824f1f6e7be6203af1d60908fc665b5511e97c505b4dd201b0ac2a587e184ec3f3e2cf0d1b343901b8c6a3b65e30eeb665b41efc4289018d8cd760e41adeb0ae16be1499aafd4ef8dfd82a0297346b6c4a7c422570cfdf556fb46f105828f0f7b1a91015fd880261983c232d7c72d80f0130ba7fd0b490a715b0cdd6fe245b92bd0fdcf91234d8837d5b896454f3b43f2329c0ca41c69dbea5d00e4a1a35b57ab447480fb81c0483841c92441f2f1d3192fef16fbf4e1b3eca00b311ed4bb29a00519de0f279a789a3054b38194ce699adb1baeb09248878227d67184f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hcc8ee3a4b1dc614c32f622ad3768d6fdddbbd1b697ce787570b5d2ee4056af41228a56a5286632f90f93365760ebda2597d86336934c647d0d017f968bec5584b0e73661b84f7e667eea50b1f67e2a9963d79c6df7bcc42ba1640202fd0f4bd520382a81e48d0893210c6305c36589c7ce90748f8944854f17440d840a87bf3a251ab04287a0a5a70f5837190dacd8482402e2ff2249518e3b0368817fe76066fbd6672b8c99721fe461dbdff78628b52ecc624399624c2bb3ab6532276e1550bc209197a251a84d02291a8728e33638ff0e2a1bd5a17e0d45e270f91f6e7880a69b0a9818e1cb04ad3743fd1cfc648cb2befa0103292467dd87cb2c6d85e96d960f7675cbb6358839fbc7a62ebfabbd71102132892ca6e10efefa730d1ea14311b218fb4d7e2db6f21e71f5fb92990f3225ba058dc0a53361c17d0425cf171c56d20cd1bbff77176d69e712314d67b0bb9f5d9249ab4b6b0fe221e36a46f933da9dea3740022f00c3e7a0a2dd4c55f16c3cae577ba5d560cde787425f0ada0e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf749511dab5c6cb32f1fc6d2154583a93c674a063b7098362d954dc776df10849bba511ce8c6ee7c0b14ba0d4e76e266e682320471757b77dde012d553d48d19244161a6ea3091d891b38b5e4b9783ba260cdb2aad303e65eabafbfb4bd38257035c35aba09ffab8d26ad7c0d2b083309df52330729f2d7e668fdb38ecb5bd92f49736df259588cd7753867de1766d92f78bd4f3be5f7982641d9c0cda7b0e1ffc106e390434e84e325880f8e9bf692dee29f17891cb1bbec14202c98aca47c3e713a0991f7ffa8f7b220a03708acade76c4dd29279393c64c1a65b6ed524b36116c215920dd3bde0bd6a2532904b5ac7fec709209bcac242cda1eff01043d7a4e5e8f1cdccd424552b9f79dfc089945dff5061f76a48a4af5cd3317a3a71f4298b8d797015d27148504e78890b1e41a2e1af51f2c8e09949c404c895943dbce1d8a3ad7b153b44e17a7b94ed8aa3b52fc47da5717ce1f1846cbd84cd9c8c9d18e06f0b41d0b9369a59d8c29231c947f326a794c62e06731a4e21b5502f2a736;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h74e9376508c17e1b37b307ae73c97cdb97c2a8e333e49a34052fb1c45e65042c44ed309f2f2e692c87f2b80e60fbe0686641e3354e8dcdd345861e73d4199538eac825069f32853842394cab873cd207d7ddcd1201900489d57f2937970dd8303e23072ceab9032136904c231e1a58f345edd25c3b2012a385cb2321a7753ee91f6f6f02f444b30a6bc4213f2f4cdca319d6142f1e24b37b397f3a6bf8f44afb65a6d032f5cad2eda3c36b15c7184fb39b8dd3f39fb70e4f43083add80823ce433ec223f0e4f6deddb59a9299ec4de24ec5f92f04a1af0d9fa289b55a52a3db3481137c8184d1f26c9b3d0b9dce4e2991b87e72ec01bf0c4a5b4ed548276cdb7ac04ed638bb19581c27bb6097232564ed9abeea61dc6b2dff28ac84db5378ea6d4a2850fb67aad28e17916ffedafb5f92d8587723e4caba0faf60464d519a2ee4cc1692fece1f64bc78f20c89c57445356c1dd39848d793d9ebd41609cf02dd3153009c4ee32c3e22976711db89b4ef7a7d9479a0e9a47afb2d35cd5d8e26b45;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hbc2c3bc41bdb518648c470130ac3986d757f9e1f312412e073c9aa4201230e641fa650f101d60385a1bf5b05f1e1208053ed7cafeed437b596563d86c6f152c7d07540481aff1cfe87cfbf3d31800f5be7323136a854b529d8a37920aa7e729951715641a08b7d458e3f17be23cd21c115e540e12306fd83bf752e6a6b31733400ca7dc8aef65c700a931c35590572eaf83860c61fb4f6e38f80dc105050b9af6635273b3185e1175127149894464edef3a9b58cc422d840f49d0be4ed9aebcd9884b1b18f8e728c8ba269d70b6435ba579b6aa540967f396d09d9d7077eedcc160945bc9791f243c62f31e4bfee22bb000b829abfc978c956ad6dd70735c1d0abcd0def9a584cc0ce533b38c32503ecae333015bd7cc0335c1445809157b50c331e4a9d944ce1d7d550d441821738b65b82db8a1bfe386063caf03cf19ecbfeef8971168a24e6abc8df922db25cad262e73760f2a97cfe5ca09ddf9e5797ba8508a21c3d6bc9e250bf48a5738225f08495c3d2b60651da8cd862f1d096f9b0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h73057251c57031647d60c15f05c0c4a16138e24498bc171d35830880aa3e285d3ab4758301dcc4c82b7f811d49e3e141d99c5002f9f7d425c3734232100a92670bf56a75687994abb2bd9ec00780874c8b4dbca6fb06ca3d8843ce6991583747da49da82286b102154d210e5150160fc5ad3384dd091c6a395d1e542d1507f6dcb88abf75ab8290423b6889b77f036985478846dfab44313ebe1504ab5c5e09458ee892cfd3cfc170f5848f376528bc34e80a131e199cc7c5f2f75481b0468b9dbef9e481820a8cece3def2b2dd0dc2d4f605a460a76403db51911dc95633ab338281bfffe50928dc770126183e778d0cd34515236b379e97696477a1aa92893333c4ee1db2d02c2832e5eab003e3eb3601228fc107cd19e8d5ebd25ca522524ed20dd01ce336048fb5c9087424106da9f86ec6c868260a2da4683c1b00abf15723eb8fc25310b8716d95f14e35ca58257fc1123a96ffdca804b39c6045bef534e3d4971d0de9e28b7914c633a60e6bd486913ac314ecd7ed4ad8df29df563e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hbb29a2556bbe8793ee12cff0b930e53b5267c825fa407b50a52a410e67d2451952f26801d4941d807a5a1dda02c74600e8394112a6f81f46ce6229b6fb2eb686d7d318630c41c8a67a0cc8672a1d19f622a80c79d3914fa8eadf9742112e2425fd09514daa91975e2f225a7820cce3c4ae86920a364dd411d2bd399d5a0846d5500a79d318869a45c7bc0b95a6539a2979fda6498153e81f5f2e111a781ba98a40c3a25674b3cab96a8dcb4476aec938ae8fef29551276a5f0e32c7a616f42af8dfbe127856de5cb4ca341e73161da33516460430bf2a2b8c7d54f90ffe45eb1f118e96d50123b98e3bceb803a761778cdf36fa9dcdd2ea92f14c223a54734064b44dd5e6fa34fa699a1ae530534f02f869bfef2aed55f8844db01b681a95ef7800fcc5e41bfe12a393b7f74ef7fa15ab6411d59a538586ce41eb822639a5c53f672665e744aed27b03e5c898bc58fcd50ec86a8aaddb80272a8e8794cb5b9e910a6fcc36a360d7520b131819680ca62dd1f9a6861039a9a4c61192ae4b7fdbd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hbd599f3fce2c06bd018a8f76957a741f85ca7e1aea563c175c2911b8086eb95678a41654fcd1bb3cf4a6a8890959644064a19373a57312614c2600b48d79462f9338e47e9f67e3d3bcdde57b527b2d7e34f343e7001778eeea52937a71baf9fcde12ebbab91e15b87f831e4536caaa7466518a7dfc78a671394cfb24cd6f06d4711e2a837be34c851d82e6d6381381bb03f749741cb1e9f60f048257de9ad3923938320532490a13f2710fdaedff0146a998977db45a79466e507711d4ffb6c053f5a6970a53f02bb12043039cb430570e009e7894a20c99a3637bedbbd56688c2c49fa1a78fb7c1fba744bb662763e37c744468c9fd9bca3240704ecc719ddb74666854bdd89ab97caa0e6e8ab20070385426bb3baf6d5a1bb8f8eac2b3b1de7c36d423b50fbcd5c84db60d5bce8cef95ccbb5db911038aff57b3cf2a61f5a55f719719ffe1fc000135b7aa1c9f46aca137a4cd82536d2d70ee04274b06217ca708e7e1b95a2528c324d857a0c12136c0364142d0945e17ed187427751b46f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha2fc4185de815a8114aec38311d0f120003e8038b54442d59875a97bdea079e8a4f9b35b3700c2d301808ae884002e76f38174cc1ebd4f724390caca0f8ffc4ead0bb6c4fd82536a7cbfd71359d89d440be136078fd85b394affe4d2df1b205ab7207851300419d08b8e096477d5ccce7b2a058945860881f3b31bced29b9ef954e30726bc52b804fed43ebcd201ec9017e4fc5cc8b08625cf7639caf57d71505e2f8e55f7351c5642fe70b402db75abf752df9b6ef86dc21e6b2b11bcae627df0c42a01a36c0294f2eb06a4750ceb3482630003c625fa090fa70909d1ca4c39aa0c0a52b352f72f3f0e512ea5b1e8ddeebf75d7cedf12cda56e8c9d2ad9034107a2dc8b2fa066cead8840ee687b39d74a6c30edf8efb7fc65a00c8784cf1ebe20da8a490f45d55df00583a546c9b147ad772743cffac3fee5b84b40c6932fee30d7573d49b8835c215a79bd774a133621200febda93ab6344203d2f6446950d18020c8c64ad4cf7e9a03cf4f1c1ab85002b83891d72e2020517e1c5f1088418;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'had327f22dd39e36894b84163a89b087bfa8f6d99d4da0afdd83bf8898caaa5ad643333fbf5c88c518784f622f5d8492827443e5ddc670d7198a9d8aa64cb98378a1a8a5885cff9e587d4bb870ee91512f094db36237167368655f91032389a46d3e6917b4c7d673eaa6b3a8c8b278ffb225fdec745ec09dfbae8b3490e8c60dc72b3a9b483fc08c0643cb128ff8419133308b43200f06f9ba20d9329004405dcb538f0876b3ee7cdea54cc6a764f83926869e661e0cd68ee1d5a121971d339a6c7e2d859e51ac4e4ee238e8b7f1f30c30930f035c345cd02ecf443ad8a55bec41c5b73cadc776afefff817fb4bb26d0f62575b96d3db3d759ab3bd6fb66ff132e4e0693665cba225919bbb8be2dd785fb102dfd74f292aa1b3627a6dd64677d04c14f2dfabf81eb377aa52371f3083f686478ce82e7c5432f1d033146baef3b8957037e676b70660a1d661ca2b4b62e1c988173de9f424b4b725b3121ada74570f2b47863f72f1acaa9aa2437a0859403ba1255a4d5163960a17163db72f29db;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h79412a524e1e2732e5f3bd41e9cbbc563cfec2438fb24ab34b0e929ec3aa0399a43f487b690eb5ebbe6bf91fff7ec5190df37823027505056e50e6db2a01d4e82028729c211de28feb53ca804c0d9ca362f2856870fa1b6e158c812e6cd60bf17b126c6bf70d504deb3549bd967e176122226a26876ccb2e7ef26c7eaa404d79362c0a8ca9df43020b6e3b40f0d016d656508d98aed910dc0396100d6677455b45d837b0d6a7147283e772ec47aacecb089223061c72a7270336527a81c1613e6d7624d95942ae9f3976f90a7c52a9abbe3fd588cea0b589bbc8d02973128d719e322603a9d3c9cacee700afa0e28b6dd9777b258d2a835f5c2e6cb1cb5a2165137dabf62f956e41ec4118f4254aa6b4ac4c2cec28281b9dae65c9515a3f6c29a39f6c114c099d242ea105aedb224bcd74bd23cdc67643aee11cb7d6f6b829c655cde275e9f62077361129abe17a3c976fa882cae677a931217a19a0fb59ae8899dcb1a56277125d1bf41bd3e9c1076725597727ba79decf00cbd13f61476ffc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h81eec59b61b024a2cc6d485a387a70292cfc67f3b1e5965a8cb561200bc0515aa3e8644c0756934f9685a70c2231cb173579488bbfc0f84b0b44e4cbcd17ae92643e4137cbb297e20dd57f00908c016a447f64fae32a6728a8033265948c8673c94fa22f49606b02f22dfe65e4bcb7643d7cb49f26ce56832e8967302245abeb07badc96a249791381d8e77d2d2fe02ccff79c6283c2698c690466f039d94373fc0c30fe38c381b06e32d44ebab8966b4e6688377f8847789cf785b98b2a665afcfea977d9c03e125ec271ba73ba756310a8c93d74f6abf049e70d9da13819e8025bf8c9e28bd91801544cd3365ebcd98c3cf087782065c40ea0eec6cdaa30213265c3168bd0c722de52c688907b22ab0c56164f9c0fc74371ecd66a17158e8c69822572a137e79a05d2410177bd13ba01611cf02bf75bf58c4601442fcf6c5b0c3d8a1690a0e757dd42c6de3cbb1886ab72587e1f94711e08cb06ea045002410ddcbaa1fff0bfd077ad7dfec4fd1e63fc483544080b6a5210e5b3c06c998106;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h95b39fa59c3853f3782dcf65813a9865d70614da9e78204823cca39fa0671b74658480b00d4ca3991523be46e74d32486e74e92e483c7d8a6ca9709b617e0179cb09cc91c4b2b72d4d0ec8b6444b1d443ef97d7285e376f46995cdd709e506e8590e8adb098d0d1a9f180efcb868c199fde6a0c0bf3331f1eb0128eb8cbc3d840b3dcc7f77af4b10da877e8900546afa780a98d4f20ea92256249ea9604602de9f58e1ee64c6305b93416715ba6f801590276a25300520b0ca8da17214313f3348a7b26eeb1b43339548b4d24fd4980e6b54e4cf25e37eb59a4ba3cf05ed4b6a45d8e94727e7b73c34bdbc6e2a0afa37f176ec9fccfb074c1ec003a3be349e134a99079f66f82e42b129cd333c130652adba9e4d734411e9c022018b156155f40369ceedf18270042d1ce195a0fcdbe071f935d711ea2c450d863c5888aec7c41a8c12b9c433856caee05aa6d58b3e9f72bdfc1aaa835900829d7ffb816cd070ba3905e76717ae8a60470ba590df2b8851c3434c969b605e31018a0069222f2f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h71282c2260e0cad89c88dcbd800a4dfc614810c7f9f07b22af6ad016a898f81ad729fb2abc24fcb55fe3d638c6267ae89f2da8d6210c75eb2bca3f87c2af7e3be1fb08388d8eef7fc2e9b3e4eda8092e3920e6ff21a7c0c4c4abd07e1e24094164b5efd53c49d263531faa5a81eaf5fb4b8f4b2ebe5ec4b8bcd542ec724a2b99642359909efb0425e4109e3533cc39d15c1cefaa4e72b9879d7aecc7e49e75fafda8b5f43a4190b51ac83608477e51e51e0b8173eab373401226ccd1387486a4ceeafa1330b42a569394ab557a6afb6cf77abca58c91ac4c5c4c49226cb6604e3e52c7cb33da188f8248e06fefca6a68c873e661923f56b4524e4815a1aa91e7188fbe31212404d6a4ff695fbf5cab06916f32510e543c8209eb9f370b14f0ad763a30d7e9e1b4600f01d0d4627578520cc084e56685d4261a7d0d87738c2f19a415437c268c3efd34b2299bc36e5ac2647b469afd7090a59c392d525b102ca25db2199ce956af990c48bc2f709568deb5eef6c35dc5365280d5f9f2f0d919a3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc34cd765606e3360e7bb0b1cb69d8d1bd9bfe0a91b14e9c7f3b8545ddb3717d81023d78ae3960634480dd1efddf76d4f714ceba65d9cb492f778b0fd741a95a81d98bd42b7b5ab1f58a6d735b65756527c2e3060dfb53881d760deebf4419fd231a6168b52513c9be22b922a4ea74ca2744e2223917cb9bd06562ccbf832ccacfcd42870887331b6a946f1423943bfab62a3326637f446713b40ee8ccb3270df4ed8902b61cfa5f9e7ff9e5d66a94fa6d5271998233d76a8afda10ea43af45fba59a7e118c0b40a2344e490849461be466687a0bbdfdace5299d17de7e27fc1433660cac9a5fc9504d4c094851416074576541118e06337fb0af53edafb2bed5193681064f0461ecaf86a14f81522f540612b2ebb0753a49f38f35209a646ac8b356cec8be4156d51efae154a7d20ab7732277ad3eb3e63fceaaff35f5a9b0860caf48f84575105e77eaa5f372960078a0bf14bf231af205a0dadc0a33c840810c3178e8cf24786dbe867f49c5b9d10e0b49769f6748d830c8d7db8759a671bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5f341b6daf7226817f8249e30000dd76e5994de2c480bb0a9aac9b34bae7b64b9e94e1197a12ba5352bcfa91d329de9d84e74df8706878517cc0c20c5f831c733254b7e66db7b36c22b3e51bb3209ec3752a1675ec8ff2d74fece64c87c748f480f435366019a0722e0b8df0082abb43e6f4f4ab0e17eb7d829ef4bbfe22ab993eb5d18ef4d6eb5e6739620359d7acf76419717e9be908a9eb0cbc16c0a66c90c7a485d574f1484affa53d43feb4448d71a94e50bda347db876ed87612b4811a5663caf78773eb38fa02e918470ecc2f178c4a79a115782f846e08fa71c77828af1188544d3b14c952f7616de89b9920c9b35dac7dbe1ebeead879ac90178fbc50a2c9fa29fde74b6dbbdfba91e9d02eb9e93bc9dafe952dc0b611cf1f3df78e085ad43dafa03d305068edb91432e1bd79547febdf62c891d5aaa630ff75482f518b14b35d630c03006f66fd26621f235d473278340ead94c93a9a7bc2ab809f666d5869b4b6ecef7d46f9c104672c203284186a5b7038c61b318e28a50554e0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h8124b2dee37a25529b8ea4689d93708f7ca4494d8b83b08fbca601d3bcf0adb76955d1021027ccb6a0920f311502fd3d1e34bb18a132790dec14bf5d977f7fbb9653ce6e4d5f1726bb43e52434e2741bde67292c9e5651f24c7b7db042b7445ebc366ad64eb48d93993dbc96014700c457ec1b37a4f0de2fb3f141150f8211e1a2e336a3a765de6d8212cc33cdc482fc556257709a057c72c6902349e46d4e21a3c9ca4adc46591f4450e637f09e71aa82b2e7ff6b948e29635d9756b8bf4729f9723aab0c26ed3c803cd6725cd0b6bac9715d661c567d6f994359cc95cab7d8fe537ec0d82d49043d12f78d242cbad4988235ed72c8d598716a2e836a19b601236fbb4b626f0a415a49efeac8a345c97bb499e4dd653fdd8a23e6d556c2ba4cf63cfcc07d265afce2e9934a15be455a6fb04a599cb927650fcf07140d15ff71adeaf17190df24af77000768bce355a47cc32778c5964414820d88cefd986e78865f23d33eaa86083579d86cbcc159791c6bb91b606c2947fc85e8b4b045d694;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h95e9e1d5020ad8e852305cd580ebbd2a05f786782eaabc22fd510072f426f325fed7ab0f7d84c39abf6e6d2dc6fbca903d69d16b33e255683a2e22fc922ba4db885ffa5e2492572e5cd9faf522edb0ffb712172a5e10b29243034aa5c66d7d0f6147b198186293a8881912b83a6a439b332a6ae273bb4498bfa3e25bbce4fe4584b9f0f82dfc5e8d577716d2a9466ebbf0e346f6761b185761e707b1b530657fcc2d3891645dad7cc310b4f416b14f9202070b76734b5d529b410b1e9a8dc7d00ee538c7f784c0de46ddcd962d25e794d024b92938341b63134e570ebb23b2861c6696d63e58fd9a3aaec9d5d20cfe57dfa4a7b11bcca70dd488c31132a83d17eb67fb98eb8c575be567261496c839c9b760f98c343224ed79598f18b893f3c5ac762648a2643a47e233334168cb63cecebad709c5309fc155d19a5866c24162494dc36c826f73667de67f9a144e80196c5f13b4b58146ca41ab9141ac6490c0c764ef8ad3323b05ae45d4bedb73a322b8bb409ac498db4eb139208b85e2a9ce;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h7a4bd7e9d69ce81188a75036256ea298bffcb8dfaddffab0f24d446fefef89c91f1a16d067494d11ebdd3fb6a6a344bbebd471e46151137fdad562d4ef38adf34aced4f6251bf17b37841dcf77c086847ffcbff17a6e3aa82e1194f77b5cb1880e7bdd88d8b929490b669afd1cfac9657a745edcf587bdcef9cfb80a9c6b56ac1cdb9385dde0ad5bb52e33df02bde425f3168ee76d2728ed62f4fa1d0606c6b915ed816fa052c6d1f1d777e5cd73bc694df866a35393cdc6fb8165a4672d6101ea074cfeffab44245ddfbffb6fa8ddbdf83513d82e2e33f4f1e59e0ec51e1c19b71bd7af4808f758c89fde52d215fe6c2c62cb1f2a310d11194625679f86bc65a3ba6509e5faf5658cff3154c0023a1bd205c02b742fd9b099d66f7519090781f3feab4279c06088061467f6a3dfd8a8716c0c1c08e56b27faf41f4f85574c55d89acfe900ca43f277d4d946fe18b96cec840d7bd2058bf8a12fa449c24a1f24b314381bd6b2abd6bd965f2d997ea1920c66ad8a67a04a7f49d25e114ee5e7df;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hca560c6bc9508a0a4f0bfd2e7649303df5c6be538c8564672773af6798baae86346fb5e999f3a48156b516097390b7d20de1e7b5843e1b140b0b573fcac334b48c787802c9b212c9b303a646e5be2e2b1f55f20dabf2b742b5d942ad869a5645bb4419c2beb68404a72fa49f83cb4594a464c3842d32fc178b0bd45e38619b176d386e5d7fd24b4cb5f95064397a96f8fa2a722ba4440e99ba5c4c80b8480727f18ecefc3febad3af2b88b35c45b6ff96bf00c99769630decef7a4dfae763e5083de3fd8d49a90f822aa6590e8f2b9f97a656d426391d4dfddcd1f88ef6a67e0755de49fe7869c857b37ca041f41b912dc0222541a879645fb70542f40643469ef26bf1a4dcb9fc420acea4f393182a7b657aeb02e6aa2b3be5d8b326abad6bfe654a82eaca56d10c4aac875ca9334a6188bfc07dcf63f039e774a690a5484de5946ac0f7284812c3a8970afb8441dbe9adfb2aa523107557f666fad0cacb3e08c8f4004df69d9a20186f2526716ee293ca3ca5168be8f502aad0570f484edae;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h11de86f63d17de6545d25fd349a305963b5209e75b40ff700ffa9fb98765a9367180e9b7e074888d97e72cdc87750059829c20c5944f4ac7e63a7b92eea58ed3deb3af0194ee8ad32df190d85b2c989563c7a10127f5d74f6b6ab1013cfef231e7d0e2fedf98212f7f99bc05656c5a768c5c14a3fce13782642a72d13bec7f615dbb11ea079c4f17433070249166d3e055f5169b2f7872925e8d50dd44d80d112cd116df6daf377368899fcab63369b96950d223cfbdbbbc454067f4423af676da92c04e439587aa013e4e5eee1df7bac9bef58785aeb61c538225616e1e86a8687c2271695a4c67609745d5f1b90d9480bedbe42d06532b7a8b34a3d9e0a2a5ae04505d7e0b9b0a4f405ebf2a676648dc443a70980beced9f55d7425d962bfff117d883e4c005b50c0c4d147abc3481607d7ec88edc1b5f0f4a1db1246cb9a6b8970314971892b51a0c80601c27400e450f07b455ee978c9a1ba7e9795495bfc07c7988120939f1156e26ddb1b785c4b7d23b3450d1879ff562dbf21c94b07e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'haf613f0ea3cf1848b7d2e8ffd689400100854dd229f9822d63037b33527a028f2207bd323911a3a90ad8b53ae9159f62496e7b4894d350250f986f8df824e7deda18e37f01c78667fc21cd7d6c5876b44187a563df443ed3e45ce0015bbc059829a6abd6d41722fa9fc0a5bce8138c9607ee98c54a8e1c74e04cf37758ea40683c83d8331b9f5fc9fe193a9fc072a6083d38b2e6f941d527acfeeeab55672b7b438f2588dd08270bf0794784a58c3d20fd70cf6cf97c0210d7ddb93eaa0301a1d4ef64868e76c2779976add37a9fb53a283e26df77d1f7bebf1b23864778e53dc5f4e4c73005f89b123a33d44ddb7520af6649fd6fc018b93ff24d0c1942686588716b8c44b302bbe0d69ec778ba128be8b726dd5615f424a6518e2d9b3c53ce4b9eb53d977964d0d728916fd8d72cc1d7bf60a603f9b44b3c0819f463db0675b6aaf2f1d8c8781b93698c4756c8fcdac2a7b3265bc0028d9217d4179593deebfa90bbeceb7a3e49e04c06a1202fc986a50cdce47d4a3e316593c2260004585d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h73a4de17b7b7f14386f51b3cbe0deacccfd2d5bff2f4c926dd57b93d98c8395e63cfd12a9060f9477e29735d7bb5c677ba5c015206ab55de616ac2fd882968343d425c6c8e9176b9b140ae915f643e2bf0f27d2795ffc2fc6fa94995955499df29a28ea7be9d53c84d12eaee541af4876f16356148d178d33dc63452ad1c8a97da80d8e989131a034e9c2656c92be1dfe3e9346e4c9ceac995e5f85abf12de7130615f386d01b1f9419d9e911ed523db36a94e098110145f618e90d9f33f93ca27125296319507bfaec191aad88e4c29835cb87c6cf3137294e6d6dda961ca148c093872fd2c07e6439042acc59d115d4f1b59949fd2e62d003992d91bdb3924919882cb2b35d36e5682412ba737af84fb0bc7dd2be1c7de9fd534ad49e4bf9244f57ce4c5f3bea9c486c89c356d5edc5fa81dedf1be83e9969f253c37cb4e6c2c30f0479489c2e2fc7b039b87313b8c5efcbf6576a1ebfc9e145c7e8a343b00e453663ed0b8579655764ae2d385c10ce94cd3661e00ca57f12bb76bf98f52e2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc8ceb81bc2a77486f61de2bf40f0dacc927e26775cc342805ca46db4551277465add5e0b27f2fc6424ae6bb6dddd746ad445afb8bcae4cff25a85051a23ca4d588303eadd15eeb54d7da77fc9806fa30dc0d37040829c9152dbeb564dec5c705f3e679fbc37284419f3cc2d7f4aaefb4321e1ea8ef81d710a6095b1a4b41e2fe3d2b02de6af21abc5612c4fa6ecff0eefa263df68f8c65ecbc3bde459ab8e69813e9bba7f408ec873a9d149bfdf7465e5f9296b7580ad8d7ae24ec33e5204410a1ce876062e43a20fd326561319980a519fed970daf797035fd4f64c24589148ae1a07e83b9e53e2ab36b21fd68ae82f89c4400adf08b093899b2b06c24623d96ceb1de74a35a653c1a65a653d85a17809db7177677ce3bf6cf622e598adacfacaad18b4017342fbea5887ab90fb7166b2b8076f2d4b17b28f4afb5bad4e661a63ba068fe0a8361e31c6b303c1edfa65b32b348e730b82c29d2693fa31c4b0a93e083d42abcb09b9b41aa12e5b7fb0cafeac70ec267b4112fcc95f0e1f917e8a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hbd0866056c4bbf101713f54405280958046dc1b7af58b13df2fb29da30cc8abf9e698cc7907e3c229b7efa0bb05c47aca8bbc9708b30c92f91932881676c6d8ba254b6e658151adbe937fe121c248fac54b9d45859de577a6f278a126adbc6a8218c7f2617663b4177b60f822e45964c8d2a8067859c4b8ed4484d62432fa23e16f95612bad100df9f6f05beed4e46df2ece97ba88dee5a16ffa8f8069d4540090abc07bde9676f9d6d5862e81fd70b96c192cfb9f82699157ec6e5bee7165babf3c862dfefb0fe284f83088f3867a8c65b6f2788496dedd07376bf0daf0e0aec586b0b3b7f788469b0cf46897984fb45f4e6686a995c02819f336b63cdc90d45889ef41d8922b8ec37730c0e0d694c408500722bf039a2ba46a15a7ae21fa78fe3e97dc9a8c8dbb2079d1b5116ff833bd6f9c794dc6c3641306d39826a7aca0d835fb96f6ddee8a8805a86f2318d37b00eecd1680a503393d1bbb4c1ce24bb07749a74492b6d0bf0c02542f8431025f2ce5ea5ed08491621fdfdf22b72994f2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h64cc1eda3db9785cc1e84cee916c5972d7d35501a23b66e415cdf4e3022d02dadb5fb7cef8c789fcbce47c173f92e3171a2cf5a57a8d8cd6263a0e07126d778793b75b73c9b55b3246c7ad132518efae79b9033754e776fd3bcc540cc4c1f385f82fa1161cd334d0466c8885b32b845f5819997b30a181479213bf067088558e74457d61f0fbdab479a0997c18b993f15883c0f2f35d6c6e2d93593900719f3f134870994e74c90fb0ee30dc97e6deb00f7ec9834259915601cc1a5fe99e0bd594e817622c351a3e171a2831c5fbaa30ffac4cf472f5c0e09dee5b8dfe5e1d72df1c80d85699bfd05197c8286afba71b6163e775f5c843ea5850a80cb820a3a755aa26dbd859cd56f839bbc15f98feadb2fc7f9d7349f322751c3cd7c38bdd58fac20a48a02592d236d267001fb8b55f81fddcb2399c76c5b15fe6cbba9bc300ee5cdbf214a05fb389e9b361df94a820a610a7bf3966e756b9534706a13fd8397bfeb1a6a697adfd74ad328d232a7736e39b8b4b6b49864b9ef84eab2080b3b6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h45b9166864710463fc4db11b5dcd5420471fd50d2e59fe15d2012f965deba4c20fbd1e77ecfe6d48e20de398255b4bd4125a3c56c5a281d667027b6e6656f382ec5f9ab6b46e6b56de6573e448a8262a591d94bf5566c45ff258e567c1a3ed209b63d131d6e7dfea47a89b5b51e72ae5dc986b362d7de92de4c3c1dcaea0bede968d0ce6e81ba96e17d5130a4c4e02092adc80355d76f77d7f89e923a109993c2fe003db142c18cd8805f0c454d94fbde47e04225e9bef247067d6ad26ea86b7079a6943c38e2e087bdfd0cca42806805d24614faad539d5f9d077684ab80862ed288e60dd2414f6c773cf21f2802cccd5980ffcd3cc780bd6d76096e4a330992555a6a781e5e4ebeea6d627e09b0b4542819a41757fbc39901b50e42ac59bc257597e020e26f05541c81636decfc1059b26ee438f3486e6296da4efcfe78c7ef52da82df20c6c10ea5a9a0468c4bc7e36897bae9e86dcc1993aae0da773f6b84fb961e15b4236952f277151b55bd553d7725c29e9744a5df63b5171604783d6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf5ed4617e0df7d240d18e888a3d9641a891ce14022a776e06abb033f04433abf21f878d89399acaa8a0809e247033dd4fc905a155902e3ae3eb2af54eded880c123f27329b8d8bf2be785c3e727fff63ce5518b126a40207380fc7a436d0337f0bec4da3f2ce018957790395860ef5c5d34778c47def8c84c032e10993a0b6181d0d5ac2d74ac8503089f37051a120632ae2a241cad837c428ac0b5df7e4fb39dbf9822eabd6c1180d15c0eb64e6f3c79383b93187e69622f7ab4e0de6b7e74c0b85a693d1ec06088fa02853a9f528f52fbfd7fc5e2ed866cc1c0f1d4b39d6047b93b05c8da7aee8741f2b01ca51d8fcecbf335cc563375b11ad0364e9390bce9d6f426d19b12171cd20e96fccd7295921bb9a51f66dbb3846d0916548d5822854267fa331c6f07a461082ebd4b386e2da901deb454c94254f2943596191e7f20c5a6dc7b29c7a55419102f22cf56c3b067a728ae6b308c1e08c05a7c192661343711592ffa7b27e4f2467c071d6a4916834022709821cf7944967a64e341e0f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h1ec8a66f17bc802db336bed0da72c0bc2e5c3ad1e2536b82bf2511cd40be690160e5f695bc1c8b990c5a09737d0fdacd187fba2fb2262063b7b5a2b1707cd75d1715a03be7b23d46bc3b2d34aaf6eed60c5a3a795eabcd97ba5901924f4c7501e38825ff2ad4cd0f96133d00c3128efc17ddd677cb702c3fc50e50fe2e1df2cc95d58465fc7557736ad5df5f44937ade229daddec57cc271859a9cc6d029963c1271cda92f1990907054428629235e5630e846429b114d3a3d0e7d172ae11fde104f928511f73910878ac21eb79dd525dd765b9f6f0a5ba0e6f7e76f4c6c7e6ef877bea90873ba5e1f6b47a8a50289d5ae6193e86894e4d77b690854dc4d72144773a96af1f9a11da0e57dbf35e0f5c271ef1ce5a00dd1113fa7a7832472757d20dde14c16a579a7cad09b66396e6667e46ac2453074626d6864e57b939d78bc527ea746765ee387b4be5f556172bb79a012efb9376dce7cb48c21af1b08d2aa60fb332b9d7d6184aed05a93717292ba1dae3cc8713c7773b498df708e289405;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha24c9a5b1dd522267ff544831a04d5de959d2659f4de9a3ca3c5b2eedc230b79ece3c10f00d18de234e40e00fc3272ca018d88718ffd32b8dca67e2aa9a582b03b7795d1107eca6a27029a433991648585436898dcfa736319422447c2d4a8a33794425b9026bfe7c8b74f7d96988e7afac9ce4851cc3e4dba855b8b8b52b81277d87e52e08837b176051c8ba3a03f7dcebfc24874328264ac825e73d02c4980d1d9adad8207c724f28c7cf70544e77aa7fccc84f9938fd71e0248febb118bd543f2d0854675b5112f20340077a35e96989749b1a9771d10aab1eb62b3afb2322f2e235f9231ab76ce3997fdd9ba9f30c42038e66c3c7d855b180769e1d800737f7fde1b3ac1528c60e57517de9cc74b874e8b65c3f4d15c6a977708ea33da2de48029146eb45be996feecb1cf3b6f0bb07c98af34025c1a1a33a224dc881126670feb27b216112ce96b4336297436adb6011da6453d8b99f017b9d8aae16f4547048a9995d16f9967b8e26030da1bf1e055ac6edd5a6adbb1ed6e3f9f04545f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he308301546d2c842a307585e82435a608d1247a96f5457161168f5c3754c9a622e3e2a1fba810d957b31b0f0ccd9e8bdb7afa23d2602cb5110ed921c2bf52ea710a79207c59a31a6a84f6ae79bf2d7eb771d4a10e09312533f9340e7696eca902f35b6ea8a17e66dc8e8abaed8adc493103446846aee44ab1c66c344e93ad1491c492fdaf0a1de96f7a0873e367dec5e05f775984408851d94628f8601c4af4eab6c889eef16089c678b3a1f58a76f4dc8076924a32fb02b1f81d165e298025217f44b318256b3a9587d9928b18a52f89f74da5c472f0d864e772fd34193ad0e6c94a99df8a8a31149a9317149263b7edd9c51d7780b1bfb27906851c52abdd5448d17fd18be3b88241c5781853364e19f2883b4646e6f96fb2ad646a11bad53dc11b230153af78164516b9f8a91dea194cd96a6c7d04e79d1cd652994b9ae08afe83924320d5f5cf5386f5fb33a026236e6d4ed84f97ccb99238a67dd4f69e6cfee76b96d0b877f98adcce6f7a3e26dcca2d99c2ea4c1efc9409e15c59dcf12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9a337ea0d7f3ba00bab794b930657681c2053087192303a08cefef858731dff50435c11206294d93dea3b2f32aeb835501057247dd0fa5e89e5e1306d8dc49b1f3101485c78a8565432fba37471f913101c6dab01092797d12fb51dfa8aa097023df36d21680d9acdafe8bb7aa7be1bc5c76ff3dc3f77b97baa35a27b4c02ef476f51138cc9048a5558a3aa44a0ac0a4cbb3286c9334e35cc556a642d280a4af0b0473d3767f8aa2a6822294c78c13e53f1988a0574bd326866380499fd3f9cfa6d6c65caeaf65fdf9299f8cd8b819875eef25c8b05be5520437d6be05794b1dfdf573a716b40848d01a5284d3b47800b6547bb9a62bbc8dea9b8f98620b12701709b086e1d2e98d45b421bb5b79193f96a0aaad768f21077e160053fe359492cbcbb0264ee27aabaf2c464babb8245b9971f61e41baf51de018177f5cfb34f9f59eee565a03287045bcff1e5b690698fb7e66a4bd2247bc16141e175c96ebb46eccdd628a200ef697d2a7da51fd0bf58757d46fd194733f92e74466a0a420b4;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hdb81402054c05cf99d8933993eaf5e551b6e179e4c357e71629ab7f6b1cb2b233c45c83d17c1d5d002d9556fe05adf5d6f56ffefa718f7a35fedd254fbbc79b8a892b3e79489290c3208126b4a2425aab14c67d8f96d3ecf0d47e9fd3be303ea3890f35410333b261d1fa81ae98ae4f08ec7af760bb6aa9e646911f7c0da298878807dec047a9f851b88520d6e28ffcde8fed6cb1546bc75693ce8c7cd6ded8733f66d6b9572ea60ca9265ee884b18c7d54f654fda5c6ab30a6414a3e7af0b659d796660307cc61e21c883c7124ef825b90873ebcdf668e1d37feb7453810b3cb0aabfdb181c3f844a4506adede063fca482a04d237bb4988cbb9a66c071486fc64ed44a2252d0f787a4ae6f66645ab52233e2cc1684557b101ef13b437490913e09ab3fdca091783d9cb0e16f08ae68f5f125572f2f32379350e624911b5e863f5771af0155cb92c4a66e77afb600cd931f5cf8266b7a753a6f7306d0cf3c7414ea0f02e6243b2a1a06103ec185f1b8c360b30e9f315742b68fe532aab1a39a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha9f20c429fe0bfa98877f6a1bc76073b5a435bc4e0e520b3a91ed4e15bb0b455986338f36a4432c99a600780e0ef56a7f450de563e9496381d1b66b40bb8e3c5e85ed24bd2d79f045a02936de275af258e57a6b5ec8a99135b4c9fc93006fc56543faed61c201df748c8a1206c7bddcc736a4fd37fadf3e58ede2947886b48592916ba81546bf650bc0fb36d3dcfacf0cb5f1c8ba833f65452dccda1668081f2efd3618bab934d636e269075023d210e1064ce5f5532286b2f03d31a49efcb69f3671440f57c536e096352b3b8c10e5593d5f6f0b163e3eea226e2b429797c30ca3a0e89badba93fc4439036eb58197e0c2eb84b3320f131481e4e20f3ae5f01731583a87b8b8c86719cb592c6f1753def80f5b7745d725383671003641f7ca834bc0da5c929bae6dd0569931f410a191bb3b4ed256d2315e4e4a4113ea22f61b42960a78680d9aa761f84b1abcf301cc28cb473a6d61f8f52e34d2217b2a56c22929ef95d0452dd86abb0cdc336a91a7b87a4005a18adff00a84d5693c75fa9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hb789ef3f87cf2489749c5ec5bd95f0e86091ba96de4c91dd4c63b94647813594453bbf53b887e1c7b9c2f427d12937971264cda98b12369f4819b0635c504e161dbfebc48a7a5414272a1370ea86de7f2c64db3542c9a5f9791af8117117d09335e3babfb115ef77fed2bcdaf8c7f036e26b4885e715b9079523d6df79ea507ed2542b9afccaf744bfc86969086f1919f7af774a8b150339614bbcdbf75345c00d6d057c2bf05690458d12f59f2103cf0599564fa121d27651d4f5e4242e861d0e6a3f7623203a0611c2410718ff838a2a3d34772e7f5ce689f0419d3b1645090ec3019836b19c07b6aac2a14af9ebab9da20d677d150704cd025149ae3b59aa0fbdd4aedb0a5698d6a12e046c99e7dd786ebd3511a81c3e399543e608ea568fb4ff288455232041495bdaf5454eeb53fba524f8d686433fb1e62e97ed44d1ea13732a4ca59d2a740ff4e19794e9120cbd6e45d44e8c383fcdd98eb4749504748e11afd91bb930527398db50fb3395b7e31ac27ad05826e3de189aed07d8f75e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hefdee6381a7aea9ca2885e4fba8b561ff5d5a5c1499836b8eaac0148c5c6ce5e79884164f31a1f1abedd6afef6505c838de9b15de9052f1e9741459a50d428eb518bafbf41294381a25d766b524c1c7047b87bfc7cd94be17f04d6e411dcf1bda200468891d7e05603d0fea146ae3f3b5b70bc4dc9e6fe9ca19d86691bd617f62a39e81e66a43cdbd58031ab8b097a111e1bed84975b556a14ac33367a5049577f70e807965237fd3a0e403f74538610103886adef567779740f3348c98de600c47fe6119f0c7868752b78e5866c8300036e7c71187b3c6bd2bdbd1bbf76b7fb3ca449ca8e698b9bd458932e1899b09ff01baf7057a6973f28ffe20123b9d81cc312067c8cf23921f2458b0941c8a563c590c4b31caade3597021027b52a04f920f132b71540768b6860d37ea62a6fa42e2195ea025bd3e7beee9cb9fe219b8e19bd8d28b13b3db0ced7a8dcd6b20f056ed6e285a6ab76ae49ec20e6865fa122af661702efc589c795fef00e9f8f81a24501ef091523cece198822d918c5d0fc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha22efd20200ce8f4545d7e820e56cfa6fa4042a43ff5adec14f1b8a964e80ab8cd7eb6fce3c1704b3a2affad7a728e75b65344727c8537bcf53b286c1d9934229e73aa3cd16446ed60a7d2af08ba7ecf73a4fa36763830a47dd7407350a95395a399e9a06fe489d8bda79fdf44e5ab454ecf59396d35a5f8c69b2b31b3340a161e5f254a6f0975389cc1db003e81a5a657c9ec29b9e2c7746a0b79f5f80502cd64ee7c9b0c2176b593a2df0604d7d7471bbc470efc14c21783ff6f1efc62c45f25befc9928eaf63bd801b4e43e6094e091f05983969046c85ef62cca1ae62e822e8064862eb0a07721daeace497a1bdf88c63e2b4531d2a97879ad3ebca0cb2dc3c27ff70ecbb39c85bab16d7c5424d0e82f56b770453bed383fba46de4598b5dae681bf9684b83d25e018afa8061012d0837c92ac76cff7b2df9d914fbcc001c7037a5045f16f4a9c973eeb2bec531e5b5ea009c5311adf7027e2a730997b72be92918d2b37b13648499fc2a9bbbcc0caf02696deebf239e2d3add9a8715c4a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h563189755645d15fc0bf4aa99380a9987ea081f7754ca6c93a0c9a4652fbe1120606ba2df474a30f8eae5cab557f9cfceff599fd074b066d151889ff0d70c9692890a0e83e56c12ba2fcca138dd2866253818079ec3a07aaf94e8a54be31f65cd9dc4d9e518c2a28c4a54fe1606956eb190c23047d3e0082665e0685357bb7d5fe4c62eb635e133d1bd6eb9451d954c3f5b09e37ff6f8d0690bc8b2f1a568b4cb129181a009745a0360aa3265646fe02db4e10ed15dfa955e6624f7f2560e9efb7c1c1418fa45e1d4c27868e888884850c03096ff0f36c6518e498c1bb91fd8f38cde5e65a6c772f7bc163e6e015598f438a9787f2674259019beb7492450ae8dbd771795537046060949eda2fda92f20a4b11cef17e17fa2e9e5bfda29eb1b8b4a3e071ce59fbd8fda859cd4463773999b609e13e35f429cc930d02d395977b4cc31b4bde3b76484c2d33750c9196d2ea49b3b3b6362968b815884980bfec300a2c302fb09e6df76b70503b778cdcc6b718ecfeba1528ae3a23b0beb3368fb1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hfe0347dca72c92b6976ba2df406b4ee74daed13ead73abc01ffa264cf0c356863211d2bcc15a20a4f4474cde6dbf47f49684738a71d4f4408fba5a03c5457a5e8db3569c17ca205c14412f31d5efe72dcab7c66938c0fe6eff1d60f0bed38d02fbf5bb851744d1fb44a1d8a35f4c68e9c95ee47830963f419beeef8d5b6137c77e8f04ca60f06c48c562fb52251709fbdc60221b6622d1e75eda98c23708a2ce23e19df0ee70ee4114bccfda4c3cca08e936900a2018e38b500f41df264ce9c6252bfe626a99a940d815f1eb8eb215eda535dde5b2eb506e8376703addaef9a6be2bf655452a73c46b11d6b24a4bdb993b54cea1e85d1c3387071332df6928e9e2fd7aa1c228d0515cf6fd6d1d118c705a8f9effaf2f551d4207b42462cbc62cfce6dbb4a624f8aa6ca2f1b96d5c2c62f84f082c7aeb9e366df30e53aee8805cbd7dfe1afb8c89a1c03832c82643a2982b91a5ff2c0204e48e9190932dc91c651a1c7bea5cb6f16092d496fd4f5dede37ee7d71d9f0db613c98a01fef78596da;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf7dcd44819d4360dfcd15c528c8f89ab1c1422e15d494adfe5a8671caab430830f78a966819b533a1681b37c212b6b3fd8add3b7bbaca6e6038cc88f0d632144772ffdc049ea90056d1743169ccf185fa33aa5c9d3d50658a0c408269bd7b5cb43cc9efd3b3b57c4a94cda06f796b3cde317361e5c866e405fb06b5eca4e93aef8ec87172644238acea9fef5c0bdc9e5b3eb6d99497eb10268bd311c6f18ce3b56474f65cb690cb2251b310a6d028785d2f17ea9f1f9000e123ffdc31a599c4df0f4160fe7449545f238282a9e5395bd2e2573b6049c18fd81c4a238449e5906e6478c6f2ccc4aa0de357a90305eb6e06c9e359c7df336a483e0432b641a53cea099aa0439b3ed5d8416bb2f3124a47db3af718307349562785b7af78d64cb488b9745ee01dd64398bfe035cd81f911691ee41e5b074e0cd9bd69d9085ee452203aa67a093392d22d43727e0e4ab53e205d2ee2ddfac746f960d5a9a71912f3e43c498d2188bf3e7289cc09712f1c2959e482b6974d3dc4e2e5ce0c084b5e68c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h6d7738757ad8d8911ceb0859a829b25ef15dc191be416ca2cb54147ec48e1f1fbfa0067685f982eaa62b61b52ac793b7e20369ba9ba2bbb4a94f6f694e2ef6d4f5bc2cfbfc9ed231cc4e1193d6f77e28b120488ddd788630bb24d0504018492d9aef7a1f0d9931e04c182350e46d5d68f605b9a44bd14629c1805e1add1e4243a66af5bbbfd55c442a5d85aac247fd0c4e692a25ec0c4e898fdbc2574479d84339cc510650fcd681d8db9f78ec75ba0cbc7055d6d66fef70bb1f3b79c5314dde4c98391eb8c7188647f7d73ef1db9e7f7fd1985078794d5fbd7998ddac80dfe5ff74315994e28f22ddd1e0594419b9a265e0d1bcc8aff15315cc68bf0738551d4a34246af84aa6f7e5b29e1046a93e5f0e413e4e46b30866b9f5b21a0079d2921d4cd67236046a8722197a999c5bb71a672a9af9166506c89fb40182464add911c92560caf20c8e7928e5c622992f5362d20d6c301df3589eef9466b9429b19936d1d2dd4ed9c1412c1a094b5b22992a3aada85d68cc56d426e76c39e5773706;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h25e6f8b3ef6fd4740ff5e7458a3a3702764fe3b9e333e219fbca30e36a84366c1fbb98d066084022a29979441bcf72949bfbd720d6441957ce6667bbe78ac4d0b18104f64d8fb53e2d8836eb0b75d9aacfdba530dcc71bc90d571f780ff50bd95ec69f1fe8838080136361f63286f02fb16e6938f08d5757a17a53b66df44a87bcd4d04894a04a5a39bf9e896c434f50782a20623e801824ce49c684d2ecdad0b7ddc00a2682b2e74e713184a818e174ebe8a31f9e309195a853a8b19e86550717bd6b3140da99879e761a1884b1a87c676de82bb64676ba39d6c83c40550b15d7960ec0bbddceb134cd2164da1e5aad93fc9174ac98835b9527a71aeb5b9dd37da33c8ae3a352f0809e31a4135a0f5fe40fc69ab395ef273d5df709002e085d8c0005d847a93a7b950882c1b46bfda9e8ce6d0f5f3484940fdfd671b565ea256e932cd413f647b0acaf9e05bf42d79e83dc3a197398183800acbddbb7a174feadd32481218104efdbe0b9c4228e56fbf0f2fa2e21cb9ffa099600a12eb6c607;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hcf6faa8d148b276c143ac5d07e0142dcec84af64f3eed7fd527a98a910e9e8dbe9768dd9200fee73d7234af0987d5bc862229c409dcad6369aeaf94747cd57ad2b24f9f05597fd54488be12791d90ba1abc136eaed1e097d08f5c0e834c0727230a2c29f7114aa401529f03d7b9fd244d9df7fe46f4ead0dde057cd45249843aa4a764d4e2e23b850d1a5a69aebba0afbc5fd79b3ed57085c8c91984aedb63756aaa768d26e39e0db7d0287c589c2659bbdf53540816457866f33bf4e6972f7beb4d4ed3f75bd97a860b2cca7a47db014bda4ea90b1ed695069d2c695cea8326c158e5d49b71f776379e1ec6e1dc5174dfeb01f28d80aae421705d25e5cf4959b1f1c52fcde7b1d832ef7d489970939e25d041204b2fdd1eea40a91226c21c65ec72ea1bd9eebc9a856bf475eee5d0d1b164b69398a25d04553519c150660d99e319258294c5432cfc3c46c2d482fcaa195d111544ec5c4479919b47ce8dc8d218e731c8404548b8bd81028c9360e96ec6df06b5227d4d06adf83dedae39744a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h8d2935ba79d4c3a5a145f97f02ba8405c3776361b5db2fbc5fff0ac459cedf91a3e674eacfc8c8473b8b1279f939c6b3c9e6c3844f6d449f46e57f149ab713b3aae3f1df51aaa5f61527984ca871100b16613df224d4841f85e98a8024fcdddc1976187207b80fc4320410f60ed9709767f907a9a22826d666025be82562dd43489a149ac8fea64e78a58465acc8c1ddb3e4623a14f6d1ff924236de2cd0378571719ba956eaaf9d38ac8bc0c3c8094ccdc0dd3578bcfe3b46b170935f7073416017fe4fa5b30bfea67879b2012044e91b11a88530b233bf69518c4bc361884e42c8e78eb59cd8d7f37e3e6d8c11c7a99375b8cf02f8313fb4256298b81d1c01bfd24522911b667973a020170f893e935a41600abeb2bb29af3251d13468d6be143fe23c33af55cf3b73740a477c0dc8d5e4828a041bf8fe1d954266c8f399073f0b737ffef3d799221a50a211c57c804ef3359a6085e2fbbd5cc93a5b61c297c5e05e50d13dc472091cba681faa725299e086b57965d0f83247240aa481287f;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5082d1eac97640e9cf7672dfaee597d368a5c84e4b19b8a9eea3aa280d4784599992cd506e9354f8296fa1423cb74f6d1b69f2308e7ea615cd96858e8f1d9765a5f83ce71900cc824f86797962f9014834e1f4ceb8212baabbbc8fbcadca8ff40a489157f5bd08a009c8a86154b9e8d06ed6412f4c54cfbb2e399b89b975b8e1d253831f31be6befd57baf948e27d033f969fc8ab7d37713d378b4ced56377c6e1bd7797f71219500005cceeea5b723e4a08a83db022427339ef685841fde999eda59c3c6120f03fe82dd88f7bb281705f40948a91880e6b1c4280bb16ce3739e38e9529df3629549fc449433f65a111d2aaf7c1453bb4375d4f871d1742602a1c8c4685edf2a27ca0fefc290c9c047f394fd080e015c8654783fb032d6a25e82451e4cc9725ed5b6ffa8ca86c73a6d3e2d233aade2f1ffa2f421762cf468bddfcc45cc8b8716ad08dd8902dfef15a6c271e6bdc141ab5df99611d1f6c629b86daacff334621a1d28f9d1b2a8cff3f77a3f1e4d6b5c69ca651c43c5bf7e9735d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hcc1c4a6350cc67b95fabd62b7e59545f1f3561364b81c692ed2a64b5f70c8cff9a452ceb696336e597ee92169996636ec61583dec9577def01e4816ea534469b90a404bbc288fcfb3b577c6c130b5649a5b7ec27ffe361dbe90e9722516f9f456087f37bb3c3defffc90d10bb73df8693a0f919852a7050006024df984f5fec7a97b18aea247394ff341044ec2c01e61712b13dcfbc9b628edf842bc989b1bff86802c16d404b46f9149092cc89d2aed35fd769bb97f2870679de2ca7c3becd7dd01ae8658f8cee85979efaa61ab00c23da79e39e4795bf80e8d6ee70883d9da8de0bcb7318a0d6bd62c22a1b6b4e8054aa64df2cd5e5e33d5bde5406628067de21d6b8b735b4ae1ba13950f1751ef7c5398e188de911c56588d04e3705dff1f271dbbffc6c81bac813c4e854ee2a548a763369e41f25f8daa0a5dea8d859e170a7e3e9d217963533e93b45514b9ae845bc08c37770df051d4ea96c11ab385fd2f2d8c97a25eba3b45a88988c8fe52fb17ff0880b04745051341768d37cae45c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'ha0ea7f8c54a5997d62187637f607b015167e04e420835e6b5024a0433c6c854d06c7794bc2703e52169d964e75bb1bbde04b6950de9e78a44058232c12b2fea2d1caa609e04793f3cec6dc8e66de2ffcfc03598af128bf335e020eceb6187b63a822001833131d30d36831cdf6f7fc891712bbb470fec6c6783fadb025e07c4e3cb8240879611b42290dc0330d9433b81638502bee80ecbe855b159f1fddf967d227829a76072a66dd6262827b32f5433c2dc637ee1a4807a58177112c343f21145e67c929dcf24c86c864d772ddf4a547bb627a18c7a5276e52ec6112a401965dca17c2980baf82a865a4cde9c16e669beab0f35b7b2448b044dd9cf13da736df000539b10b3c8af5bd7a2a83182663be65fe2d6425bfbc6fb4b574a97b83d43d0c3dc42274c8586257d8ff8cd89f195b6a7015a29889a98ca29407d08c27a8d97034c6d0561957fdc30938c84a05a47135129c94def0d48647ee8ea303ddfa30722e124c8bd6751cb3d281a8223934c68a7eba338522243a3673f4254e6e1e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hec568b51175f277c35c487b6ec7fa7a25aa2eb784d7a628a9681fa3ea673c78fe6bed8413ffbd6df0e3d31557d4783d5665f91f802401572ea43e5cbafcf51e211ad1f2c233adce368baf990607343c5f7b2d2c30c36588899cc650afb7974b390557c8a8704e01dd46e124b7ae2de2e808606475ea3dfc97180d20c6d71024026806f4c8cdac51f1c27132324b92e303812a50a599013ac564d9a8f8ab0f6c3c88d1026f935a0dc103e12c72044588d30fe8a23f485003f2b546c44829c63312b5d61cdb566e37f0c5f2b2868ae148399a524ebc22f03fd1939a53961bd5ae8294957ab10d2701250f205f855493ed32855fc673ed4f19a77bee253c16d61501a790c6cb6c5daa9fd662f76b4c810c9cdfbd58df8eac28baaad1c92dcd69898b378d53bc7383d4d99a882749431373e28654fba7ed786835157a04e38e239a218fcd40882655401a1e811beff4569efe45c49c9c2fc426af3827f25e03a8d0502c1b54f65bc8f21c1718c5ba28c2c169cc02db4f23c4e5a0094d62c3be19d96;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5b2e5442e00fadb8fac703c986d087dc019d3fdb0380380095e703d52928edfa74bf06636cf936f5ef6d98b423cc36a9d398d9dbdcda382ab174c3185b93bb8ef0f8e32f80b847d18544856708e2ca3f67953236d58db115b4feed411ed7893733847ee6e0d449de254d226d1d0cb919a1e2a496c1b791697bae45e08376b9968095b13018318faeb84bc2bd6cb1105ae9da32ef9c1950e44bed82990af7644472640580dd2952466c80005c7365d3fe9407793129917ef5ea74d37e8f5bceca4a9f890411a5c1b38d6ddfa396a55110ba7aadbacbf3f103d2f9bbab722c551e5cc04419ffed6bf2de397d5df828748f93a09a95a41df0c2e304f359ad899acaf1c55bd199864296222787d86a5cece7f7c773e69bd311c0f61d8208a341ab24bfece2e96db023689fb1102472c2ceda49531ab84718e23bcb27dc3befebc47fef27b5a7fc7f220d02a6cc0c48e787f02efee6c4c72a5ef53ab41ccd926a6871e2dfbfef0bdffc4f873f30e0ebe3819be33f4a0ba98ea872bf7263e21d41d3bc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h9c52b781c6a01638118db3f0fb9827c45477c82843001474d37eff8ae3bf9c95d485dc8f0ba44d26d5025e336778d946cfc4cf93a5b6f26561d46414662c9c0f5467654ec4338ee15160bf7c26efd1f249c7be3cd0d1afbf02c8ce5559d7adda868df37103650246d715775d491d8f0d7a232e3468e5bd884500c4256e67a925e2ad4cd3a5dba1c2cbb1a3e4dbbda6dbc69c7d2b5088c8197973cbda2611da172d9832ed0de9604340cc7f0c6bf84eb150d87582f80908847299838210941ce52fc976b67f20a79c7b398a65a441ea5db596b3d03611938acfdbb7033c14ab75b4c914a6fc293a7f17170beee52f8d3aba22a9239a8d866aa21f81e26baef629e89bd25e19a894ac68cc0cc37ea984dc3f076fcb70b777de1e12d0be1ed0518eb6466f1c4999ccf9c88f592868441002350b9ca28ce1be7e12dea23c82cea0fd81ab37742ec20a6d0c2013232f177d0de2f870996e6f5dc7dbc3ee7e926785014e23789001babad17465a79c5c59a900c68353500bf17152ce2f613faaf1d0b9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h861f84da412d67dbbbe74ce038845d393790f4466a2e3a25c6df27af9d3ae6480d97919870c935e0ca68e82061cae8e98f99debb8f426dd8b3257b49e3889622d07a3ceba60cb9b35697868481bb4ffa90915b21f0ba74c159142236fa5f8bec9110945aa252d8a621a86772af709a02bae3dc6c1fd39e598c9c0ca5f8dc4a3f7512bdda9d77575734fd05501df7aa696e7747b7a5061a2ee84663c53c330a8f0fd20497bdb4544e6894d1fe4ba9716514abefd3397d02c2df85a8087c8178d3d870d384affb72daabdd3d712460431e194caca6c344cf7cf9f5a2df8015e11da3c6743e8ea90eb78af67882d095938d5bcc2ef7fa15d9db5094bc22f1926ec901b4d27db87262ac4cb4148c51e6adfdc634c60b956bd5c02e9f3a7d0d5ee7d757efd6b08339bc538d870f1fc5e0e29048d0f187ef7b9b867c028045e9841e4ec19fc20fd8bc1086ca5701b63ab94091adaa8e56b670f38ea865368aa6e25310df0262a4888cd0c250ffc8ef490a86b6a68afd35d881ecc17ced7d9c2422411c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3d12253dd57bdfa4a6e09c87719fe1b5a9e2f05d984066f615a82573a3f0a3ae21918ecc0116ae0bd6c84e436570e32c25900826d49b214f4210e19b3c84decbec1f6a8e07b429fc9fa710d32b7903eb6e8220eafa44b6111d819484fd1dd959b746d2c623e912d2bdc4623d207705e3347d1bd1a5213d68841418b4c1700e1dcd33274f0a76fd84f9219dae190abb15cbfece9e8df351d7d8696213a3ba3adb24eac0b379115951c0d43c64cf00cd7ddb206f8a76bfef47066a595d2a3a2f1fff0637d1dbc0a8ea815a6706550a394d67271639cd4e2a4eddeb2726f542b549043215c1638a8f0a1c2afc331b936f8e565ab9f4085656d9bbde9ada5f1fd7418ea076e388c08c1eb3f57fd6924a8467d7947efac9c841c1a31e32f1def3146f44221b3f0230b210d3970e6a7f2d4d0e572e6434f1631fbf9754898fe874f1ff67bc364efcd53f035d1a6da561ae42d0534b53239afbed495db811cd122dfbddc43a9059a4eea84465cafdff43047bf12790f1d0d19f5fbfe7c0cbfd56b2b0d8;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h71d192eda3ffe509dffa792139770a4f29816de3baa87956c25d69296fe562a893d662c04cbdb41b7c75154b74c23f0ae45b846b6d832f4042ad63fbd6dba8c05069ea369fa7a8d37fcc76bb72b57fb907dad61fee8ca0621efd069f96f62736a05f4cc398d987cfb94baf00d9e6a26c1a4a7e612a212692cfac543b5beac5bf51dc0b8c159d7f2b33c79a2eae466f70dfea92f619a132a8604a7e2a6fcb503b5e1b5f08c75e4e402e5cc96f1824f7adf8bc80aa2b6e8c6f974f5ff80854426d2f22a5f7eb50d9dae694d287e02d61197f45aa2ee5c3b7350486b8dfb56506b84b63704c8154a04044cc97e3018383225a945a7b27bab86a0a91e45c963510ac9306f7f1561d17bb3f13cde3af653f7cb4ad416a008494fb54c6043a847a4d344af267744f04f487771d0ae227dd42dcf62f462de7ee8d8bc0c0993c9ab3461cf715653167e8b76680fa16b0507edb0197b17f958e260882a099c8452150d0e4d0f13b761e69b8737166f90beaba7174ffbe92d35405f478b07ef17b53c9ed2d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h7c843d7afd7f30803bbf8fd8972075ad0109302a38561476b519dc4fae8d032a1e2ac3dc8a0fb29b0e65c1b4622b088c6a44a0dc6aedab321545c42d8b5786ae640d979aa41a4ffba29013e05ce13886817dd04639b60d13f7a107855dea6c7e94f996318f83660b49aca2339163a5175fd99c04f822a7e238f49529d9d9954fb7c5734a64250452a0cf3dfb4758499aebd15045bf9552e8e8044da259194447fad99d594f94cc828a76aba072d36032c3ec54fba903f9676dd959d3a9786f9f2061ece78048162390ea686d947a544ec0a0e0b8c3c55a445ebb7e226881777342e328c8021f58df21fe01aeef23054c9a8db82a894c9fb487f3a3edc7a4f87c7f7212b9cb9fc51f523c2f527b6f9cbd4793ec7fbe1c2c4320c4288b7c0e8683b2fa5fa4c5c7fa5f377ee322a3bcb6c2547d44da3c7e92ca9105a232a79efffbccbea0fa8d90ead43466a0177602dc239297d6893bcffd670883108a61d78943708c685d0063c139049ba518124ddfbd23ccacfea63d6d52260af2add353947;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h309eb51ee3cea5d04e2fd263642478ab6a6e1dc1322c578bde2898dad960c9e421e3794552596a22e5df0ee04df75da02826bf00aba961c3ed5a6c496957c01d69b92d04e7c2580b94861cb12d857afaf41e785d78f9ce877e9f7594a57760d7db01e227f7b8a4af2cc3ec818379c527a28d272207bdcc27ec8bfd03a5458d162ec976c961ed415ceb00b785786e68e288b88d16993fe18102f172c308469abbacdc824287167718653fff9fda27d7d0b6bd47ab622a93ca4773951064f8a33a26b1a5ee53900e4ddcb2131ed1d23642ed7675464f6dc2a24ce77987fc697883937bb4556cca75f2845ce9f2fc03b3558aa7e9b1eaee0f3ac2481e59666605b611fae9c176f9dcdc08c5e2c6892baaf0ae2209d07833a488dc553f6e7c007accee4e9f07e79b0beec68a92d8f5e861a31384764d0d595923a53ef6a897f1067952db3d2a8ae52dae398cf0e3fe2f4159013d3a7d70d8e9db5468f9bd275a42fab8c1b4e15b9af99fae6f37c03ab1aaabc1801e47b8aeeb9b876aa1a264e33765;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h37f97df22ff7771f1fc2f27d787f16306b0abee157affd6514e7d661e1c325187100d8edead2fe8af5c92e76729e8a11efeee6d3e68fb59159ee297378851ff749120332571bf587a1e305cfac4f6094b541959aba48fe04fc9684508f97caf5d2b0ef2ddb67f2649735c640a672b9862874d6ada8381787458a597e5bf9c221069c66341a37760fb6c0a8ee28912d1ee0fe24dc20536d77cea22184bfb9c837e3e44191de21a8a7b8ee7be83da195b29960845392820b53ba514ba1c8bb4ca816da105dad1a9ebbf5bc73c2fa590dcf5c965025bfc70ddabed9dbbd2216f04d77a22a69c4d6f008002744d5e584c3b533c887051476cc2821627a08ba93350f4f1311e807f0f64792be32faa3de736ebca31d5fd0e796ab44388b35696a36d811774104c10a6285d1b095123a5bd822fc796435709f639a522f17da99ad6142795170597166b408e7c9143921d534269cc970dd4d1f4bfe397cfb7107c1e4915a42f47c346cf701eb4555e98e6fc8f0d15c1bd479137682ba6f8aa159b29f12;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4e4241b9391bcffce655d793e548eb1d73db120c2d4f40e0382b6e8b159c34dfe9b879f764c7d8e4f339010cab2acc8187189f3401bef952944c0efad2892c6075e260faac5c59abeddeee176451aa8c7418eeaef2e310f25f28856706214944d78f884b28880e03cd183927d3a63511957753e55219c7b5d873d207c592603ae37cdae12b94ef33d50e4c0c27355ba645ad135a9a3c1f829dd79ac80fba5b8c9b613c6e609f5f3e06d958028b2f2a3b4249f53e4ed21a836d6bb2988549447a45142863eabee7e8514afb6c77c17345a004cf0df7d62cb78b2368d064998870b7b91fa53b8da689ed1ecbc3af9e8ef5f1afba320842542f0ed3e31d8d6bcb206d39f2642336b1cc1fcfe20aab5c29427e54d4e629e3dd5c12375bd465b8301a4b7178c60b2aadfc95bf2a178fa2b6a70ff809275471d97b3cacf3575f931be466aca7bfd057c20da206e82ac3eb02be0ae4423969b88897421b91d3f9fc8a883d3a8f05bfc8b86d8f8c17e6ead76a23b37a363d85e27e615cf3a09ef9bb3457;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he0f77bbc4812c02b21b3a3ea106577ed9804817c2cf2695ba20cee22c573ac96c39f704083ab82014117f559199a804a0be1b21a7f676cded7c81cbe846d43bdac70fb856163b5418104069e92afdb9c63d5d524e1918a1db7adace153b9aeb3f9be745111431ff7c9cffeed53bce304afe5880f2cb18a5808bb09dc4f062c074b4293729672cd5aa6fcec70dcb5ec42468ce150a82b55f263f92f17c14519441bb81cf9c039f953b181c68fc4721cbb4dd7aa47f0fc261d7e5399649c04d163c517bed0faba05991ba96c928c28348b50d2032e3f578554035d78562dd91eccbf37dad77e9f10726bac1cbdc0b99218367eee273ed07938e767a583616166d9ca550d861040e1aec3a2075476ecd5723bb1664e3eada30645e5e5f0f6dd63f3a3243965c8b7c0e6ea8a04d4acfb08cdaa0e00f91af981fa675ec48232882d6300050f544c09783e52a5b5a9df09722d31adc42b705a3b30e8f1658fb8be9e220fbb8f0f6d1b66a7afbd4552dc7777637b34ba76e768fa4dabe4791232d64c1b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hb363cd2f396d535b68ac1a2e18343c03c7ba2c70c9b2ae5151bf1c9d485de2ff9e03342a176c5d1d82528d4d4510129ed215a0d10a2c580401ed28166f9a4090677fe4f843cb9c610a34c081d1b82bec85cbb94a4eba54692f73ad9c5e3f9f7f0711a7c1cbc4620f892abd77747ca1c9080c730207dfc860b7fcc8840f1892fdc0d80bd4c6aceb83b6cb6b782c14aedac10a89b66cc80c11b8d428c8f0ea4a3a9e8233d657d899ad53ab885e7a3ab3e277aeeef0e5533bc9aeb5e7b8e825a758a3a4be64edea8ca739047053b34f8220733e12181d0d48ebadd7f305c4bc39bd20c86435d39d2833dd773ea0bce691cebf0c0d11427ed4d7ac5039595b0cfc2f5d8b7dde0d4576857a72d38fcca87a597bdfdccf1f800e9d57459e60842d8f9d09d6a63cf1458b719bb9edd259e998012b5c7137688a1420b43f0417511adb276dd747b5d40b1b1acdf4364d322ff60a534458dc8b7dcb19b1890e5496499918bda922eb3631a0b3e820595d56901cd6a57448b10315477197ade2869bd648d3;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4ea5b956f517fbee831132f374a48c6601d8fc681c6700c8d59aa944c67e25eee6115c2ee365be642682586167fcb9932425af64bf80492239e1ec1f231613d60fabd77b85b41df4913c34d6f1d417fb40ebe2cb0ec594b2f5c1f2b82b99da6471837c428c5ef1ae492f2e74dc0f8ab181f6f36b6021add49c648611eb666241ee388d561bb5b04b9e273803c806451f66def4a10a7d7e13e81f94244b98e15d0b4d83736db1500772975af4e7a48fd9130229429d233499e2bb82adaad780826f8d130ae95c3043545ce4424c8f51b0f5d368250193ea96392bb6c7035a39b7ef8b4fd807f43d87aeb8fa25ed417e094e44d461a43a829b5695a3a2b8cc8378c7c99ba3f9769a1cb84260a5a8e05288a5d092ffdaae59a501d8bc17e6fd2c1aba91e878b38652065ac2429d42258b9edcfc9f72383c3237bcac5346525e0afb4e5feea9c59d806c889d91a0e082378bbdd910fbd77d1aef20b5edfef734821bdfd524d33843ab141c72d0eaab3c0af98dfc00496e7b037cdcaa1d57b449850a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h7cf8d7933e175ddc7735006a1d27256b44e9ba0bd32c431ee5c960afaadcbe9b5e6c84a3d5f193d7d8ed214d1f95c6785bef990e032db89b300c0c7987b7cbcccbd19cd5bc9ddd3e4d6caba1bdca03809ae16fcf0bb1f7c104f7e11294b92075acb40b39de9345ac32f2238892d7ca570ca9b0b958c5df9074406b0fb665f6a89da09deee5b4fa8b1e1fa0daf405ee15c04433d6e2bb056890f9d9e14e3838846f4586b48c6a80b35602c690bf0e5463055a5a68c310797f9236791e062df8e7d235c1d3b9b4c556d6a142e2451b48fa139573a6b328bdad2c021ed6095d24069c38532cc0dac0ab191eaff798d0aa1ed2dcfdce66df241cdeffc57a495c3d38d40168ef2540634336847fb3ddb44aa606a34f92361a1e761c9eafeb266f3b7b6f47efaa023767bcb7fe7104431ac667a59e716bcdbeff4bb618752a94e7d877a75bbd2105af0c434a561a11b0977ca1904b28ed9e1a6746c1c7edfaa7f8f0e4bbc154c7dd8521772e36f7832a2480b81666de9bc951d4a24c238f23f2c65173;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h4af8b17333d9e963d676dfc755dd507c40f6d0617550acffc47ed399ce18db23d65639abd298c7ea5f5e7fa52e7cab05c2a9eebd94ee049dd99eb8f111dd2740d832e03fe7c6b538f1b982b60f631b6be40b7db6abb2e3887a097f7ece4c564f75910be0097c9bfcd71c8e989a929ec0a9df0929cd7e55715cc2c2e26f7162f857b8875c753728e766e681402584b0a7959d118291f697b48d2749bf4c5cc85d14cabd52444b99a6c1461658452aeac6e295292cb3af98fa6e06d77b798751a9c69204b229e6503133c3944672b4eea474591461275e0d56ef9cadb14d0e234c5eeab3ea1da4898b506dc2ae3639765f67f76fab3cfbcc5a26ec11a3b2081663e68bbdd9ce0c0e602442e77424d6a59791685a3df0cab1d17eb35aeab86b6213258791c3dd6f7bc3619252445a2ca89d79864ea8a397f4cf3d70672724a9c73ab322673b690069ca61aae7167a48a8a5d5d43a11294d1d844cae63a64523e497c6453e4283d4a229d66ee7c10531f92697512cc467d2ada552906241ad885ba1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd3f11b0a5a27d912c18e11e67837adbb663e670d3b2f46cd6454d2a416befaa96ad013853309aef277cb3782230f620fe7a04037d283dceb640c4446cdf850dbae6d0889f62ed487d218478da689e0175de6c9896a2b886e2f61dea4c64fb1d588a81d37fbe740ea85396a78496cbcf3458f40f6744fae800cf980dbf6099a2845bbfbf3c5c53839c73e5900412c2d4ab67047841db12363478356e19573dad271e3ec55d3d1b5a7ec31d07d1067eaccc5e82a1a04e6e2b75b76615873756f77504c0b0dbf84955edc1d224bcfa12cc8467b5a68d2c94230ce4681b71348bd8df8808835591151802c334725284ec7f9f17a73b846286f9cb99e35b4c67c14c3d8c6570f6e02806cad038169944b4d26c1497b924756be43f82e2270318b009de7d713886561d8768e0a325b6e25484f10133959ce46bbf4cdb2b313a85c28585e4e446491df127d42d3bec8f6443256ec46de1db5c445e6fb54278381c14b48ebcd32b6befecd1d654ad00841ee6aeeaab3fd866c761140d80b56e0d647ca23;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hbe6dd5e96d58705d06bd3fbee363d5fa38d49cd95f2d4ba3f4055ea0f30cc2d0f5b6455da3b32dfa1e4873a703f23e41d1c5f438c76b1f678aa750922f52f4a3d43fef8e39982077c8e0073249c06e9bb544a7c3b1a77c34f248f3df40695d1f4eb3781ebc2ee60fc6317fe3952ec0b8bcc50ad983101301540b577232f578a297fb33a24e938343770df669680fd4adb55444f57eec9b18a7727b1682bf33337aa8dfd4b0a26a001fe466bc768ae4f547a573bfa14f1356f0796453f5014023419b69bf505a2da75b3cc2c6cac5e1a09257ae362aa68e912016ef1d82d8e155f19c0aead5e9fd70d2a9a2255590e7934e632ea7ca9f0023f868b7c68d0187dd350e2da91107d08dfc776638e57f16968c82629dde18a928fac53df367e38fb7ab99cddf566a78ef6d713d200801c9c2e9d673dba6916aae587909f6a2eb56970874999e9e0a7edb7f58df02b45056f88677062f91b9cc2da7ec394a18c55b72523f91b7d5f36cf579d8ba05d5b2e5cb5e1f751956cdec2f740c61377e998d11;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5ec682dde91dc97c8885c508ebbb9aa9dd8f076ff9ea7e4efc6e719d9eccd49aac6c9fe5b2b8d1a63b31611ae41246cb5424e4169f3251432abba08d8e86c00166a7de5f6f233ac7e9df6ac8bb255c045fc54b2207b3b2d4fe6d771deb2b8bae721da825d9acd6c7355bb82a8c3491a56fc2067d67e6ad914525107d3bf08c3956df14bbc7b4471fe6c48589dadbe9efa710e1711a59eba608a65bbc75db20ee7203fd6022e4af68de9fef471a9b14b3c352a806e2dd08e9c39f2ce378a106d25a4a16e290542b0818a5e3e80856c435d2323494763ca89175089ed577f3ac775d71c030452132861547458cca5cbd08bb6bfc92da5a02064d94edf2bb972cb75011c695f0dfb40ae27873dda9ab13fb73e2b16a3551a13fcb3c920bfa19e336dc260a8c4559da051bfb0196cba649c5041a7955e4a5decff92158d81620daf7428ed9101f2b5f0249df5834363f5615bfd26c67bb336af7e976bf79ebe57b5b1821e84713d60f9e1ba316db53450a3c4bd30608dee8fa0890d8f3a07176629e;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h5428d791a1fa1dbe447f2c6cfae6a3bc24ebf44da43bdf50b401c1cd6962b1b798f6043a9c982460a6de297ba517bca597d98e6987c2b82ef9e5daa594a88e592a6a022c1c366c989f242ad5adf3a05e30e056e42db6049a5e5f34fbe35847ec8eb33494c9748fd48fe6157c1e7ad57f2db9d8fc7c55d37f83226c6c0cfaac98df81c3839ad1315b4b4f2668db7470a1765e19c75a8f1ed13466e04ef063a0efefe1be672a35c7db18e72b36241797992438df63f8c4018a7ade385497e48c611994077cd38c4e8d0c77608d1b73e65a2808ab1efb04e65dc09f37950692c2c4b9898c0d0bf7001625c22517aaaa8239dc78534718880c6ecb2964948bbe0ce6ec59d41ddad72605c8a01c2985b825381e198abe50207c696cc19b49b8fc540c3fc660e4b41e40a195b3af432d89d019c5dc89a7933d444619e519e313655e3fee2e666b6daa4ce1f156a1913f5731ea95ec9c5afb6c60425ef2b45e4d5e23a38b87e508cee58504661829f48c093e16c2691bbfd74a59a9e016d355e8679c47;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h7a05b903c6098574e4d18f2c1f8ba24582942e7cb23a8982047c62b7a6ae515dbfd11f616225a9a83379b1ed5cadac11fb8b51cd869097ddbfcdd7d45704edb09b8b3be1d9bb3731406d93a6816d2007860f15c1da68624df88bad5737ffccd3415f99f82eb8685c7e5407322396b70b81f92fc65697aff098271fa336c387069cddad3876f5922fdd3a9d8c0ed3a11ffc28a7fa1ec9822e2569c23c1d66d965e095ea0c873ba45d12c0989578948da1ab18e1777cf55778d44ba2a6e7d33769c954f12a35a7a8d1ad36bdf1d6a6060f182ec6f774d41f4a3f61d0f09c1d0ba81d2aa1d5e1738657767add9b2fb39e4fa687164ee2561e8909fd131433cdbe2cc5b315b84339e94df5a15a5a436fe20ae13dae0619f375e36c8b089ab1af79995f30d4d11b2966d018acd2e1409ba2207465d9a3ef39337961870bf04b4932a4e2579e5111b72ead1cc6c45cf831488c12319482b4d6eae18033dd0307b34a1ae05747338268dd3e4fa15b45f76ec4f87b84a0486342c2ae9f2870afa77091ab;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hfa1c63f4b8ff508d7b94c54d6ac02fe0c37deda5fab2af813f4061116da30030029132b0fb82006585980cbbc58dfedead867c2b1e8a941d4d7d508e744ab99218d996a047bfe73412cf351ab6b4c13c974d19e4af635b32ce1a8a80753656da703c9e13129344893e5f97f5ca3fea60941b38a6c5e594392fcf3bf4ef9c95f8f26c8138bf43461f65b04a6274f6839db27f003a64a0489140d057b9e63607c05816ea7b4c1e87653c6a7451a7ef5d01d9f3655f5802db4ac9dbda51fe2c5fa89919a4baad5c99aa1cb0e79a3c65286912731c58fa1acdc26df27f2b599df6485d280b57add0e3d5be2e6de0a5cf29cbf33996c655332154b24a6d75d9777e73db1313188370ec7a0ccec85acebc4ac35d96db8760a535f7169aaee6c86cf57ab3ea32ded02a8371f3db236f76e2e447ead5fbc2fe47c75b1cf3883bf12c737af9fc3fef70bd9440b99c4008a976e27d8ed12679b48d0559e7f6ccc715b4a27c6e070970875604c1382f5b58060540d4976fa017a03d3d500c3ed74a0cb86175;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf7b0d8635f1af03a92f243194f47b8fc7d8e7518acc20bd276c93c7349b0e379ad9360c0c688a06b06b75da0e29100499c7919af76c929134e2c4476a5ea8e2f96b59a2e51a333f3cfb727946d44f2ba386dfd91c3e1ff0b8251230215975e52e67e7869a7ec02f8acdc07b7038467fed5c0ca8b056038f718acaef4b7e4cf127ac94be3e31f49d96a9795ab71557dd44bfc9ce7c38c7ff0cefaf1bde280519b84529775449de63dbb8765957963b27b7b3c9c96eb4eb8c9e3fe7280c4b0cf4c24464b1c9ed165fe05050e7dc0195dc2f099af7f525759ad55d6305e0f156208dfd9e339625d38ccb2bcead498a66f497980489f87bc4a293c8b987e6bb1c16dabb6475d5cf239ade642d35ebf447d38a4d66440af1356cf51bfbdc0408922032accc43561b1832a979a9efc209e4a8bd346aebc4a210e452c44553f6db0ccf1f804690b8c07cb5ee40ac7e01d864f895d4273675a3398d38c20955c6007b88cf10ba9e6480555522d8bd0d4d10f07dbcc2fedca58f3fe8c6984fc44186a7bbe;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h12ae82edafe5302fa622b1f2101de1bc21d90ae765b8b5dc689a83cf2fcf9cd702113314fc7e580a31c418b4cb6536bf8b3b18c3d4e0aa76249eada2ef0380af88cdb76f81a7c76a7cbe7594e1d99f71475bf4c06b2573edc98419b1ed717c21de1852f2eddb5beacffdbfdb787f4c8b67854dd719d891e184419ce669a726b784f911fe9d5a9ac48942ccae7531798f1542bdbb72787807738aaa9a5bd92226f32283055ee2619f3f91db6c0fb4ef5c9dacc50add28f85aa5b499e694af6215b13dbc46ec7b3625696113f6ef405df7e3c3405412caa0c23146ee33f96d974fb6c00ceb6445f015c0d409e8bf236a1af80010d51b30f36f667c3def4bfefce107eb46144c3207952d3f18b1fc7ad0d0b6a2f15bfc2314481757de8735f300ff600393dd3e6a813f0a3bfe6046f61777a64827376d29239f2db2334cbbe2ed655dbc64796cb29910b5208a6b9d5b1f89de9f3b1938c73ca366313ab21fd86475e08d6554f0d73f1e1619777496badcaf092b4a5a3367168cc817028899ece63a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf9ecad3a06b38f1f362fa4ea7fde89695d9054adcca54a7442bd308696973de60d0e762d5b2c6db66271c870fdcfb31fef650a9b0347ffb37b294f831ebc235c41b3ef76287fb0115deee640cd1da64c3c92528d715c8a6a00f0a3d948ea19b08dc80418170768ba8bdd157b7bdc382c47230b9f3cf5a0025b6af9cec34a9ee57b0bc6e9e5f5ef96be31ec4f6bf3158952b67adca97de6f328b096e343cf089a467f12a3e02cffd30678e15a3c67ecd98c0b9cc78d1955dc7a74a76e12b076638af0eb22b9b7d4c043b1fc27a34826f711761a270714f09d066d923cb3fd2693a3bf775885d019b5091ea12a636309bc97c9b1df35cb2d973ab3860cb7f12b5c8a245393cb83e4421173c1e338a3bb61f45375c485b7c833a2bdf6ae3440a8463db912b5733b586f3c6dbdf4045f71e1dfcc132f1f887f3195ae4aaadc0e0c1f22644d289521f5e0876c0f8b18af6b6c56e23ea62418ae4e4103ae462571775b142d1f12fdf46c30c313edf35f7b575368a349ef69e7deca86be7b5263aff30d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h411d63e6be2014a7d5210a5a5ee7af121579398af4bbc45eb1a078d163932dbeb99a36f1face424cbbde8a3d6e6c60ada714ad684d4e4b4f3ee94db68d7ce166d895e8f93e354bcbaffffb106450d60dea41d017e7e3a647d3dd00d0c1e305ba5aea91b68b372e19a566b2d319a22d36aad3ed8f4e90289ebe9224ce201dac1a64c68987a7e84ea618c39680d3205bfe6796e1cc7bb3804c19c4492b1924ae116a2d4f3ae7571f11c36f8db9885a96837cea6d58afae33abbb4ddaaf76c348de7244619c19bb736be96d5f770d2e52b0bdd9de95081d67cf526a5bad231f5d1f3aa38491f5a93cd9ddc108a9a8fa556fdd1d90e2da1065ab32465163aab654a099d5778cff2d1c5f4d3639d7281a6ca7a007cb1d60f570ace775f3e1a1fbd1f0d3549396e392fd08f3e99338c78953968e6e492f88b50f0f2240f0d864631aeaee6ce84139f44493fc3fdfad98e3266248949aecd43d49d0e99746cd9f6be7036104b9b92bc61d93444d18ab76f9b544b00f95a99fb866e2c7effdd3fc7e54bf;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h52f1b72b0b999580884723e0635f2cae877ee7679a3058104be1df7fb1e4c10a4dd499d011ee0109069c4c9490cf9aa63626ab1443bd245802ba8f2b2e77896f81ab55e00a099d5196a8c6b1330741338948942ab949c4b9709c76628cb3e83c9d6e962be420fcd132e14055309b1782400753016fbb5063391465cea590f46c679387dbdbe6523b1de5be8c5300f68e7635c0ec175eb37a67d6331076393603d958f2d5490b238262bc947861d08f5011144fed154e825bcf173312c4fede17e8318757842cd414eef17ffd947bc0d69a405a6aff76d1c856a3118b9866d38769705f9dc15714cfd191196a165d022071e70d342a6dbc6ac8269854b6f22ed9fe4f84539101fc39db7b51d47bbac68ad49ecaa8d8be5155cb7b41f501e5bc4dcdda0cffd8880b57694f266bb35212fb1eaa54aaf659ea2f2dd53bd44109ea4f9caab78a43373f8dae3315a5e68f20e29805dc33e16275279f10f213adc68b148b84adeb8ce3a143e12c9071813ca435c9486cb0a66a65e0e30b90eae8923a7b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hc09e0f67a44460215ea9ce267797cafc5245c6efba785554b5b20d0bac1703f49d098b8eab00e74482c6b35335cd21fa7a92511f5fae5d7f5397f3f0dc8df2f7e154c40478f604902091b68afb49edc4d27aa05ecabc17382f620ef36e3c86471a989bbdea97fdd241f32990226118f9823488f602016356c155f86596e577bab31f0e999250b6276e2e7d0425874a37865a3a0d64bdd7651e2f9761021cd7a6bdf30aaed8957bc38305acea981b1d73bd50d9c4197439b9e3dbe9e6d9f3afe6f6652908affe38f9b2486f75eec7b898391543501f9f6383fb39073c798634f6c3212cefe9303bdd73998d36f1c7c43a6fea09b58473e34e6768a3af7c028529dd717b9418cdca6bbefefab618f7f26ab7d3fbe47ca6ae0743945706772bff5e3bd5ef4902b77525d64080df2fb99ca502fed4aa6134755700df333a52e336bcc680e0ed2a0c9ccc46d7fa25ee53933f5f6a344172eec8cc1c2ce1841725e3e025fdd40087e6e1f2d42439f06d402bb252a23c15a6368c4170866844cae8e67d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h13fecf4d9160243c4aa84e6bd885206992c9ea54bde4986cc1863c7a849587ca328c723658871c59d9a2fc06679328e5b99ea3a32201005165ed24a69ab524e7cd387835c1eeaa17b822f07cf5527cdc5ae99e1cef189c5eaf6fc0507303191b36aa558bf63bafd7eeff70a2c24f71650b6e7d1f7c7d5cd6bed20785668fbdf63b468d90df4dcb2d16af19f0385bdcd0e5c7cce7ac8f1fb058b3a9b9ae6454612e11035af94f56847a33e151721658f90e14c9c522a04d57ee4d751e8a8befb0772d72a0416ce579eb6c3166453267ca339fc09c820ba8c1a0abb4840d3dd83a5b41aa4d9b092eb1649a8e7ec2f72caa5b195e2d4e7658672cf7dabc74ad943830c05047b8d527fb7698155cd4d33d1b6c20d41e5f21cb338fb10e26b4250b413bb9cc66e6d428b644d5968a4da440ecfefec3d9773d31050b713832e0954dfdec6f5936c6bbe17ec94e763b7c541ee7783c322453265e486f602c79eef109e675f744b3bea2ce23f6bbb56390901bf63fe1acfbf923478171d95ea8120f37bd;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hb5e7ec2e01219af1c60d349e8e679bdb2a1fe8d9e4dd1309a5a96906fa779c2e3fa3ad3941437ded4ba3d470abcd3707ed2bf9b6b9531f417e75cdc0013ac8cc2b3b492111700daf53e6792d71fd29e22ca6911b8707dd01a8d589b2be63ebac8daffb641c68b60e9a069aed6212bb2114f521fa268209742e7851973e870c52f58657555fb18d0a2b3ee17e17eda36deb8694cf2ae4622a4c8ae92c5deb60ebd95235bedb5e063c5671baf9561dcd3151d4b689a8a42feca5c735db3250bcf51d3e2a620821cbb4b6a672e63965e0cacec5438da8d014c82bf2d8001592f9012523d396bfdc2d94f5e15bb8fa21a1e6f58fb595183c36745643155c2818d79e5761dde1e54746511619df792f70948a76333777514c338c8f9389c94377eb3073563e3bce5ba7a335f9aad2f1730cf4558417cd34a74dc1648eb83ef70879a8edbc7b26f9e875cf0c11f573869696011531711ceb3e62a02c3037929354c3c1a82add5b91345eef32af34523cb04ba3d7a3e14b1faaa973fc3dd94cad7af953;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf3d4ced50d807342a5e8b14cd4c5502ad1c9a995906f107d20502df033043f2037fe262565523b98eb9c0232c3c83b03e501de59f756192be61a2241e1c5db8203809d0d7e987423afc5dc24e3163b0c12c62cab69cdc8a42c666aa317b384e1387fd7039897e7479a2ed995760acfde884889c7d5654147b586e88fa95bd6659570e2ec4448ddc308c26e3aaaff868c95687156e9b4e41c4e3bf2def7fe0c8287f92582bb5360e3380f85ef87b803a257855eb7b7608a2e039e361f3053506c6081392241f5659bf6b77fddf8fbc702e9865a200408f996f558a10c9b5b62b72f66eb920093504573e7d5b0a653a7b28262aff7affc55900be52c4edc5685b36ee0dadbec92c5a6cde8017d28b876e9706afb2b5c7637e770d3fe3f2d91bda5170cabf51f33ffb8b6b890c52065c210c357a1f23e3c9ff96dac8089d7bb3708fc0afc14a935e46bc0e3f5d3001e507b658b85d4883c31fb100ed40df8189fe83c5800b2016e19f0c409ffe409d2a158453b46957fa843b6b131c52933dabfa7;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf60cf7cc580dd5f3494e004b3db5fe47fc8b504fcafa22af8571fcb970456837e18bdae6123441aa8222e4896828dc66db7f866d5cd56d8bc21c2a4c9c2c2a7d5e791c003d61feba181e93a5f87dccaf1574ba88e6d6f279676c2ed6d3976d1e18726758c847820d0a21d959cba482382ad9a2a6e8cb22d426ef41fe1c9ce3217e351c192bb3f811eb4da21101a69758cddb849c780c673e690c5067b4772193f74b7bfe39ce005562acfb51eb8ad7f12695b735201da1f016dcabc862ac33e8246e2e00522263f8bb72880a9373765afebc22a774a0c0a8826172e59deccf09a3dfc3ee062ca9b55a2b5f8d11c2076dc5f2d72a563bce92a65f908a8c94814c44d6e2d064c6f89e4d9e8a316e14510877e4794eec4d4320b7dbfa5e338507880757b70971b5c7d1ead9039813c12d370f5e6f8da4687185a631a3710efc595cee67056d29067568a6da39fdc46e552753d7257630e62a134829070efbe95381ef44a472a2270c3ceebea4e04406ac2ccebd1f792ce2c9ebc5f7a40ca94485d0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h14086b1de77a9859aab9ca72d9f03972769ea7c5870488e6b40db544dc855dbf17a7a63d361afd307d1e75bf86bf8ba78bfb6fdebdf71a6bc7da81ac8b0b2dcacce313e3a85fc3daa4e7d6841c7f06d2dfe66b1303db0b85e16cd12937098bfe1cd5548b6680b5e14fbb52bd9cfccf6bee6221e42cafc8c6a66fba6a641578ea83f8efecf40244343bce6fddd168888e0a8f0d5fd0ad5e37b813e28c1c24186b8b7ae70db7d2873a45ff5c67bfdf8d673d5037c4ad9724cd9be469ac19c2ff329c35d5b8ddef6cf3fd84507297d5afde45ffa08ec78c5ac07106cc6b19d6748dadff69c0b2ae7d0d0b6a3ae252b7ec925934187573e60e4bb815fdb512677a166145b00377cdf580d3abb5e2b381fe3692168cfcca128818cecda9e04e729c54766e4cc34f40889b309c774279e0851497bde22804111e4b8d56aa9d2435c952901b24dee5d0ac6bc1ff25be7d670e7655c6373b994727e1a8d21611a471d2dcd3d6a9e9e05e3d50e5e02311ff31b12ab412ff41f743c58b826db8d7a475d6b2;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hcbcd2eacfb945965b1c807335e2e6cb2f5b9773f8932c649bdde3ef932cb286ab8116b30cee42108188354851d5808a118c4cc81dfdabda2d97cd21779f8fce23ba2a65fb1d838e5963f90f8088d75e8d84488c970891bb0be3713867b0242d4a717c7cd3d6bf11b7bbb9dab3f4f9186fdee38dbe556386fd9f80f2d10bb69b18a3333becb92ce578bc0bffb44d00e2049b41c70a8d9a2f0e1786a0a1081c2c240ed694c0bbe863868949871287a93923e77e07b37fbb270ff24f3564f8686a1eb04374bd1976c0d0e89768edd8998388625977abdfd67ac30d3bac32ecb74cbb4350e689a469f6aa4360068880620fcbd0822b9c0b214c9024c4e5e6773c7a87112a5d5764e8f6c9c43c482ee4ec85549cd72578cdd256f087549bb59710210822ff9a0c0b12f46dafebe7a9f7349b65f8c96646d3556226964d6b00ef639390320d2e7b0bdebd200f5b8c78758c4f721bf6deddcbe348aa264f5e3c060b52729b5e4d539c77e4c37df65b50a4193e366a0955f32702d2b21e37874207e946d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h382e79ac1243bd8a594bb8cf41dbe4c2c87b04709e9d54998b2058cba1919afa6c57d6635e933c57208f2270d993953934c50c59d5d1ee5f554284ab5ae3a0886f01cc9e275aa386e8a9d4cf1f6405cae0b12ec86701a56da33be60b4092a760048bbcdafdddcb2d9a192ff6012ce4a1b3117be61478557aa4b7aa56267b4fa2ec1853abd88c623cdf02203514678fcd4a5181873b4d99f7977e9fa6b97508366241d40f7e295c0a6bdd6bcc2f21c147fc3dee9c8d4b6118c118ef2d87f32635a96e205edf531c72b6d70b4ca6efa81aeb759b8db195a6b81cd1eb74d59514d6ea1b9b98bf7805267caad057743c1907b0e44351e70cf775966cb1c6035baed0601e108ebcdf60afffd1a2ce16a7b670d5cfb7e1d1b8c56990d3fb4ed458c3e5c75328e3f94b778eac970cbd77494c1e32c6f6305048338c3230dc9bd51d670466944c5ee04b3856619099ab2828a5c6e2798d61233aa69fc8e371a3d2174f694ca0e720f7e0509816f117b8ffe2632784a1ac843c018d3c0df580aa10399ccc;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h69cfca4b12f95e8dac0b9f6fd827f082aa5a400de93590d17ae2a48f55513bf2f87d6c43ff1bc558a207af7f2029d6a04088159c5dea6814a98884d67ae55bc7eb8df4a369fd5f8c1eb11f232c1e33a0fb10525c2d45bae63b6ab54e0d619a18b6886b48ffa75b889a470c343713224a69c8bbeda055adce624a04ad40f79f23cdb8df70a9610b395ea7c4e6fc7a483aa408f5c70c9631d983b961bf740bc76c5804babf676e04eaf5d8e40021d66d414b097ef5384c0e9d3a0cfa29b41b01d9561355e360c09993f4c843ebcf0dd9c62a511163489b3f7a8057b65a500a8df61daa23b0ce42136346fd5889400a2ce0fcb6d06c160a59c65fd53c35ee1257efd4db5e22a3be1772c59f46b2f0d5490d52f55a068c9ecf96f2f66c16464bf57ea273be4e18ea76fdf856a3f5a78d56b3a5466edb8d80d7d9487dd88333a126941ed493852a46eb1bb676bec1eca976cf17ac8909c2d25b7d860f88da623eed30ee6d59a6f4c4754e0cd86bcd050c1b86ef5782dceda6a95afc6555b3414a0333;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hdd350e54e2b179fa0b0f61d73a7c161a0cb0339d32b4351959188705e9c8cda0071f3416322c1ea38610722a6f8b25210b89d7a429a250cd476e6ede49263817a80e653f68ae53b99748030a3c6167f5a45c6f9ee5d64293069fa1696ad0cddb7959ca0c4c3434940a578654a719b2ecbcaab8dfa64d8f22dff5d9d95efd2fa5e9a3a74466d822df6953b41e11d6fcafbb7c00258ba5cf3baa62664d63738075bc23fa4dbfba6ddf0172c700c9f3882c8d01a60a976a6e11f88ca93e0536c881943abba0e73b4638d4b8927def3fb1ff738ec239aea4512d4e03a9e668f1b592a925f85d542602f2af6fdfc21f634906f3ac3ff0453be4b28d59b5ca432757834e3f22a795277ff0b137552640b86b02002c5358e640098b91f2a67ab770a04bce69f5e17873820a823e5c75c188f60b7045c4f16798a7bb2ee6c0ac40a828c3d0f6c024e3b3b9a5dc84d50a68cf78ae79ff9de34afb108c7061585243a6ffca6903afe9ba5a4576918f1c44dc64c98d9ecd9395351088e40b6f343a42ea7e15;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h78d9372659c9adb509f7d2c3d75957a3b7b62aaa1b7e9c9bf5899cd1835d62850b3358c5aaba57e5f8916ff1b2862fc564d9355f54579375df1c1449b0a54b0c6be4e4da08f684ad3fde034434437d3299bdf5d8bdc4092b43693ce211b43c9fea420b0426a27484159124d7e8341faf7523619644b4e3b73f35e664eaa743671852894b9349f58e6480cb30b721ce55f3d1fa199e91d3b45d4c573bdde25063cf74391b40cf31eef2bd00db3d76777f7e2ab14ee722a8aa6e37393bcde18ed449f86699a44dab9e6c2b5065776a3fa56abc0bedb135b8c47b35c8f297efaea365226329bcd2666a5aa765fddc89dc8c7266e7f65c995f4387017ac02f0b7ad581df4926906e65c899ca6c198bcefce20e521804856f441ce62ce7943587cda4b0c17fdd8e95460c56691327c6dce59f5207c519b313c4aa4b89c7dd75896d7deb209182a16f0f6a7a93b1547b2ffed03857a8777286334c3150b8303650cf6e41dd43346768abdf4fc3531d4667dab114506a04461489f48029963caef7726c;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd08458fd7769f94ddac0e329d4fafbf3e2dd170fb7116664b7c309a36dc6c73b9f3d2f668517c7eef0a2cad842f339d63cb0fd10a42a59ee2cd504d846b8e1759c2bd2028630f317a494f4a47afd12d7f685f0bed33a5623a6a8648f321c38c48c1658d83d7643382d47187de272447f3e50f9ccc32b55d6f1eb992a0609b6d12df5365358089fd3135122fd8a94bfc1a6c16c5ad8282baa1310bcacbaccd9d73873a9d732fd2468507204cb14836d2bf8dd2d063717fa15cc4de04c2d321c71576ef69f66d416f0d21af42abf6c10e194a856ea5974befe6096578d8dcf3d4640dbe16f3039bc9c960fd2847e32a5dde4f0ad34f465e1669ce0809b9d5f709dd9a107948e0a7334d33498b6e7968bb9702913f1431d8badf3924918306e2f155485f1b287fdf4c2202cb1bc6803eb72da18472705e3f4af7be8f121e847d7cb91c16d608f86af4a4516475b1ecc9880f9738210b12022c43a01779d61d6719f1399e6f2258ea778a1553993412a5e0e69f93a859ec6ca56968534736fe128c0;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h6487106c75132cb302762a28183952c6ebdebbc2fda88485f2f24e4153ba78ff16bde609c202fed4f2d858c58c2bd623fe53b2b436423edc2955dce78857baf8b0baf99ef538a86d9cab42f309a1a32eccbaf5103a8436d04eac6bd668bdb0da8b681fd1b7f69adcf8517465f7a34ea7b6e55911218ec6a9d7f447e1a98f9ccf79b8943659335eda88bd7203d4e52f90749c120ea96721c5fd6e2ee3901629a4286b0a1e98d4ac141099b1494e6d66cd7e3daf31047eb3ccaab045e2e2290154377fb2577c8f0500f38553f956cfb50b2481d95449d0f0694bdeee9abf5f06f86da498397d6e0b26694ce7443c9b83b30bc7ab0d2fac4d93f6e6c1fa1baceec892bc85eae21fc26fb1e52cd9865e16ea6fd0844abb7bdf9a4bbd3223e7f5e406c4487d224fa4f4e6f6ea61612aada572d1d856dff9d86fe55834b6f2665612c70c5132e631f1056fd4467ae7dcbf64c089263b06301fb9fdc695d0f19b3d0b0a4317ca032875c96b6d3fc822852e3ee6cece5665758228acc63c8d3e4b469ae9;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'haa043f5e681ec17dd896ab8a966682b277f2162e05fcb0e7c107d2a2c8aa16f29676fe7ee76b0e4bc8ea4df74c5749e0ed639c3dfe48b146fdf72277c07463c3b68e9501d83d4acfe2883e9ce575e495aadef089fe3a2af036a3a8222ebb0e59bb0056086ac04a0b13ea701453acf7191623e668612ea388eb9464a6bf0c1adcd80f62fd53ba30b35df509c9f98074bd6c70658e62c8216d2702371be79b2b4b08f6ddd998f4e4851080f6d07ad927c265b02618076e13114d076db5f36aa28a38161cb50f5d2b439f569dcd93dfa948e28a999b3ee6451338fc5e50f71ef07cafcf6e69c1279e2c1b195017f9a4912ad1d28238c12cba457895ab6d8c8c3966ed54809fc09eb3c435bfe3714187752337ab8d85b223c6d6d4968d4228f25111100929e8dcee0b1c8fe751ad6e0acc3d2c72f3799702d771d8e8ec756a8f35268047ca348f7a7ba6c37de8eefabacfde888bc95bcd39cc47782c89c4502473bead668ec874628bb0384cd2300a9b06c0cbaea0b34ab02c2af0c944f8f156269d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hcbcbbc1a0c6e882fd7f5798280976ecff2a97d08970031e8d15ce86a4abc0df4f3be5f48279d9ee90f0e099b7be0bb867047a164658884edfbefb767f5ddfc32218479939a72987c9f70cc1a55b6bad4013446703cb2c0f79d421ce3660992c17226e9860b26407aef512a496ce4f0df4d80425a943923c4e2fc71832166a5f20bd9572bd1549824673ce00d0be3dc286fb94efb9e646b3f21e97dee11425cffad84a85349da0b33a469072276c734475d7435afd6322a3a29e0214f4aa64807053e417646f20be994ab22d908154404bdee4a42d395eaff7de42ffe7092d14932b6159f4f2ce23eba2a74c59c81cd3ebf9c8adecfdb040730b0cbb2042170daa503f51ae45d67aa1d9d5db40a8865beab55842dcf5b13fd16df685bd251f739a5b7c63d9da196126a755f902a047e2f6e854c6f2ac3840e6dcef85c5611dc3e557c750a6c0cb12e531d5ae9476e7cee26be65c8e448517d436ce395da209412c64385d830e5e1943a1542f0534ecb2435c056afc34b5244500a4cc6f15ed99d;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hade71fc35a3b5e492fe975b600fe18cf79b1378233735b9553e764cbc4e41827b644fa665a563812d6b12027bda6483cc9fceab11c676a7bc13b3fb2df0d20033feb56414398465415d8149e84cd5134cda9e4b236f96518e4c1fc89b1397c758e732c9965a987078072115e4dd219b960525179dcecc8bcdfdedc90f692a391ede4420e6739ac879e46f58ec4b3e8c6c3c6e251baa0c4d977ec0e503b64f35ff3c5ff0e0730d860b5e6fb42d926d0d4637571936ef65789ace3594089e9113ea0ff080581b29422fe3b636a2db5939c60059770705d5d433be191e730897166148f2a534ebf775f31a2584532311bc9a33f6c9dd617fa363b1dc98d6b8c25afff6afbf5903a9e6ce997153364eda604206845ae636e808307c425c6fc481f8d519a91efef5861782588b7bf0fcc8a78992d98822c0a4acecbc55051df273764ab3798f3105c7e5f3a52d81601c5a415e40b09d3b5372ae830930ce6c49c371443723c707c365f52b7080d09d5f0947c637983938cb063dc53890224c84b2ca1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h83f62dad0fe4a7d8fe4fdc1b5e12e5b281cc52e26c78bbdb7c070be8bb7f87adfbad429609adf295bcdd35f6eb08a6b6813338363030ec4b91023f1af9010bd227988ad65a6d847d18e0888a7eeeec7d799f600f38e70a8ea53d08dac07febc47c32be886a68e6e7418b61d98c17904195849639f26d8ffe672094b91a58e8a1f51e402b481407feba2ac750ef239a21d76914c2bb9b476eb1ad5ddd35c66c817a61713609d3339b4b6a6b66b66dee35fa460c699fbae0e49a0d34c5007f6ec2578406dbccfba0030a663522b2815b1a82d899bcf51cbad4f49973091091ff45135347e5ea763894331b5603979fc88c287f647aaf23f0de0176b8071a720f19afe0fc4d003d70ae13b7daa3d724b71637c4384d3d2bcf59ac1d298caeb4585b801bf925e1d9c2f501c1f1e15b9c2dadf8620022cda486d05db8d120131c3a2abcafe33eb4dd59ec07cdffeab57da457a1b7d43560b220792b8c62b1bdeede181d9f257fa4bbae7cbde985b33b1a27db6588922d4f1f73ddd1c9ec3325ae533b;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h26016fb298a3864d0f535ff0e1d470708b4d085f6cbf33d0491939ec1084351819c0a46fb62097c2347c6ab434bd3b6c44ab1671eec8716214c5758910e6291ffc4c8c1b938c7ee5aed261cce7de9da17bfec1d9618e050b8e082092f0666154fe7131ba4965de9c6d1ae86f6d9fd4f00b49b61540ead398bc4f41220a7a3fcb101c96cb1872b1d15e85a37b666a488fe1fe9d811fee8e550001a54e100536191bd1e7ecf2a56c242ed0044c75c3193d8b6727dc8f290c770b32282dd156d83f880e481f00c0f806846efc5338eccf657c6b64a9fb0e94a8007fd46b88519bc5a4b091abcba054aa1398fce3b61bb56f6fcd0ccea8e1a249268c06526a4cf54b0e82b8756f3174a4ff7895886fe03eb0b7fef53c3d6012a549ffd259a76898ccd3d681048650d3b4b9911621d50f77ed1ef3528ff0b277071b52ec8843c89411e2ee767f713962ab224fc520ed4d091048438cf23cd6f5bdaf5f35eec0c2e9775ddb987ce29f3a09094241d58e57f53bee39942ee7b8ad3ff71e31810ef8f074;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he33c525d25bb801709afab5924022e69c7babc23ba7b3f5ff8fc631bcbfb95c1a03a118b50901ed2661c687b71e10c64379cca1721aa6019cbaae3be0c13b1d6e99440234bad05c2342519dc98535606c552aa11d6f39f5068bc8212ad2c5f769ac183d10a854703d9eefc648aee35f7076dc9ca3c73a64254a5c4634eb3dba6da1c06c3ad0cf57f2fd95f7891d627bdc5e1fd1800f93afcfa40edbf8bab6ec0e049bd9214e5c9837cb84a2033dc9e11f4d73a0d93721eea09a45032a9427860d0ea6c33840d83cf6951018a4d997c3f3b07c0ee003dab0467d9c97b05aaefea6c8796859bca61e184272dec96a1f7ed7a3b5b51e49e2f5e33d3da42f9c50213707b075ba8e1288e7179446df7a8ce7bf12f923efa287c43574628c08422a3292b35fa341803d3976d21a20dcbcb66e16579d106de8ada56080192ffd098886377d4a8d92072da38c689c318bf220cb1d413a9ec68b0e90340bc5455d50583ff47c67b43f4bdd1a96aa06746c22591996ead09135bb52857d9b126ab781437e1;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he9e8ec462ec102a3684fa75a584dc1332915a523ce67b75fda3b3d34ec0b619122d268c2cb2411f5e40d6fd109a37e45dee867880de0c5a7dbff0bd6db435691a0a6ab31d7f8c3ccc7cbddf51d616ca38cc4287ac5f7c5db7f7db080b8329712c9224ad819569e03826d3bcdb0bd352d909335cfddccbbb7e3d0a138b8468e774ee3009629b5b068d496fed61ee0b01310b82e976b232866c56709d6e342f9ba0ef6cee5cc93f1cd9c33ee3f4a2f847eec8dca2057fd545c93be07d792d4a288ce327e7360740884981dd2a1e96cbba5b0d733bd2af39f98bd3e58b7cebb673a19e2567e15803cb58ff064961fcddcc842f56c2db9b4b6406c5b7ae89e7754e9e40c1886e7efca502a8344096aebcce5b5b9c8a5425b847420b6499aa0bd80446c16b9ba00a4785a8b732efb45908882a789a71562627dba437cf06ac6c381e3c165e262c4b263bf0a6b785833783443e6b17baedd993dffce83982e08c39246cdb34e2cf92f024e04eacb1cfaf7c5a755ed1de656cc919ccecb82a4c6986e57;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3fef8387d00e46bd9e545b770cffe721dd3b0eb14d985db2ca938c64bb01340e154b6a21ff3f3a15ff0475d4f77d496585122b448bd72d89f5dbee4a110bda92f675147bcc6242ebcc79ffa9fe823f187dda948ebed251e89d49d4fac46ff539cab11841071f686e659d425ec654a9ce2686a54cbd4d062971cb3d2a2e429516083ea6bad62f773c79eab2c732aead3ea4015d052642126915a2511a51d93712b6b09ba45eb34afa65a4d07f7c0f1a55e67f2167e9d5f255358e75ca69fa5e28d8f8337afddc1bf88bc5f83c515d2c142c17a66fc7310c7d921f7c5fa7dfbb8f0d1f30ac7d51649252fd6863bb78122ca652c894a44d40448233af991ad7a0ef1dbe7a751a4760d36702dc27fcebd8190f60e257e6d72d9829d4aa31828692fd82bccaa96b2add9cfcd05b8165306b534d2463430047100fd148cc34dde6c22a833d9fb1f11c7d90db66867dc86bf9265e20aaba4bb834c5e41764ff73b8e9bd2b792b5a11a247612a3d715ab634f52484d69b39606524c571b2dd21a1a9255a;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hd22103f87c6a2c9232cd5a0013c88d99902cc31aa9986a32ff46fcd6a02cb5290ae67e88e0ef4f48d277f479bbc1ea37f9d05750996e1acaa6d4d9d538d663ce80d657f5203fc6e3bba68da823baa876e702ddd6c8fd53e0f3c1a328e17fcc29fabcbd43e64c24a7de1bccbbb4eed01386afc3f55b432358c8598be5892f2e98ff4856b66f379f822c6862e9604c8da3d8907033aaf495e81e6087ae253f6c13b694fd86c8a5dca53d85abb564e512e654b45ee91ab6b16b62e345454721aba36db80f1966b3c83a7487a66deb2a676d4ed074880f49119f4ddf9c511148b3b9a2e5312fd1e41a6a4b1fed34bcb1e404e0a3ad71fb91d25df2db1f62e3a7410bc37389b8e0bc0d0e71bf1d45533d2750e51fdec16ece47ea3ea8da0a96c2c0bd0d0320eb92b16ed39e74eacce96c557c9932dfd2399051db81a0f27df936b4510266bb4354b15c4484beb7961ed29742856e242f108a885a5bca930b94593dcb45a5049c039f7f933e00a7fff1506d52eb151dd8630a1d4eb7cb69e66085b437;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'he9b397ffa4cf3c16fbca8bda097b015e5a6ea41703ee5b9298940613656e051f56e970a43bef3d05cc1d5301bdca9f17a572e6f6b962c2d816a1b7a8ed02047388bbf05930d82594b45ff60c6378f43421f5480d25e0044456c93bf66664edd6f588a44fdb5c19fc56cca2f94f489af1e35981ffc80d752df3f95bc506b9e304931624b595828c182ea23187cd2a118dd98274adbb3ac9a84d0f008a4009549a99b14eaa87058e80e487fa36ccf3f660a090f8a2990952fc46d64390b884919a793ff79103b1a1ad7f2f418426bfdb089930a7a01db14e508a35fd82203c64e590d33464f33f1221ca4fbad4bb04d0baaa5decd86422b079444b3bec777986d82dbff7bad6f302baf93f315799ffcca60d40249c2acdf918a41cbc2d15fcfacff28b473be4d0217f6c79a979b6ce983ca0f5c7f179021ca268a532d34fdac2511e2d2b3259df454f3ba1557120edc1d2e2375bcc06b55546a56a2eede5ee778507d8dda3c95f8f7875a0c34e67c79592420662bb8158164c2acf414cf49b5cc6;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'hf4218be461af4943df9d65d32df253642944fdacaf0ef0ae2cabbfe3cfd1823fa98db00d82c7ce805a31103ceef825efb665ec629abc48c5f1dbd48dbde76975ae90cdac5d080376cd51ecd88dd855b59dfd8c7685193892cc9cd97c2fea3201233a8afb0d2ade9d2ec4c84254753928d206acd46de99e050947254eba3136657a278684289ca8dd7ede7ba733c2db10260ff1d27f595f433c8b9ff0cfd78eb34ecfbea378eeacc8365c00add2662d210ea4c45592a732ee8592d3559fb7c7c469ca9e89ae92374aead367d5bbca3da67019fb3017db9be26bd739f9fade0c8e86032336c1dfd26a61f5330c4c78b12f71524b41f5e82a73a865b6ac86ae91b441b453d25f8fbc876e14e36a7251eb572132cd79bd45ab24af007c9b1694c794f27f8c6343e59e40cd80cab867544ff0e2dc778078bca14345dca49f51f9f32a2ca5f27a1c9e3ee98c1444d94b35c517d870cce05c487f9c5dffc6b6294a4087d03c1accf76bff015b9ad67f255eb9b55485d8000bf8cf68a9301098c921a397;
        #1
        {src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3072'h3bd55933c3be9563038fbeb55e4497dd5afbdbd22a23fc1051f8f99e2f0afcef30482cc374acd8e94b5c374c7a8dcd56649eb49cc8fe3a0c506579dbf2fe7f70b41bd419b07da9c9f77c96dfe91a2f509f0203963adc42c5aac3e4b520d2281eeec6356885c75817be89357254f5325486c34dab0cadf167d0992195bbe2d162c7e4851d89ab18c437ec830b05311959372f3e1e21dd94b52516ec5019c9d918713978c5c22571a727e04f44b45a24e259f3faba93ad80e33a024381c71ea45c5d046d98f0556006d95f28714605f429ae883841d93f04596f5aeaa251463a72615f7938312bc76f58b819b5dc07423b6d52144972ac00389ebe46b62eb2e883a9a2bfe55f838a0527e31001a115dc390335c3184f572ad43fc0d63492436ad4ae78e4d82b625cecb22cde4c7a8e84f02ff26beea17ef3ae7c8eaac1d06fa65b7eb557dec6d0da163d05669a0194b0358fa434f09368e5e02e396d9ef58fe55d98fa66c627280e09449199fab1bd2010a9345bd33943363efb05c802929933c;
        #1
        $finish();
    end
endmodule
