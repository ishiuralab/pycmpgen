module compressor_without_rowadder (
      input wire [25:0] src0,
      input wire [25:0] src1,
      input wire [25:0] src2,
      input wire [25:0] src3,
      input wire [25:0] src4,
      input wire [25:0] src5,
      input wire [25:0] src6,
      input wire [25:0] src7,
      input wire [25:0] src8,
      input wire [25:0] src9,
      input wire [25:0] src10,
      input wire [25:0] src11,
      input wire [25:0] src12,
      input wire [25:0] src13,
      input wire [25:0] src14,
      input wire [25:0] src15,
      input wire [25:0] src16,
      input wire [25:0] src17,
      input wire [25:0] src18,
      input wire [25:0] src19,
      input wire [25:0] src20,
      input wire [25:0] src21,
      input wire [25:0] src22,
      input wire [25:0] src23,
      input wire [25:0] src24,
      input wire [25:0] src25,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [0:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [0:0] dst27,
      output wire [1:0] dst28,
      output wire [0:0] dst29,
      output wire [0:0] dst30);

   wire [25:0] stage0_0;
   wire [25:0] stage0_1;
   wire [25:0] stage0_2;
   wire [25:0] stage0_3;
   wire [25:0] stage0_4;
   wire [25:0] stage0_5;
   wire [25:0] stage0_6;
   wire [25:0] stage0_7;
   wire [25:0] stage0_8;
   wire [25:0] stage0_9;
   wire [25:0] stage0_10;
   wire [25:0] stage0_11;
   wire [25:0] stage0_12;
   wire [25:0] stage0_13;
   wire [25:0] stage0_14;
   wire [25:0] stage0_15;
   wire [25:0] stage0_16;
   wire [25:0] stage0_17;
   wire [25:0] stage0_18;
   wire [25:0] stage0_19;
   wire [25:0] stage0_20;
   wire [25:0] stage0_21;
   wire [25:0] stage0_22;
   wire [25:0] stage0_23;
   wire [25:0] stage0_24;
   wire [25:0] stage0_25;
   wire [8:0] stage1_0;
   wire [13:0] stage1_1;
   wire [9:0] stage1_2;
   wire [11:0] stage1_3;
   wire [11:0] stage1_4;
   wire [20:0] stage1_5;
   wire [8:0] stage1_6;
   wire [20:0] stage1_7;
   wire [12:0] stage1_8;
   wire [12:0] stage1_9;
   wire [12:0] stage1_10;
   wire [11:0] stage1_11;
   wire [11:0] stage1_12;
   wire [13:0] stage1_13;
   wire [20:0] stage1_14;
   wire [12:0] stage1_15;
   wire [18:0] stage1_16;
   wire [5:0] stage1_17;
   wire [9:0] stage1_18;
   wire [16:0] stage1_19;
   wire [9:0] stage1_20;
   wire [9:0] stage1_21;
   wire [13:0] stage1_22;
   wire [17:0] stage1_23;
   wire [8:0] stage1_24;
   wire [20:0] stage1_25;
   wire [5:0] stage1_26;
   wire [1:0] stage1_27;
   wire [3:0] stage2_0;
   wire [6:0] stage2_1;
   wire [4:0] stage2_2;
   wire [2:0] stage2_3;
   wire [4:0] stage2_4;
   wire [13:0] stage2_5;
   wire [4:0] stage2_6;
   wire [12:0] stage2_7;
   wire [5:0] stage2_8;
   wire [6:0] stage2_9;
   wire [4:0] stage2_10;
   wire [3:0] stage2_11;
   wire [6:0] stage2_12;
   wire [6:0] stage2_13;
   wire [5:0] stage2_14;
   wire [5:0] stage2_15;
   wire [12:0] stage2_16;
   wire [4:0] stage2_17;
   wire [12:0] stage2_18;
   wire [6:0] stage2_19;
   wire [3:0] stage2_20;
   wire [4:0] stage2_21;
   wire [4:0] stage2_22;
   wire [5:0] stage2_23;
   wire [6:0] stage2_24;
   wire [7:0] stage2_25;
   wire [3:0] stage2_26;
   wire [4:0] stage2_27;
   wire [1:0] stage2_28;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [1:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [7:0] stage3_5;
   wire [2:0] stage3_6;
   wire [3:0] stage3_7;
   wire [3:0] stage3_8;
   wire [3:0] stage3_9;
   wire [1:0] stage3_10;
   wire [5:0] stage3_11;
   wire [2:0] stage3_12;
   wire [2:0] stage3_13;
   wire [1:0] stage3_14;
   wire [1:0] stage3_15;
   wire [4:0] stage3_16;
   wire [3:0] stage3_17;
   wire [2:0] stage3_18;
   wire [3:0] stage3_19;
   wire [6:0] stage3_20;
   wire [1:0] stage3_21;
   wire [5:0] stage3_22;
   wire [0:0] stage3_23;
   wire [5:0] stage3_24;
   wire [2:0] stage3_25;
   wire [1:0] stage3_26;
   wire [1:0] stage3_27;
   wire [3:0] stage3_28;
   wire [0:0] stage3_29;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [0:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [1:0] stage4_20;
   wire [1:0] stage4_21;
   wire [1:0] stage4_22;
   wire [1:0] stage4_23;
   wire [1:0] stage4_24;
   wire [1:0] stage4_25;
   wire [1:0] stage4_26;
   wire [0:0] stage4_27;
   wire [1:0] stage4_28;
   wire [0:0] stage4_29;
   wire [0:0] stage4_30;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;
   assign dst22 = stage4_22;
   assign dst23 = stage4_23;
   assign dst24 = stage4_24;
   assign dst25 = stage4_25;
   assign dst26 = stage4_26;
   assign dst27 = stage4_27;
   assign dst28 = stage4_28;
   assign dst29 = stage4_29;
   assign dst30 = stage4_30;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc606_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2063_5 gpc3 (
      {stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7]},
      {stage1_5[0],stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4]}
   );
   gpc606_5 gpc5 (
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[1],stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5]}
   );
   gpc615_5 gpc6 (
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22]},
      {stage0_3[14]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[6],stage1_3[6],stage1_2[6]}
   );
   gpc425_5 gpc7 (
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage0_4[6], stage0_4[7]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3]},
      {stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[7],stage1_3[7]}
   );
   gpc623_5 gpc8 (
      {stage0_3[20], stage0_3[21], stage0_3[22]},
      {stage0_4[8], stage0_4[9]},
      {stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9]},
      {stage1_7[1],stage1_6[2],stage1_5[4],stage1_4[8],stage1_3[8]}
   );
   gpc615_5 gpc9 (
      {stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14]},
      {stage0_5[10]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[2],stage1_6[3],stage1_5[5],stage1_4[9]}
   );
   gpc615_5 gpc10 (
      {stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_5[11]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[3],stage1_6[4],stage1_5[6],stage1_4[10]}
   );
   gpc2116_5 gpc11 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25]},
      {stage0_5[12]},
      {stage0_6[12]},
      {stage0_7[0], stage0_7[1]},
      {stage1_8[2],stage1_7[4],stage1_6[5],stage1_5[7],stage1_4[11]}
   );
   gpc606_5 gpc12 (
      {stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17], stage0_6[18]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[0],stage1_8[3],stage1_7[5],stage1_6[6]}
   );
   gpc606_5 gpc13 (
      {stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23], stage0_6[24]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[1],stage1_8[4],stage1_7[6],stage1_6[7]}
   );
   gpc606_5 gpc14 (
      {stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6], stage0_7[7]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[2],stage1_8[5],stage1_7[7]}
   );
   gpc606_5 gpc15 (
      {stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12], stage0_7[13]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[3],stage1_9[3],stage1_8[6],stage1_7[8]}
   );
   gpc615_5 gpc16 (
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16]},
      {stage0_9[12]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[2],stage1_10[4],stage1_9[4],stage1_8[7]}
   );
   gpc615_5 gpc17 (
      {stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_9[13]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[3],stage1_10[5],stage1_9[5],stage1_8[8]}
   );
   gpc606_5 gpc18 (
      {stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[4],stage1_10[6],stage1_9[6]}
   );
   gpc615_5 gpc19 (
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16]},
      {stage0_11[6]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[1],stage1_12[3],stage1_11[5],stage1_10[7]}
   );
   gpc615_5 gpc20 (
      {stage0_10[17], stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21]},
      {stage0_11[7]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[2],stage1_12[4],stage1_11[6],stage1_10[8]}
   );
   gpc606_5 gpc21 (
      {stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12], stage0_11[13]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[2],stage1_13[3],stage1_12[5],stage1_11[7]}
   );
   gpc615_5 gpc22 (
      {stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18]},
      {stage0_12[12]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[3],stage1_13[4],stage1_12[6],stage1_11[8]}
   );
   gpc615_5 gpc23 (
      {stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage0_12[13]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[4],stage1_13[5],stage1_12[7],stage1_11[9]}
   );
   gpc615_5 gpc24 (
      {stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18]},
      {stage0_13[18]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[3],stage1_14[5],stage1_13[6],stage1_12[8]}
   );
   gpc615_5 gpc25 (
      {stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_13[19]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[4],stage1_14[6],stage1_13[7],stage1_12[9]}
   );
   gpc615_5 gpc26 (
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4]},
      {stage0_16[0]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[0],stage1_17[0],stage1_16[2],stage1_15[5]}
   );
   gpc615_5 gpc27 (
      {stage0_15[5], stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9]},
      {stage0_16[1]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[1],stage1_17[1],stage1_16[3],stage1_15[6]}
   );
   gpc615_5 gpc28 (
      {stage0_15[10], stage0_15[11], stage0_15[12], stage0_15[13], stage0_15[14]},
      {stage0_16[2]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[2],stage1_17[2],stage1_16[4],stage1_15[7]}
   );
   gpc615_5 gpc29 (
      {stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18], stage0_15[19]},
      {stage0_16[3]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[3],stage1_17[3],stage1_16[5],stage1_15[8]}
   );
   gpc1163_5 gpc30 (
      {stage0_15[20], stage0_15[21], stage0_15[22]},
      {stage0_16[4], stage0_16[5], stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9]},
      {stage0_17[24]},
      {stage0_18[0]},
      {stage1_19[4],stage1_18[4],stage1_17[4],stage1_16[6],stage1_15[9]}
   );
   gpc615_5 gpc31 (
      {stage0_16[10], stage0_16[11], stage0_16[12], stage0_16[13], stage0_16[14]},
      {stage0_17[25]},
      {stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5], stage0_18[6]},
      {stage1_20[0],stage1_19[5],stage1_18[5],stage1_17[5],stage1_16[7]}
   );
   gpc615_5 gpc32 (
      {stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage0_19[0]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[0],stage1_20[1],stage1_19[6],stage1_18[6]}
   );
   gpc615_5 gpc33 (
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16]},
      {stage0_19[1]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[1],stage1_20[2],stage1_19[7],stage1_18[7]}
   );
   gpc615_5 gpc34 (
      {stage0_18[17], stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21]},
      {stage0_19[2]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[2],stage1_20[3],stage1_19[8],stage1_18[8]}
   );
   gpc615_5 gpc35 (
      {stage0_18[22], stage0_18[23], stage0_18[24], stage0_18[25], 1'b0},
      {stage0_19[3]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[3],stage1_20[4],stage1_19[9],stage1_18[9]}
   );
   gpc606_5 gpc36 (
      {stage0_19[4], stage0_19[5], stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[4],stage1_21[4],stage1_20[5],stage1_19[10]}
   );
   gpc606_5 gpc37 (
      {stage0_19[10], stage0_19[11], stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[5],stage1_21[5],stage1_20[6],stage1_19[11]}
   );
   gpc606_5 gpc38 (
      {stage0_19[16], stage0_19[17], stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[6],stage1_21[6],stage1_20[7],stage1_19[12]}
   );
   gpc606_5 gpc39 (
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[0],stage1_23[3],stage1_22[7],stage1_21[7]}
   );
   gpc606_5 gpc40 (
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[1],stage1_24[1],stage1_23[4],stage1_22[8]}
   );
   gpc606_5 gpc41 (
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[2],stage1_24[2],stage1_23[5],stage1_22[9]}
   );
   gpc606_5 gpc42 (
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[3],stage1_24[3],stage1_23[6],stage1_22[10]}
   );
   gpc606_5 gpc43 (
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[4],stage1_24[4],stage1_23[7],stage1_22[11]}
   );
   gpc606_5 gpc44 (
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[4],stage1_25[5],stage1_24[5],stage1_23[8]}
   );
   gpc606_5 gpc45 (
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[5],stage1_25[6],stage1_24[6],stage1_23[9]}
   );
   gpc1_1 gpc46 (
      {stage0_0[21]},
      {stage1_0[4]}
   );
   gpc1_1 gpc47 (
      {stage0_0[22]},
      {stage1_0[5]}
   );
   gpc1_1 gpc48 (
      {stage0_0[23]},
      {stage1_0[6]}
   );
   gpc1_1 gpc49 (
      {stage0_0[24]},
      {stage1_0[7]}
   );
   gpc1_1 gpc50 (
      {stage0_0[25]},
      {stage1_0[8]}
   );
   gpc1_1 gpc51 (
      {stage0_1[18]},
      {stage1_1[6]}
   );
   gpc1_1 gpc52 (
      {stage0_1[19]},
      {stage1_1[7]}
   );
   gpc1_1 gpc53 (
      {stage0_1[20]},
      {stage1_1[8]}
   );
   gpc1_1 gpc54 (
      {stage0_1[21]},
      {stage1_1[9]}
   );
   gpc1_1 gpc55 (
      {stage0_1[22]},
      {stage1_1[10]}
   );
   gpc1_1 gpc56 (
      {stage0_1[23]},
      {stage1_1[11]}
   );
   gpc1_1 gpc57 (
      {stage0_1[24]},
      {stage1_1[12]}
   );
   gpc1_1 gpc58 (
      {stage0_1[25]},
      {stage1_1[13]}
   );
   gpc1_1 gpc59 (
      {stage0_2[23]},
      {stage1_2[7]}
   );
   gpc1_1 gpc60 (
      {stage0_2[24]},
      {stage1_2[8]}
   );
   gpc1_1 gpc61 (
      {stage0_2[25]},
      {stage1_2[9]}
   );
   gpc1_1 gpc62 (
      {stage0_3[23]},
      {stage1_3[9]}
   );
   gpc1_1 gpc63 (
      {stage0_3[24]},
      {stage1_3[10]}
   );
   gpc1_1 gpc64 (
      {stage0_3[25]},
      {stage1_3[11]}
   );
   gpc1_1 gpc65 (
      {stage0_5[13]},
      {stage1_5[8]}
   );
   gpc1_1 gpc66 (
      {stage0_5[14]},
      {stage1_5[9]}
   );
   gpc1_1 gpc67 (
      {stage0_5[15]},
      {stage1_5[10]}
   );
   gpc1_1 gpc68 (
      {stage0_5[16]},
      {stage1_5[11]}
   );
   gpc1_1 gpc69 (
      {stage0_5[17]},
      {stage1_5[12]}
   );
   gpc1_1 gpc70 (
      {stage0_5[18]},
      {stage1_5[13]}
   );
   gpc1_1 gpc71 (
      {stage0_5[19]},
      {stage1_5[14]}
   );
   gpc1_1 gpc72 (
      {stage0_5[20]},
      {stage1_5[15]}
   );
   gpc1_1 gpc73 (
      {stage0_5[21]},
      {stage1_5[16]}
   );
   gpc1_1 gpc74 (
      {stage0_5[22]},
      {stage1_5[17]}
   );
   gpc1_1 gpc75 (
      {stage0_5[23]},
      {stage1_5[18]}
   );
   gpc1_1 gpc76 (
      {stage0_5[24]},
      {stage1_5[19]}
   );
   gpc1_1 gpc77 (
      {stage0_5[25]},
      {stage1_5[20]}
   );
   gpc1_1 gpc78 (
      {stage0_6[25]},
      {stage1_6[8]}
   );
   gpc1_1 gpc79 (
      {stage0_7[14]},
      {stage1_7[9]}
   );
   gpc1_1 gpc80 (
      {stage0_7[15]},
      {stage1_7[10]}
   );
   gpc1_1 gpc81 (
      {stage0_7[16]},
      {stage1_7[11]}
   );
   gpc1_1 gpc82 (
      {stage0_7[17]},
      {stage1_7[12]}
   );
   gpc1_1 gpc83 (
      {stage0_7[18]},
      {stage1_7[13]}
   );
   gpc1_1 gpc84 (
      {stage0_7[19]},
      {stage1_7[14]}
   );
   gpc1_1 gpc85 (
      {stage0_7[20]},
      {stage1_7[15]}
   );
   gpc1_1 gpc86 (
      {stage0_7[21]},
      {stage1_7[16]}
   );
   gpc1_1 gpc87 (
      {stage0_7[22]},
      {stage1_7[17]}
   );
   gpc1_1 gpc88 (
      {stage0_7[23]},
      {stage1_7[18]}
   );
   gpc1_1 gpc89 (
      {stage0_7[24]},
      {stage1_7[19]}
   );
   gpc1_1 gpc90 (
      {stage0_7[25]},
      {stage1_7[20]}
   );
   gpc1_1 gpc91 (
      {stage0_8[22]},
      {stage1_8[9]}
   );
   gpc1_1 gpc92 (
      {stage0_8[23]},
      {stage1_8[10]}
   );
   gpc1_1 gpc93 (
      {stage0_8[24]},
      {stage1_8[11]}
   );
   gpc1_1 gpc94 (
      {stage0_8[25]},
      {stage1_8[12]}
   );
   gpc1_1 gpc95 (
      {stage0_9[20]},
      {stage1_9[7]}
   );
   gpc1_1 gpc96 (
      {stage0_9[21]},
      {stage1_9[8]}
   );
   gpc1_1 gpc97 (
      {stage0_9[22]},
      {stage1_9[9]}
   );
   gpc1_1 gpc98 (
      {stage0_9[23]},
      {stage1_9[10]}
   );
   gpc1_1 gpc99 (
      {stage0_9[24]},
      {stage1_9[11]}
   );
   gpc1_1 gpc100 (
      {stage0_9[25]},
      {stage1_9[12]}
   );
   gpc1_1 gpc101 (
      {stage0_10[22]},
      {stage1_10[9]}
   );
   gpc1_1 gpc102 (
      {stage0_10[23]},
      {stage1_10[10]}
   );
   gpc1_1 gpc103 (
      {stage0_10[24]},
      {stage1_10[11]}
   );
   gpc1_1 gpc104 (
      {stage0_10[25]},
      {stage1_10[12]}
   );
   gpc1_1 gpc105 (
      {stage0_11[24]},
      {stage1_11[10]}
   );
   gpc1_1 gpc106 (
      {stage0_11[25]},
      {stage1_11[11]}
   );
   gpc1_1 gpc107 (
      {stage0_12[24]},
      {stage1_12[10]}
   );
   gpc1_1 gpc108 (
      {stage0_12[25]},
      {stage1_12[11]}
   );
   gpc1_1 gpc109 (
      {stage0_13[20]},
      {stage1_13[8]}
   );
   gpc1_1 gpc110 (
      {stage0_13[21]},
      {stage1_13[9]}
   );
   gpc1_1 gpc111 (
      {stage0_13[22]},
      {stage1_13[10]}
   );
   gpc1_1 gpc112 (
      {stage0_13[23]},
      {stage1_13[11]}
   );
   gpc1_1 gpc113 (
      {stage0_13[24]},
      {stage1_13[12]}
   );
   gpc1_1 gpc114 (
      {stage0_13[25]},
      {stage1_13[13]}
   );
   gpc1_1 gpc115 (
      {stage0_14[12]},
      {stage1_14[7]}
   );
   gpc1_1 gpc116 (
      {stage0_14[13]},
      {stage1_14[8]}
   );
   gpc1_1 gpc117 (
      {stage0_14[14]},
      {stage1_14[9]}
   );
   gpc1_1 gpc118 (
      {stage0_14[15]},
      {stage1_14[10]}
   );
   gpc1_1 gpc119 (
      {stage0_14[16]},
      {stage1_14[11]}
   );
   gpc1_1 gpc120 (
      {stage0_14[17]},
      {stage1_14[12]}
   );
   gpc1_1 gpc121 (
      {stage0_14[18]},
      {stage1_14[13]}
   );
   gpc1_1 gpc122 (
      {stage0_14[19]},
      {stage1_14[14]}
   );
   gpc1_1 gpc123 (
      {stage0_14[20]},
      {stage1_14[15]}
   );
   gpc1_1 gpc124 (
      {stage0_14[21]},
      {stage1_14[16]}
   );
   gpc1_1 gpc125 (
      {stage0_14[22]},
      {stage1_14[17]}
   );
   gpc1_1 gpc126 (
      {stage0_14[23]},
      {stage1_14[18]}
   );
   gpc1_1 gpc127 (
      {stage0_14[24]},
      {stage1_14[19]}
   );
   gpc1_1 gpc128 (
      {stage0_14[25]},
      {stage1_14[20]}
   );
   gpc1_1 gpc129 (
      {stage0_15[23]},
      {stage1_15[10]}
   );
   gpc1_1 gpc130 (
      {stage0_15[24]},
      {stage1_15[11]}
   );
   gpc1_1 gpc131 (
      {stage0_15[25]},
      {stage1_15[12]}
   );
   gpc1_1 gpc132 (
      {stage0_16[15]},
      {stage1_16[8]}
   );
   gpc1_1 gpc133 (
      {stage0_16[16]},
      {stage1_16[9]}
   );
   gpc1_1 gpc134 (
      {stage0_16[17]},
      {stage1_16[10]}
   );
   gpc1_1 gpc135 (
      {stage0_16[18]},
      {stage1_16[11]}
   );
   gpc1_1 gpc136 (
      {stage0_16[19]},
      {stage1_16[12]}
   );
   gpc1_1 gpc137 (
      {stage0_16[20]},
      {stage1_16[13]}
   );
   gpc1_1 gpc138 (
      {stage0_16[21]},
      {stage1_16[14]}
   );
   gpc1_1 gpc139 (
      {stage0_16[22]},
      {stage1_16[15]}
   );
   gpc1_1 gpc140 (
      {stage0_16[23]},
      {stage1_16[16]}
   );
   gpc1_1 gpc141 (
      {stage0_16[24]},
      {stage1_16[17]}
   );
   gpc1_1 gpc142 (
      {stage0_16[25]},
      {stage1_16[18]}
   );
   gpc1_1 gpc143 (
      {stage0_19[22]},
      {stage1_19[13]}
   );
   gpc1_1 gpc144 (
      {stage0_19[23]},
      {stage1_19[14]}
   );
   gpc1_1 gpc145 (
      {stage0_19[24]},
      {stage1_19[15]}
   );
   gpc1_1 gpc146 (
      {stage0_19[25]},
      {stage1_19[16]}
   );
   gpc1_1 gpc147 (
      {stage0_20[24]},
      {stage1_20[8]}
   );
   gpc1_1 gpc148 (
      {stage0_20[25]},
      {stage1_20[9]}
   );
   gpc1_1 gpc149 (
      {stage0_21[24]},
      {stage1_21[8]}
   );
   gpc1_1 gpc150 (
      {stage0_21[25]},
      {stage1_21[9]}
   );
   gpc1_1 gpc151 (
      {stage0_22[24]},
      {stage1_22[12]}
   );
   gpc1_1 gpc152 (
      {stage0_22[25]},
      {stage1_22[13]}
   );
   gpc1_1 gpc153 (
      {stage0_23[18]},
      {stage1_23[10]}
   );
   gpc1_1 gpc154 (
      {stage0_23[19]},
      {stage1_23[11]}
   );
   gpc1_1 gpc155 (
      {stage0_23[20]},
      {stage1_23[12]}
   );
   gpc1_1 gpc156 (
      {stage0_23[21]},
      {stage1_23[13]}
   );
   gpc1_1 gpc157 (
      {stage0_23[22]},
      {stage1_23[14]}
   );
   gpc1_1 gpc158 (
      {stage0_23[23]},
      {stage1_23[15]}
   );
   gpc1_1 gpc159 (
      {stage0_23[24]},
      {stage1_23[16]}
   );
   gpc1_1 gpc160 (
      {stage0_23[25]},
      {stage1_23[17]}
   );
   gpc1_1 gpc161 (
      {stage0_24[24]},
      {stage1_24[7]}
   );
   gpc1_1 gpc162 (
      {stage0_24[25]},
      {stage1_24[8]}
   );
   gpc1_1 gpc163 (
      {stage0_25[12]},
      {stage1_25[7]}
   );
   gpc1_1 gpc164 (
      {stage0_25[13]},
      {stage1_25[8]}
   );
   gpc1_1 gpc165 (
      {stage0_25[14]},
      {stage1_25[9]}
   );
   gpc1_1 gpc166 (
      {stage0_25[15]},
      {stage1_25[10]}
   );
   gpc1_1 gpc167 (
      {stage0_25[16]},
      {stage1_25[11]}
   );
   gpc1_1 gpc168 (
      {stage0_25[17]},
      {stage1_25[12]}
   );
   gpc1_1 gpc169 (
      {stage0_25[18]},
      {stage1_25[13]}
   );
   gpc1_1 gpc170 (
      {stage0_25[19]},
      {stage1_25[14]}
   );
   gpc1_1 gpc171 (
      {stage0_25[20]},
      {stage1_25[15]}
   );
   gpc1_1 gpc172 (
      {stage0_25[21]},
      {stage1_25[16]}
   );
   gpc1_1 gpc173 (
      {stage0_25[22]},
      {stage1_25[17]}
   );
   gpc1_1 gpc174 (
      {stage0_25[23]},
      {stage1_25[18]}
   );
   gpc1_1 gpc175 (
      {stage0_25[24]},
      {stage1_25[19]}
   );
   gpc1_1 gpc176 (
      {stage0_25[25]},
      {stage1_25[20]}
   );
   gpc606_5 gpc177 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc178 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4]},
      {stage1_2[6]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc615_5 gpc179 (
      {stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9]},
      {stage1_2[7]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc207_4 gpc180 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage1_6[0], stage1_6[1]},
      {stage2_7[0],stage2_6[0],stage2_5[2],stage2_4[3]}
   );
   gpc615_5 gpc181 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage1_5[0]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[0],stage2_7[1],stage2_6[1],stage2_5[3],stage2_4[4]}
   );
   gpc606_5 gpc182 (
      {stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5], stage1_5[6]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[2],stage2_6[2],stage2_5[4]}
   );
   gpc606_5 gpc183 (
      {stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[2],stage2_7[3],stage2_6[3],stage2_5[5]}
   );
   gpc606_5 gpc184 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[0],stage2_9[2],stage2_8[3]}
   );
   gpc606_5 gpc185 (
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[1],stage2_10[1],stage2_9[3],stage2_8[4]}
   );
   gpc606_5 gpc186 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[2],stage2_9[4]}
   );
   gpc606_5 gpc187 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[3],stage2_9[5]}
   );
   gpc606_5 gpc188 (
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[0],stage2_14[0],stage2_13[2],stage2_12[4]}
   );
   gpc615_5 gpc189 (
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10]},
      {stage1_13[0]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[1],stage2_14[1],stage2_13[3],stage2_12[5]}
   );
   gpc606_5 gpc190 (
      {stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[2],stage2_15[2],stage2_14[2],stage2_13[4]}
   );
   gpc606_5 gpc191 (
      {stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[3],stage2_15[3],stage2_14[3],stage2_13[5]}
   );
   gpc615_5 gpc192 (
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16]},
      {stage1_15[12]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[2],stage2_16[4],stage2_15[4],stage2_14[4]}
   );
   gpc615_5 gpc193 (
      {stage1_14[17], stage1_14[18], stage1_14[19], stage1_14[20], 1'b0},
      {1'b0},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[3],stage2_16[5],stage2_15[5],stage2_14[5]}
   );
   gpc606_5 gpc194 (
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[0],stage2_19[0],stage2_18[2],stage2_17[4]}
   );
   gpc606_5 gpc195 (
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[1],stage2_20[1],stage2_19[1]}
   );
   gpc606_5 gpc196 (
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[1],stage2_22[1],stage2_21[2],stage2_20[2]}
   );
   gpc606_5 gpc197 (
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], 1'b0, 1'b0},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[2],stage2_22[2],stage2_21[3],stage2_20[3]}
   );
   gpc615_5 gpc198 (
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], 1'b0},
      {stage1_22[12]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[2],stage2_23[3],stage2_22[3],stage2_21[4]}
   );
   gpc606_5 gpc199 (
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[0],stage2_25[1],stage2_24[3],stage2_23[4]}
   );
   gpc606_5 gpc200 (
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[1],stage2_25[2],stage2_24[4],stage2_23[5]}
   );
   gpc606_5 gpc201 (
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[2],stage2_26[2],stage2_25[3],stage2_24[5]}
   );
   gpc1163_5 gpc202 (
      {stage1_24[6], stage1_24[7], stage1_24[8]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {1'b0},
      {stage1_27[0]},
      {stage2_28[1],stage2_27[3],stage2_26[3],stage2_25[4],stage2_24[6]}
   );
   gpc1_1 gpc203 (
      {stage1_0[6]},
      {stage2_0[1]}
   );
   gpc1_1 gpc204 (
      {stage1_0[7]},
      {stage2_0[2]}
   );
   gpc1_1 gpc205 (
      {stage1_0[8]},
      {stage2_0[3]}
   );
   gpc1_1 gpc206 (
      {stage1_1[10]},
      {stage2_1[3]}
   );
   gpc1_1 gpc207 (
      {stage1_1[11]},
      {stage2_1[4]}
   );
   gpc1_1 gpc208 (
      {stage1_1[12]},
      {stage2_1[5]}
   );
   gpc1_1 gpc209 (
      {stage1_1[13]},
      {stage2_1[6]}
   );
   gpc1_1 gpc210 (
      {stage1_2[8]},
      {stage2_2[3]}
   );
   gpc1_1 gpc211 (
      {stage1_2[9]},
      {stage2_2[4]}
   );
   gpc1_1 gpc212 (
      {stage1_5[13]},
      {stage2_5[6]}
   );
   gpc1_1 gpc213 (
      {stage1_5[14]},
      {stage2_5[7]}
   );
   gpc1_1 gpc214 (
      {stage1_5[15]},
      {stage2_5[8]}
   );
   gpc1_1 gpc215 (
      {stage1_5[16]},
      {stage2_5[9]}
   );
   gpc1_1 gpc216 (
      {stage1_5[17]},
      {stage2_5[10]}
   );
   gpc1_1 gpc217 (
      {stage1_5[18]},
      {stage2_5[11]}
   );
   gpc1_1 gpc218 (
      {stage1_5[19]},
      {stage2_5[12]}
   );
   gpc1_1 gpc219 (
      {stage1_5[20]},
      {stage2_5[13]}
   );
   gpc1_1 gpc220 (
      {stage1_6[8]},
      {stage2_6[4]}
   );
   gpc1_1 gpc221 (
      {stage1_7[12]},
      {stage2_7[4]}
   );
   gpc1_1 gpc222 (
      {stage1_7[13]},
      {stage2_7[5]}
   );
   gpc1_1 gpc223 (
      {stage1_7[14]},
      {stage2_7[6]}
   );
   gpc1_1 gpc224 (
      {stage1_7[15]},
      {stage2_7[7]}
   );
   gpc1_1 gpc225 (
      {stage1_7[16]},
      {stage2_7[8]}
   );
   gpc1_1 gpc226 (
      {stage1_7[17]},
      {stage2_7[9]}
   );
   gpc1_1 gpc227 (
      {stage1_7[18]},
      {stage2_7[10]}
   );
   gpc1_1 gpc228 (
      {stage1_7[19]},
      {stage2_7[11]}
   );
   gpc1_1 gpc229 (
      {stage1_7[20]},
      {stage2_7[12]}
   );
   gpc1_1 gpc230 (
      {stage1_8[12]},
      {stage2_8[5]}
   );
   gpc1_1 gpc231 (
      {stage1_9[12]},
      {stage2_9[6]}
   );
   gpc1_1 gpc232 (
      {stage1_10[12]},
      {stage2_10[4]}
   );
   gpc1_1 gpc233 (
      {stage1_12[11]},
      {stage2_12[6]}
   );
   gpc1_1 gpc234 (
      {stage1_13[13]},
      {stage2_13[6]}
   );
   gpc1_1 gpc235 (
      {stage1_16[12]},
      {stage2_16[6]}
   );
   gpc1_1 gpc236 (
      {stage1_16[13]},
      {stage2_16[7]}
   );
   gpc1_1 gpc237 (
      {stage1_16[14]},
      {stage2_16[8]}
   );
   gpc1_1 gpc238 (
      {stage1_16[15]},
      {stage2_16[9]}
   );
   gpc1_1 gpc239 (
      {stage1_16[16]},
      {stage2_16[10]}
   );
   gpc1_1 gpc240 (
      {stage1_16[17]},
      {stage2_16[11]}
   );
   gpc1_1 gpc241 (
      {stage1_16[18]},
      {stage2_16[12]}
   );
   gpc1_1 gpc242 (
      {stage1_18[0]},
      {stage2_18[3]}
   );
   gpc1_1 gpc243 (
      {stage1_18[1]},
      {stage2_18[4]}
   );
   gpc1_1 gpc244 (
      {stage1_18[2]},
      {stage2_18[5]}
   );
   gpc1_1 gpc245 (
      {stage1_18[3]},
      {stage2_18[6]}
   );
   gpc1_1 gpc246 (
      {stage1_18[4]},
      {stage2_18[7]}
   );
   gpc1_1 gpc247 (
      {stage1_18[5]},
      {stage2_18[8]}
   );
   gpc1_1 gpc248 (
      {stage1_18[6]},
      {stage2_18[9]}
   );
   gpc1_1 gpc249 (
      {stage1_18[7]},
      {stage2_18[10]}
   );
   gpc1_1 gpc250 (
      {stage1_18[8]},
      {stage2_18[11]}
   );
   gpc1_1 gpc251 (
      {stage1_18[9]},
      {stage2_18[12]}
   );
   gpc1_1 gpc252 (
      {stage1_19[12]},
      {stage2_19[2]}
   );
   gpc1_1 gpc253 (
      {stage1_19[13]},
      {stage2_19[3]}
   );
   gpc1_1 gpc254 (
      {stage1_19[14]},
      {stage2_19[4]}
   );
   gpc1_1 gpc255 (
      {stage1_19[15]},
      {stage2_19[5]}
   );
   gpc1_1 gpc256 (
      {stage1_19[16]},
      {stage2_19[6]}
   );
   gpc1_1 gpc257 (
      {stage1_22[13]},
      {stage2_22[4]}
   );
   gpc1_1 gpc258 (
      {stage1_25[18]},
      {stage2_25[5]}
   );
   gpc1_1 gpc259 (
      {stage1_25[19]},
      {stage2_25[6]}
   );
   gpc1_1 gpc260 (
      {stage1_25[20]},
      {stage2_25[7]}
   );
   gpc1_1 gpc261 (
      {stage1_27[1]},
      {stage2_27[4]}
   );
   gpc2063_5 gpc262 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc263 (
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4]},
      {stage2_3[2]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], 1'b0},
      {stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1]}
   );
   gpc606_5 gpc264 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[1]}
   );
   gpc1163_5 gpc265 (
      {stage2_5[6], stage2_5[7], stage2_5[8]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], 1'b0},
      {stage2_7[6]},
      {stage2_8[0]},
      {stage3_9[1],stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[2]}
   );
   gpc615_5 gpc266 (
      {stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage2_8[1]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[2],stage3_8[2],stage3_7[2]}
   );
   gpc615_5 gpc267 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], 1'b0},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], 1'b0},
      {stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[3],stage3_8[3]}
   );
   gpc606_5 gpc268 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[1]}
   );
   gpc606_5 gpc269 (
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[1],stage3_15[1],stage3_14[1],stage3_13[1]}
   );
   gpc606_5 gpc270 (
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[0],stage3_18[0],stage3_17[1],stage3_16[2]}
   );
   gpc606_5 gpc271 (
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[1],stage3_18[1],stage3_17[2],stage3_16[3]}
   );
   gpc615_5 gpc272 (
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4]},
      {stage2_18[12]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[2],stage3_19[2],stage3_18[2],stage3_17[3]}
   );
   gpc606_5 gpc273 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], 1'b0},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[0],stage3_21[1]}
   );
   gpc623_5 gpc274 (
      {stage2_24[0], stage2_24[1], stage2_24[2]},
      {stage2_25[0], stage2_25[1]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], 1'b0, 1'b0},
      {stage3_28[0],stage3_27[0],stage3_26[0],stage3_25[1],stage3_24[1]}
   );
   gpc606_5 gpc275 (
      {stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6], stage2_25[7]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], 1'b0},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[1],stage3_25[2]}
   );
   gpc1_1 gpc276 (
      {stage2_0[3]},
      {stage3_0[1]}
   );
   gpc1_1 gpc277 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc278 (
      {stage2_5[9]},
      {stage3_5[3]}
   );
   gpc1_1 gpc279 (
      {stage2_5[10]},
      {stage3_5[4]}
   );
   gpc1_1 gpc280 (
      {stage2_5[11]},
      {stage3_5[5]}
   );
   gpc1_1 gpc281 (
      {stage2_5[12]},
      {stage3_5[6]}
   );
   gpc1_1 gpc282 (
      {stage2_5[13]},
      {stage3_5[7]}
   );
   gpc1_1 gpc283 (
      {stage2_7[12]},
      {stage3_7[3]}
   );
   gpc1_1 gpc284 (
      {stage2_11[0]},
      {stage3_11[2]}
   );
   gpc1_1 gpc285 (
      {stage2_11[1]},
      {stage3_11[3]}
   );
   gpc1_1 gpc286 (
      {stage2_11[2]},
      {stage3_11[4]}
   );
   gpc1_1 gpc287 (
      {stage2_11[3]},
      {stage3_11[5]}
   );
   gpc1_1 gpc288 (
      {stage2_12[6]},
      {stage3_12[2]}
   );
   gpc1_1 gpc289 (
      {stage2_13[6]},
      {stage3_13[2]}
   );
   gpc1_1 gpc290 (
      {stage2_16[12]},
      {stage3_16[4]}
   );
   gpc1_1 gpc291 (
      {stage2_19[6]},
      {stage3_19[3]}
   );
   gpc1_1 gpc292 (
      {stage2_20[0]},
      {stage3_20[3]}
   );
   gpc1_1 gpc293 (
      {stage2_20[1]},
      {stage3_20[4]}
   );
   gpc1_1 gpc294 (
      {stage2_20[2]},
      {stage3_20[5]}
   );
   gpc1_1 gpc295 (
      {stage2_20[3]},
      {stage3_20[6]}
   );
   gpc1_1 gpc296 (
      {stage2_22[0]},
      {stage3_22[1]}
   );
   gpc1_1 gpc297 (
      {stage2_22[1]},
      {stage3_22[2]}
   );
   gpc1_1 gpc298 (
      {stage2_22[2]},
      {stage3_22[3]}
   );
   gpc1_1 gpc299 (
      {stage2_22[3]},
      {stage3_22[4]}
   );
   gpc1_1 gpc300 (
      {stage2_22[4]},
      {stage3_22[5]}
   );
   gpc1_1 gpc301 (
      {stage2_24[3]},
      {stage3_24[2]}
   );
   gpc1_1 gpc302 (
      {stage2_24[4]},
      {stage3_24[3]}
   );
   gpc1_1 gpc303 (
      {stage2_24[5]},
      {stage3_24[4]}
   );
   gpc1_1 gpc304 (
      {stage2_24[6]},
      {stage3_24[5]}
   );
   gpc1_1 gpc305 (
      {stage2_28[0]},
      {stage3_28[2]}
   );
   gpc1_1 gpc306 (
      {stage2_28[1]},
      {stage3_28[3]}
   );
   gpc711_5 gpc307 (
      {stage3_3[0]},
      {stage3_4[0]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5], stage3_5[6]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0]}
   );
   gpc1343_5 gpc308 (
      {stage3_6[0], stage3_6[1], stage3_6[2]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3]},
      {stage3_8[0], stage3_8[1], stage3_8[2]},
      {stage3_9[0]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[1],stage4_6[1]}
   );
   gpc223_4 gpc309 (
      {stage3_9[1], stage3_9[2], stage3_9[3]},
      {stage3_10[0], stage3_10[1]},
      {stage3_11[0], stage3_11[1]},
      {stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc1334_5 gpc310 (
      {stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0], stage3_12[1], stage3_12[2]},
      {stage3_13[0], stage3_13[1], stage3_13[2]},
      {stage3_14[0]},
      {stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[1],stage4_11[1]}
   );
   gpc1343_5 gpc311 (
      {stage3_15[0], stage3_15[1], 1'b0},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3]},
      {stage3_17[0], stage3_17[1], stage3_17[2]},
      {stage3_18[0]},
      {stage4_19[0],stage4_18[0],stage4_17[0],stage4_16[0],stage4_15[1]}
   );
   gpc2143_5 gpc312 (
      {stage3_18[1], stage3_18[2], 1'b0},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3]},
      {stage3_20[0]},
      {stage3_21[0], stage3_21[1]},
      {stage4_22[0],stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[1]}
   );
   gpc606_5 gpc313 (
      {stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5], stage3_20[6]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[0],stage4_22[1],stage4_21[1],stage4_20[1]}
   );
   gpc2126_5 gpc314 (
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage3_25[0], stage3_25[1]},
      {stage3_26[0]},
      {stage3_27[0], stage3_27[1]},
      {stage4_28[0],stage4_27[0],stage4_26[0],stage4_25[0],stage4_24[1]}
   );
   gpc425_5 gpc315 (
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], 1'b0},
      {stage3_29[0], 1'b0},
      {1'b0, 1'b0, 1'b0, 1'b0},
      {stage4_30[0],stage4_29[0],stage4_28[1]}
   );
   gpc1_1 gpc316 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc317 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc318 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc319 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc320 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc321 (
      {stage3_2[1]},
      {stage4_2[1]}
   );
   gpc1_1 gpc322 (
      {stage3_3[1]},
      {stage4_3[1]}
   );
   gpc1_1 gpc323 (
      {stage3_4[1]},
      {stage4_4[1]}
   );
   gpc1_1 gpc324 (
      {stage3_5[7]},
      {stage4_5[1]}
   );
   gpc1_1 gpc325 (
      {stage3_8[3]},
      {stage4_8[1]}
   );
   gpc1_1 gpc326 (
      {stage3_14[1]},
      {stage4_14[1]}
   );
   gpc1_1 gpc327 (
      {stage3_16[4]},
      {stage4_16[1]}
   );
   gpc1_1 gpc328 (
      {stage3_17[3]},
      {stage4_17[1]}
   );
   gpc1_1 gpc329 (
      {stage3_23[0]},
      {stage4_23[1]}
   );
   gpc1_1 gpc330 (
      {stage3_25[2]},
      {stage4_25[1]}
   );
   gpc1_1 gpc331 (
      {stage3_26[1]},
      {stage4_26[1]}
   );
endmodule
module cascade_fa_31(input [1:0] src0, input [1:0] src1, input [1:0] src2, input [1:0] src3, input [1:0] src4, input [1:0] src5, input [1:0] src6, input [1:0] src7, input [1:0] src8, input [1:0] src9, input [1:0] src10, input [1:0] src11, input [1:0] src12, input [1:0] src13, input [1:0] src14, input [1:0] src15, input [1:0] src16, input [1:0] src17, input [1:0] src18, input [1:0] src19, input [1:0] src20, input [1:0] src21, input [1:0] src22, input [1:0] src23, input [1:0] src24, input [1:0] src25, input [1:0] src26, input [1:0] src27, input [1:0] src28, input [1:0] src29, input [1:0] src30, output [31:0] dst);
    wire [30:0] gene;
    wire [30:0] prop;
    wire [31:0] out;
    wire [31:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene0(
        .O(gene[0]),
        .I0(src0[0]),
        .I1(src0[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop0(
        .O(prop[0]),
        .I0(src0[0]),
        .I1(src0[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene1(
        .O(gene[1]),
        .I0(src1[0]),
        .I1(src1[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop1(
        .O(prop[1]),
        .I0(src1[0]),
        .I1(src1[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene2(
        .O(gene[2]),
        .I0(src2[0]),
        .I1(src2[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop2(
        .O(prop[2]),
        .I0(src2[0]),
        .I1(src2[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene3(
        .O(gene[3]),
        .I0(src3[0]),
        .I1(src3[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop3(
        .O(prop[3]),
        .I0(src3[0]),
        .I1(src3[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene4(
        .O(gene[4]),
        .I0(src4[0]),
        .I1(src4[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop4(
        .O(prop[4]),
        .I0(src4[0]),
        .I1(src4[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene5(
        .O(gene[5]),
        .I0(src5[0]),
        .I1(src5[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop5(
        .O(prop[5]),
        .I0(src5[0]),
        .I1(src5[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene6(
        .O(gene[6]),
        .I0(src6[0]),
        .I1(src6[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop6(
        .O(prop[6]),
        .I0(src6[0]),
        .I1(src6[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene7(
        .O(gene[7]),
        .I0(src7[0]),
        .I1(src7[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop7(
        .O(prop[7]),
        .I0(src7[0]),
        .I1(src7[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene8(
        .O(gene[8]),
        .I0(src8[0]),
        .I1(src8[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop8(
        .O(prop[8]),
        .I0(src8[0]),
        .I1(src8[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene9(
        .O(gene[9]),
        .I0(src9[0]),
        .I1(src9[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop9(
        .O(prop[9]),
        .I0(src9[0]),
        .I1(src9[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene10(
        .O(gene[10]),
        .I0(src10[0]),
        .I1(src10[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop10(
        .O(prop[10]),
        .I0(src10[0]),
        .I1(src10[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene11(
        .O(gene[11]),
        .I0(src11[0]),
        .I1(src11[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop11(
        .O(prop[11]),
        .I0(src11[0]),
        .I1(src11[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene12(
        .O(gene[12]),
        .I0(src12[0]),
        .I1(src12[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop12(
        .O(prop[12]),
        .I0(src12[0]),
        .I1(src12[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene13(
        .O(gene[13]),
        .I0(src13[0]),
        .I1(src13[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop13(
        .O(prop[13]),
        .I0(src13[0]),
        .I1(src13[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene14(
        .O(gene[14]),
        .I0(src14[0]),
        .I1(src14[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop14(
        .O(prop[14]),
        .I0(src14[0]),
        .I1(src14[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene15(
        .O(gene[15]),
        .I0(src15[0]),
        .I1(src15[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop15(
        .O(prop[15]),
        .I0(src15[0]),
        .I1(src15[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene16(
        .O(gene[16]),
        .I0(src16[0]),
        .I1(src16[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop16(
        .O(prop[16]),
        .I0(src16[0]),
        .I1(src16[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene17(
        .O(gene[17]),
        .I0(src17[0]),
        .I1(src17[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop17(
        .O(prop[17]),
        .I0(src17[0]),
        .I1(src17[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene18(
        .O(gene[18]),
        .I0(src18[0]),
        .I1(src18[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop18(
        .O(prop[18]),
        .I0(src18[0]),
        .I1(src18[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene19(
        .O(gene[19]),
        .I0(src19[0]),
        .I1(src19[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop19(
        .O(prop[19]),
        .I0(src19[0]),
        .I1(src19[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene20(
        .O(gene[20]),
        .I0(src20[0]),
        .I1(src20[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop20(
        .O(prop[20]),
        .I0(src20[0]),
        .I1(src20[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene21(
        .O(gene[21]),
        .I0(src21[0]),
        .I1(src21[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop21(
        .O(prop[21]),
        .I0(src21[0]),
        .I1(src21[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene22(
        .O(gene[22]),
        .I0(src22[0]),
        .I1(src22[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop22(
        .O(prop[22]),
        .I0(src22[0]),
        .I1(src22[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene23(
        .O(gene[23]),
        .I0(src23[0]),
        .I1(src23[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop23(
        .O(prop[23]),
        .I0(src23[0]),
        .I1(src23[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene24(
        .O(gene[24]),
        .I0(src24[0]),
        .I1(src24[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop24(
        .O(prop[24]),
        .I0(src24[0]),
        .I1(src24[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene25(
        .O(gene[25]),
        .I0(src25[0]),
        .I1(src25[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop25(
        .O(prop[25]),
        .I0(src25[0]),
        .I1(src25[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene26(
        .O(gene[26]),
        .I0(src26[0]),
        .I1(src26[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop26(
        .O(prop[26]),
        .I0(src26[0]),
        .I1(src26[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene27(
        .O(gene[27]),
        .I0(src27[0]),
        .I1(src27[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop27(
        .O(prop[27]),
        .I0(src27[0]),
        .I1(src27[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene28(
        .O(gene[28]),
        .I0(src28[0]),
        .I1(src28[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop28(
        .O(prop[28]),
        .I0(src28[0]),
        .I1(src28[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene29(
        .O(gene[29]),
        .I0(src29[0]),
        .I1(src29[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop29(
        .O(prop[29]),
        .I0(src29[0]),
        .I1(src29[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut2_gene30(
        .O(gene[30]),
        .I0(src30[0]),
        .I1(src30[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut2_prop30(
        .O(prop[30]),
        .I0(src30[0]),
        .I1(src30[1])
    );
    CARRY4 carry4_inst0(
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CYINIT(1'h0),
        .CI(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_inst1(
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CYINIT(1'h0),
        .CI(carryout[3]),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_inst2(
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CYINIT(1'h0),
        .CI(carryout[7]),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_inst3(
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CYINIT(1'h0),
        .CI(carryout[11]),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_inst4(
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CYINIT(1'h0),
        .CI(carryout[15]),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    CARRY4 carry4_inst5(
        .CO(carryout[23:20]),
        .O(out[23:20]),
        .CYINIT(1'h0),
        .CI(carryout[19]),
        .DI(gene[23:20]),
        .S(prop[23:20])
    );
    CARRY4 carry4_inst6(
        .CO(carryout[27:24]),
        .O(out[27:24]),
        .CYINIT(1'h0),
        .CI(carryout[23]),
        .DI(gene[27:24]),
        .S(prop[27:24])
    );
    CARRY4 carry4_inst7(
        .CO(carryout[31:28]),
        .O(out[31:28]),
        .CYINIT(1'h0),
        .CI(carryout[27]),
        .DI({1'h0, gene[30:28]}),
        .S({1'h0, prop[30:28]})
    );
    assign dst = {carryout[30], out[30], out[29], out[28], out[27], out[26], out[25], out[24], out[23], out[22], out[21], out[20], out[19], out[18], out[17], out[16], out[15], out[14], out[13], out[12], out[11], out[10], out[9], out[8], out[7], out[6], out[5], out[4], out[3], out[2], out[1], out[0]};
endmodule

module rowadder2_1_31_(input [30:0] src0, input [30:0] src1, output [31:0] dst0);
    cascade_fa_31 cascade_fa_31(.src0({src0[0], src1[0]}), .src1({src0[1], src1[1]}), .src2({src0[2], src1[2]}), .src3({src0[3], src1[3]}), .src4({src0[4], src1[4]}), .src5({src0[5], src1[5]}), .src6({src0[6], src1[6]}), .src7({src0[7], src1[7]}), .src8({src0[8], src1[8]}), .src9({src0[9], src1[9]}), .src10({src0[10], src1[10]}), .src11({src0[11], src1[11]}), .src12({src0[12], src1[12]}), .src13({src0[13], src1[13]}), .src14({src0[14], src1[14]}), .src15({src0[15], src1[15]}), .src16({src0[16], src1[16]}), .src17({src0[17], src1[17]}), .src18({src0[18], src1[18]}), .src19({src0[19], src1[19]}), .src20({src0[20], src1[20]}), .src21({src0[21], src1[21]}), .src22({src0[22], src1[22]}), .src23({src0[23], src1[23]}), .src24({src0[24], src1[24]}), .src25({src0[25], src1[25]}), .src26({src0[26], src1[26]}), .src27({src0[27], src1[27]}), .src28({src0[28], src1[28]}), .src29({src0[29], src1[29]}), .src30({src0[30], src1[30]}), .dst(dst0));
endmodule


module rowadder(input [1:0] src0, input [1:0] src1, input [1:0] src2, input [1:0] src3, input [1:0] src4, input [1:0] src5, input [1:0] src6, input [1:0] src7, input [1:0] src8, input [1:0] src9, input [1:0] src10, input [1:0] src11, input [1:0] src12, input [1:0] src13, input [1:0] src14, input [1:0] src15, input [1:0] src16, input [1:0] src17, input [1:0] src18, input [1:0] src19, input [1:0] src20, input [1:0] src21, input [1:0] src22, input [1:0] src23, input [1:0] src24, input [1:0] src25, input [1:0] src26, input [1:0] src27, input [1:0] src28, input [1:0] src29, input [1:0] src30, output dst0, output dst1, output dst2, output dst3, output dst4, output dst5, output dst6, output dst7, output dst8, output dst9, output dst10, output dst11, output dst12, output dst13, output dst14, output dst15, output dst16, output dst17, output dst18, output dst19, output dst20, output dst21, output dst22, output dst23, output dst24, output dst25, output dst26, output dst27, output dst28, output dst29, output dst30, output dst31);
    rowadder_rowwise ra(.src0({src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}), .src1({src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}), .dst0({dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0}));
endmodule
module rowadder_rowwise(input [30:0] src0, input [30:0] src1, output [31:0] dst0);
    wire [31:0] internal0;
    assign dst0 = internal0;
    rowadder2_1_31_ rowadder_0(.src0(src0), .src1(src1), .dst0(internal0));
endmodule

module compressor(input [25:0] src0, input [25:0] src1, input [25:0] src2, input [25:0] src3, input [25:0] src4, input [25:0] src5, input [25:0] src6, input [25:0] src7, input [25:0] src8, input [25:0] src9, input [25:0] src10, input [25:0] src11, input [25:0] src12, input [25:0] src13, input [25:0] src14, input [25:0] src15, input [25:0] src16, input [25:0] src17, input [25:0] src18, input [25:0] src19, input [25:0] src20, input [25:0] src21, input [25:0] src22, input [25:0] src23, input [25:0] src24, input [25:0] src25, output dst0, output dst1, output dst2, output dst3, output dst4, output dst5, output dst6, output dst7, output dst8, output dst9, output dst10, output dst11, output dst12, output dst13, output dst14, output dst15, output dst16, output dst17, output dst18, output dst19, output dst20, output dst21, output dst22, output dst23, output dst24, output dst25, output dst26, output dst27, output dst28, output dst29, output dst30, output dst31);
    wire [1:0] compdst0;
    wire [1:0] compdst1;
    wire [1:0] compdst2;
    wire [1:0] compdst3;
    wire [1:0] compdst4;
    wire [1:0] compdst5;
    wire [1:0] compdst6;
    wire [1:0] compdst7;
    wire [1:0] compdst8;
    wire [1:0] compdst9;
    wire [1:0] compdst10;
    wire [1:0] compdst11;
    wire [1:0] compdst12;
    wire [0:0] compdst13;
    wire [1:0] compdst14;
    wire [1:0] compdst15;
    wire [1:0] compdst16;
    wire [1:0] compdst17;
    wire [1:0] compdst18;
    wire [1:0] compdst19;
    wire [1:0] compdst20;
    wire [1:0] compdst21;
    wire [1:0] compdst22;
    wire [1:0] compdst23;
    wire [1:0] compdst24;
    wire [1:0] compdst25;
    wire [1:0] compdst26;
    wire [0:0] compdst27;
    wire [1:0] compdst28;
    wire [0:0] compdst29;
    wire [0:0] compdst30;
    compressor_without_rowadder comp(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .dst0(compdst0), .dst1(compdst1), .dst2(compdst2), .dst3(compdst3), .dst4(compdst4), .dst5(compdst5), .dst6(compdst6), .dst7(compdst7), .dst8(compdst8), .dst9(compdst9), .dst10(compdst10), .dst11(compdst11), .dst12(compdst12), .dst13(compdst13), .dst14(compdst14), .dst15(compdst15), .dst16(compdst16), .dst17(compdst17), .dst18(compdst18), .dst19(compdst19), .dst20(compdst20), .dst21(compdst21), .dst22(compdst22), .dst23(compdst23), .dst24(compdst24), .dst25(compdst25), .dst26(compdst26), .dst27(compdst27), .dst28(compdst28), .dst29(compdst29), .dst30(compdst30));
    rowadder ra(.src0(compdst0), .src1(compdst1), .src2(compdst2), .src3(compdst3), .src4(compdst4), .src5(compdst5), .src6(compdst6), .src7(compdst7), .src8(compdst8), .src9(compdst9), .src10(compdst10), .src11(compdst11), .src12(compdst12), .src13({1'h0, compdst13}), .src14(compdst14), .src15(compdst15), .src16(compdst16), .src17(compdst17), .src18(compdst18), .src19(compdst19), .src20(compdst20), .src21(compdst21), .src22(compdst22), .src23(compdst23), .src24(compdst24), .src25(compdst25), .src26(compdst26), .src27({1'h0, compdst27}), .src28(compdst28), .src29({1'h0, compdst29}), .src30({1'h0, compdst30}), .dst0(dst0), .dst1(dst1), .dst2(dst2), .dst3(dst3), .dst4(dst4), .dst5(dst5), .dst6(dst6), .dst7(dst7), .dst8(dst8), .dst9(dst9), .dst10(dst10), .dst11(dst11), .dst12(dst12), .dst13(dst13), .dst14(dst14), .dst15(dst15), .dst16(dst16), .dst17(dst17), .dst18(dst18), .dst19(dst19), .dst20(dst20), .dst21(dst21), .dst22(dst22), .dst23(dst23), .dst24(dst24), .dst25(dst25), .dst26(dst26), .dst27(dst27), .dst28(dst28), .dst29(dst29), .dst30(dst30), .dst31(dst31));
endmodule

