module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70,
        output wire [0:0] dst71);
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    reg [255:0] src32;
    reg [255:0] src33;
    reg [255:0] src34;
    reg [255:0] src35;
    reg [255:0] src36;
    reg [255:0] src37;
    reg [255:0] src38;
    reg [255:0] src39;
    reg [255:0] src40;
    reg [255:0] src41;
    reg [255:0] src42;
    reg [255:0] src43;
    reg [255:0] src44;
    reg [255:0] src45;
    reg [255:0] src46;
    reg [255:0] src47;
    reg [255:0] src48;
    reg [255:0] src49;
    reg [255:0] src50;
    reg [255:0] src51;
    reg [255:0] src52;
    reg [255:0] src53;
    reg [255:0] src54;
    reg [255:0] src55;
    reg [255:0] src56;
    reg [255:0] src57;
    reg [255:0] src58;
    reg [255:0] src59;
    reg [255:0] src60;
    reg [255:0] src61;
    reg [255:0] src62;
    reg [255:0] src63;
    compressor_CLA256_64 compressor_CLA256_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70),
            .dst71(dst71));
    initial begin
        src0 <= 256'h0;
        src1 <= 256'h0;
        src2 <= 256'h0;
        src3 <= 256'h0;
        src4 <= 256'h0;
        src5 <= 256'h0;
        src6 <= 256'h0;
        src7 <= 256'h0;
        src8 <= 256'h0;
        src9 <= 256'h0;
        src10 <= 256'h0;
        src11 <= 256'h0;
        src12 <= 256'h0;
        src13 <= 256'h0;
        src14 <= 256'h0;
        src15 <= 256'h0;
        src16 <= 256'h0;
        src17 <= 256'h0;
        src18 <= 256'h0;
        src19 <= 256'h0;
        src20 <= 256'h0;
        src21 <= 256'h0;
        src22 <= 256'h0;
        src23 <= 256'h0;
        src24 <= 256'h0;
        src25 <= 256'h0;
        src26 <= 256'h0;
        src27 <= 256'h0;
        src28 <= 256'h0;
        src29 <= 256'h0;
        src30 <= 256'h0;
        src31 <= 256'h0;
        src32 <= 256'h0;
        src33 <= 256'h0;
        src34 <= 256'h0;
        src35 <= 256'h0;
        src36 <= 256'h0;
        src37 <= 256'h0;
        src38 <= 256'h0;
        src39 <= 256'h0;
        src40 <= 256'h0;
        src41 <= 256'h0;
        src42 <= 256'h0;
        src43 <= 256'h0;
        src44 <= 256'h0;
        src45 <= 256'h0;
        src46 <= 256'h0;
        src47 <= 256'h0;
        src48 <= 256'h0;
        src49 <= 256'h0;
        src50 <= 256'h0;
        src51 <= 256'h0;
        src52 <= 256'h0;
        src53 <= 256'h0;
        src54 <= 256'h0;
        src55 <= 256'h0;
        src56 <= 256'h0;
        src57 <= 256'h0;
        src58 <= 256'h0;
        src59 <= 256'h0;
        src60 <= 256'h0;
        src61 <= 256'h0;
        src62 <= 256'h0;
        src63 <= 256'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA256_64(
    input [255:0]src0,
    input [255:0]src1,
    input [255:0]src2,
    input [255:0]src3,
    input [255:0]src4,
    input [255:0]src5,
    input [255:0]src6,
    input [255:0]src7,
    input [255:0]src8,
    input [255:0]src9,
    input [255:0]src10,
    input [255:0]src11,
    input [255:0]src12,
    input [255:0]src13,
    input [255:0]src14,
    input [255:0]src15,
    input [255:0]src16,
    input [255:0]src17,
    input [255:0]src18,
    input [255:0]src19,
    input [255:0]src20,
    input [255:0]src21,
    input [255:0]src22,
    input [255:0]src23,
    input [255:0]src24,
    input [255:0]src25,
    input [255:0]src26,
    input [255:0]src27,
    input [255:0]src28,
    input [255:0]src29,
    input [255:0]src30,
    input [255:0]src31,
    input [255:0]src32,
    input [255:0]src33,
    input [255:0]src34,
    input [255:0]src35,
    input [255:0]src36,
    input [255:0]src37,
    input [255:0]src38,
    input [255:0]src39,
    input [255:0]src40,
    input [255:0]src41,
    input [255:0]src42,
    input [255:0]src43,
    input [255:0]src44,
    input [255:0]src45,
    input [255:0]src46,
    input [255:0]src47,
    input [255:0]src48,
    input [255:0]src49,
    input [255:0]src50,
    input [255:0]src51,
    input [255:0]src52,
    input [255:0]src53,
    input [255:0]src54,
    input [255:0]src55,
    input [255:0]src56,
    input [255:0]src57,
    input [255:0]src58,
    input [255:0]src59,
    input [255:0]src60,
    input [255:0]src61,
    input [255:0]src62,
    input [255:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70,
    output dst71);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [0:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [0:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [0:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [0:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [1:0] comp_out69;
    wire [1:0] comp_out70;
    wire [0:0] comp_out71;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70),
        .dst71(comp_out71)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out71[0], comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out70[1], comp_out69[1], comp_out68[1], comp_out67[1], comp_out66[1], 1'h0, comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], 1'h0, comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], 1'h0, comp_out33[1], comp_out32[1], 1'h0, comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], 1'h0}),
        .dst({dst71, dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [255:0] src0,
      input wire [255:0] src1,
      input wire [255:0] src2,
      input wire [255:0] src3,
      input wire [255:0] src4,
      input wire [255:0] src5,
      input wire [255:0] src6,
      input wire [255:0] src7,
      input wire [255:0] src8,
      input wire [255:0] src9,
      input wire [255:0] src10,
      input wire [255:0] src11,
      input wire [255:0] src12,
      input wire [255:0] src13,
      input wire [255:0] src14,
      input wire [255:0] src15,
      input wire [255:0] src16,
      input wire [255:0] src17,
      input wire [255:0] src18,
      input wire [255:0] src19,
      input wire [255:0] src20,
      input wire [255:0] src21,
      input wire [255:0] src22,
      input wire [255:0] src23,
      input wire [255:0] src24,
      input wire [255:0] src25,
      input wire [255:0] src26,
      input wire [255:0] src27,
      input wire [255:0] src28,
      input wire [255:0] src29,
      input wire [255:0] src30,
      input wire [255:0] src31,
      input wire [255:0] src32,
      input wire [255:0] src33,
      input wire [255:0] src34,
      input wire [255:0] src35,
      input wire [255:0] src36,
      input wire [255:0] src37,
      input wire [255:0] src38,
      input wire [255:0] src39,
      input wire [255:0] src40,
      input wire [255:0] src41,
      input wire [255:0] src42,
      input wire [255:0] src43,
      input wire [255:0] src44,
      input wire [255:0] src45,
      input wire [255:0] src46,
      input wire [255:0] src47,
      input wire [255:0] src48,
      input wire [255:0] src49,
      input wire [255:0] src50,
      input wire [255:0] src51,
      input wire [255:0] src52,
      input wire [255:0] src53,
      input wire [255:0] src54,
      input wire [255:0] src55,
      input wire [255:0] src56,
      input wire [255:0] src57,
      input wire [255:0] src58,
      input wire [255:0] src59,
      input wire [255:0] src60,
      input wire [255:0] src61,
      input wire [255:0] src62,
      input wire [255:0] src63,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [0:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [0:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [0:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [0:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [1:0] dst69,
      output wire [1:0] dst70,
      output wire [0:0] dst71);

   wire [255:0] stage0_0;
   wire [255:0] stage0_1;
   wire [255:0] stage0_2;
   wire [255:0] stage0_3;
   wire [255:0] stage0_4;
   wire [255:0] stage0_5;
   wire [255:0] stage0_6;
   wire [255:0] stage0_7;
   wire [255:0] stage0_8;
   wire [255:0] stage0_9;
   wire [255:0] stage0_10;
   wire [255:0] stage0_11;
   wire [255:0] stage0_12;
   wire [255:0] stage0_13;
   wire [255:0] stage0_14;
   wire [255:0] stage0_15;
   wire [255:0] stage0_16;
   wire [255:0] stage0_17;
   wire [255:0] stage0_18;
   wire [255:0] stage0_19;
   wire [255:0] stage0_20;
   wire [255:0] stage0_21;
   wire [255:0] stage0_22;
   wire [255:0] stage0_23;
   wire [255:0] stage0_24;
   wire [255:0] stage0_25;
   wire [255:0] stage0_26;
   wire [255:0] stage0_27;
   wire [255:0] stage0_28;
   wire [255:0] stage0_29;
   wire [255:0] stage0_30;
   wire [255:0] stage0_31;
   wire [255:0] stage0_32;
   wire [255:0] stage0_33;
   wire [255:0] stage0_34;
   wire [255:0] stage0_35;
   wire [255:0] stage0_36;
   wire [255:0] stage0_37;
   wire [255:0] stage0_38;
   wire [255:0] stage0_39;
   wire [255:0] stage0_40;
   wire [255:0] stage0_41;
   wire [255:0] stage0_42;
   wire [255:0] stage0_43;
   wire [255:0] stage0_44;
   wire [255:0] stage0_45;
   wire [255:0] stage0_46;
   wire [255:0] stage0_47;
   wire [255:0] stage0_48;
   wire [255:0] stage0_49;
   wire [255:0] stage0_50;
   wire [255:0] stage0_51;
   wire [255:0] stage0_52;
   wire [255:0] stage0_53;
   wire [255:0] stage0_54;
   wire [255:0] stage0_55;
   wire [255:0] stage0_56;
   wire [255:0] stage0_57;
   wire [255:0] stage0_58;
   wire [255:0] stage0_59;
   wire [255:0] stage0_60;
   wire [255:0] stage0_61;
   wire [255:0] stage0_62;
   wire [255:0] stage0_63;
   wire [90:0] stage1_0;
   wire [82:0] stage1_1;
   wire [130:0] stage1_2;
   wire [106:0] stage1_3;
   wire [121:0] stage1_4;
   wire [95:0] stage1_5;
   wire [115:0] stage1_6;
   wire [109:0] stage1_7;
   wire [131:0] stage1_8;
   wire [119:0] stage1_9;
   wire [155:0] stage1_10;
   wire [153:0] stage1_11;
   wire [132:0] stage1_12;
   wire [96:0] stage1_13;
   wire [84:0] stage1_14;
   wire [131:0] stage1_15;
   wire [119:0] stage1_16;
   wire [110:0] stage1_17;
   wire [99:0] stage1_18;
   wire [125:0] stage1_19;
   wire [129:0] stage1_20;
   wire [107:0] stage1_21;
   wire [91:0] stage1_22;
   wire [128:0] stage1_23;
   wire [139:0] stage1_24;
   wire [109:0] stage1_25;
   wire [140:0] stage1_26;
   wire [118:0] stage1_27;
   wire [126:0] stage1_28;
   wire [109:0] stage1_29;
   wire [90:0] stage1_30;
   wire [114:0] stage1_31;
   wire [114:0] stage1_32;
   wire [110:0] stage1_33;
   wire [103:0] stage1_34;
   wire [118:0] stage1_35;
   wire [144:0] stage1_36;
   wire [104:0] stage1_37;
   wire [136:0] stage1_38;
   wire [124:0] stage1_39;
   wire [91:0] stage1_40;
   wire [142:0] stage1_41;
   wire [171:0] stage1_42;
   wire [78:0] stage1_43;
   wire [145:0] stage1_44;
   wire [158:0] stage1_45;
   wire [100:0] stage1_46;
   wire [129:0] stage1_47;
   wire [107:0] stage1_48;
   wire [151:0] stage1_49;
   wire [98:0] stage1_50;
   wire [105:0] stage1_51;
   wire [139:0] stage1_52;
   wire [107:0] stage1_53;
   wire [159:0] stage1_54;
   wire [89:0] stage1_55;
   wire [177:0] stage1_56;
   wire [104:0] stage1_57;
   wire [85:0] stage1_58;
   wire [147:0] stage1_59;
   wire [141:0] stage1_60;
   wire [108:0] stage1_61;
   wire [200:0] stage1_62;
   wire [68:0] stage1_63;
   wire [63:0] stage1_64;
   wire [41:0] stage1_65;
   wire [29:0] stage2_0;
   wire [36:0] stage2_1;
   wire [36:0] stage2_2;
   wire [53:0] stage2_3;
   wire [44:0] stage2_4;
   wire [45:0] stage2_5;
   wire [51:0] stage2_6;
   wire [42:0] stage2_7;
   wire [42:0] stage2_8;
   wire [59:0] stage2_9;
   wire [69:0] stage2_10;
   wire [48:0] stage2_11;
   wire [53:0] stage2_12;
   wire [63:0] stage2_13;
   wire [44:0] stage2_14;
   wire [73:0] stage2_15;
   wire [54:0] stage2_16;
   wire [56:0] stage2_17;
   wire [65:0] stage2_18;
   wire [36:0] stage2_19;
   wire [79:0] stage2_20;
   wire [48:0] stage2_21;
   wire [40:0] stage2_22;
   wire [60:0] stage2_23;
   wire [81:0] stage2_24;
   wire [50:0] stage2_25;
   wire [51:0] stage2_26;
   wire [71:0] stage2_27;
   wire [72:0] stage2_28;
   wire [45:0] stage2_29;
   wire [58:0] stage2_30;
   wire [53:0] stage2_31;
   wire [46:0] stage2_32;
   wire [51:0] stage2_33;
   wire [36:0] stage2_34;
   wire [58:0] stage2_35;
   wire [62:0] stage2_36;
   wire [54:0] stage2_37;
   wire [46:0] stage2_38;
   wire [80:0] stage2_39;
   wire [44:0] stage2_40;
   wire [74:0] stage2_41;
   wire [62:0] stage2_42;
   wire [61:0] stage2_43;
   wire [51:0] stage2_44;
   wire [78:0] stage2_45;
   wire [62:0] stage2_46;
   wire [70:0] stage2_47;
   wire [41:0] stage2_48;
   wire [114:0] stage2_49;
   wire [67:0] stage2_50;
   wire [78:0] stage2_51;
   wire [50:0] stage2_52;
   wire [77:0] stage2_53;
   wire [74:0] stage2_54;
   wire [34:0] stage2_55;
   wire [72:0] stage2_56;
   wire [82:0] stage2_57;
   wire [47:0] stage2_58;
   wire [47:0] stage2_59;
   wire [62:0] stage2_60;
   wire [56:0] stage2_61;
   wire [52:0] stage2_62;
   wire [74:0] stage2_63;
   wire [44:0] stage2_64;
   wire [17:0] stage2_65;
   wire [16:0] stage2_66;
   wire [6:0] stage2_67;
   wire [13:0] stage3_0;
   wire [10:0] stage3_1;
   wire [17:0] stage3_2;
   wire [18:0] stage3_3;
   wire [20:0] stage3_4;
   wire [34:0] stage3_5;
   wire [16:0] stage3_6;
   wire [27:0] stage3_7;
   wire [17:0] stage3_8;
   wire [15:0] stage3_9;
   wire [32:0] stage3_10;
   wire [30:0] stage3_11;
   wire [24:0] stage3_12;
   wire [23:0] stage3_13;
   wire [26:0] stage3_14;
   wire [40:0] stage3_15;
   wire [19:0] stage3_16;
   wire [29:0] stage3_17;
   wire [27:0] stage3_18;
   wire [27:0] stage3_19;
   wire [23:0] stage3_20;
   wire [23:0] stage3_21;
   wire [28:0] stage3_22;
   wire [15:0] stage3_23;
   wire [30:0] stage3_24;
   wire [33:0] stage3_25;
   wire [23:0] stage3_26;
   wire [21:0] stage3_27;
   wire [28:0] stage3_28;
   wire [34:0] stage3_29;
   wire [25:0] stage3_30;
   wire [31:0] stage3_31;
   wire [27:0] stage3_32;
   wire [26:0] stage3_33;
   wire [26:0] stage3_34;
   wire [32:0] stage3_35;
   wire [19:0] stage3_36;
   wire [18:0] stage3_37;
   wire [22:0] stage3_38;
   wire [30:0] stage3_39;
   wire [29:0] stage3_40;
   wire [23:0] stage3_41;
   wire [29:0] stage3_42;
   wire [38:0] stage3_43;
   wire [21:0] stage3_44;
   wire [38:0] stage3_45;
   wire [39:0] stage3_46;
   wire [32:0] stage3_47;
   wire [23:0] stage3_48;
   wire [67:0] stage3_49;
   wire [29:0] stage3_50;
   wire [47:0] stage3_51;
   wire [39:0] stage3_52;
   wire [27:0] stage3_53;
   wire [27:0] stage3_54;
   wire [29:0] stage3_55;
   wire [25:0] stage3_56;
   wire [32:0] stage3_57;
   wire [28:0] stage3_58;
   wire [32:0] stage3_59;
   wire [34:0] stage3_60;
   wire [23:0] stage3_61;
   wire [27:0] stage3_62;
   wire [27:0] stage3_63;
   wire [17:0] stage3_64;
   wire [27:0] stage3_65;
   wire [27:0] stage3_66;
   wire [1:0] stage3_67;
   wire [0:0] stage3_68;
   wire [0:0] stage3_69;
   wire [13:0] stage4_0;
   wire [4:0] stage4_1;
   wire [6:0] stage4_2;
   wire [18:0] stage4_3;
   wire [9:0] stage4_4;
   wire [19:0] stage4_5;
   wire [9:0] stage4_6;
   wire [9:0] stage4_7;
   wire [21:0] stage4_8;
   wire [7:0] stage4_9;
   wire [13:0] stage4_10;
   wire [11:0] stage4_11;
   wire [17:0] stage4_12;
   wire [13:0] stage4_13;
   wire [11:0] stage4_14;
   wire [11:0] stage4_15;
   wire [12:0] stage4_16;
   wire [14:0] stage4_17;
   wire [10:0] stage4_18;
   wire [13:0] stage4_19;
   wire [10:0] stage4_20;
   wire [8:0] stage4_21;
   wire [14:0] stage4_22;
   wire [8:0] stage4_23;
   wire [11:0] stage4_24;
   wire [13:0] stage4_25;
   wire [12:0] stage4_26;
   wire [6:0] stage4_27;
   wire [11:0] stage4_28;
   wire [16:0] stage4_29;
   wire [11:0] stage4_30;
   wire [9:0] stage4_31;
   wire [17:0] stage4_32;
   wire [16:0] stage4_33;
   wire [10:0] stage4_34;
   wire [16:0] stage4_35;
   wire [12:0] stage4_36;
   wire [11:0] stage4_37;
   wire [6:0] stage4_38;
   wire [8:0] stage4_39;
   wire [12:0] stage4_40;
   wire [11:0] stage4_41;
   wire [14:0] stage4_42;
   wire [19:0] stage4_43;
   wire [13:0] stage4_44;
   wire [11:0] stage4_45;
   wire [14:0] stage4_46;
   wire [14:0] stage4_47;
   wire [14:0] stage4_48;
   wire [35:0] stage4_49;
   wire [16:0] stage4_50;
   wire [19:0] stage4_51;
   wire [13:0] stage4_52;
   wire [14:0] stage4_53;
   wire [17:0] stage4_54;
   wire [12:0] stage4_55;
   wire [11:0] stage4_56;
   wire [11:0] stage4_57;
   wire [19:0] stage4_58;
   wire [11:0] stage4_59;
   wire [13:0] stage4_60;
   wire [11:0] stage4_61;
   wire [11:0] stage4_62;
   wire [12:0] stage4_63;
   wire [11:0] stage4_64;
   wire [7:0] stage4_65;
   wire [23:0] stage4_66;
   wire [8:0] stage4_67;
   wire [2:0] stage4_68;
   wire [0:0] stage4_69;
   wire [4:0] stage5_0;
   wire [3:0] stage5_1;
   wire [1:0] stage5_2;
   wire [6:0] stage5_3;
   wire [9:0] stage5_4;
   wire [7:0] stage5_5;
   wire [5:0] stage5_6;
   wire [6:0] stage5_7;
   wire [4:0] stage5_8;
   wire [9:0] stage5_9;
   wire [5:0] stage5_10;
   wire [9:0] stage5_11;
   wire [5:0] stage5_12;
   wire [5:0] stage5_13;
   wire [4:0] stage5_14;
   wire [5:0] stage5_15;
   wire [5:0] stage5_16;
   wire [7:0] stage5_17;
   wire [5:0] stage5_18;
   wire [10:0] stage5_19;
   wire [2:0] stage5_20;
   wire [11:0] stage5_21;
   wire [4:0] stage5_22;
   wire [2:0] stage5_23;
   wire [6:0] stage5_24;
   wire [5:0] stage5_25;
   wire [5:0] stage5_26;
   wire [5:0] stage5_27;
   wire [3:0] stage5_28;
   wire [7:0] stage5_29;
   wire [5:0] stage5_30;
   wire [6:0] stage5_31;
   wire [3:0] stage5_32;
   wire [6:0] stage5_33;
   wire [6:0] stage5_34;
   wire [4:0] stage5_35;
   wire [6:0] stage5_36;
   wire [11:0] stage5_37;
   wire [3:0] stage5_38;
   wire [2:0] stage5_39;
   wire [5:0] stage5_40;
   wire [4:0] stage5_41;
   wire [6:0] stage5_42;
   wire [9:0] stage5_43;
   wire [6:0] stage5_44;
   wire [4:0] stage5_45;
   wire [6:0] stage5_46;
   wire [6:0] stage5_47;
   wire [6:0] stage5_48;
   wire [7:0] stage5_49;
   wire [8:0] stage5_50;
   wire [9:0] stage5_51;
   wire [7:0] stage5_52;
   wire [14:0] stage5_53;
   wire [5:0] stage5_54;
   wire [5:0] stage5_55;
   wire [5:0] stage5_56;
   wire [6:0] stage5_57;
   wire [4:0] stage5_58;
   wire [6:0] stage5_59;
   wire [8:0] stage5_60;
   wire [3:0] stage5_61;
   wire [3:0] stage5_62;
   wire [5:0] stage5_63;
   wire [5:0] stage5_64;
   wire [4:0] stage5_65;
   wire [10:0] stage5_66;
   wire [6:0] stage5_67;
   wire [4:0] stage5_68;
   wire [2:0] stage5_69;
   wire [4:0] stage6_0;
   wire [3:0] stage6_1;
   wire [0:0] stage6_2;
   wire [1:0] stage6_3;
   wire [4:0] stage6_4;
   wire [3:0] stage6_5;
   wire [1:0] stage6_6;
   wire [2:0] stage6_7;
   wire [2:0] stage6_8;
   wire [8:0] stage6_9;
   wire [1:0] stage6_10;
   wire [5:0] stage6_11;
   wire [2:0] stage6_12;
   wire [1:0] stage6_13;
   wire [6:0] stage6_14;
   wire [2:0] stage6_15;
   wire [1:0] stage6_16;
   wire [2:0] stage6_17;
   wire [3:0] stage6_18;
   wire [3:0] stage6_19;
   wire [3:0] stage6_20;
   wire [1:0] stage6_21;
   wire [2:0] stage6_22;
   wire [4:0] stage6_23;
   wire [1:0] stage6_24;
   wire [6:0] stage6_25;
   wire [1:0] stage6_26;
   wire [2:0] stage6_27;
   wire [1:0] stage6_28;
   wire [2:0] stage6_29;
   wire [2:0] stage6_30;
   wire [2:0] stage6_31;
   wire [2:0] stage6_32;
   wire [3:0] stage6_33;
   wire [2:0] stage6_34;
   wire [3:0] stage6_35;
   wire [3:0] stage6_36;
   wire [7:0] stage6_37;
   wire [1:0] stage6_38;
   wire [2:0] stage6_39;
   wire [1:0] stage6_40;
   wire [1:0] stage6_41;
   wire [2:0] stage6_42;
   wire [5:0] stage6_43;
   wire [2:0] stage6_44;
   wire [3:0] stage6_45;
   wire [1:0] stage6_46;
   wire [5:0] stage6_47;
   wire [3:0] stage6_48;
   wire [2:0] stage6_49;
   wire [3:0] stage6_50;
   wire [4:0] stage6_51;
   wire [2:0] stage6_52;
   wire [3:0] stage6_53;
   wire [3:0] stage6_54;
   wire [3:0] stage6_55;
   wire [5:0] stage6_56;
   wire [2:0] stage6_57;
   wire [1:0] stage6_58;
   wire [5:0] stage6_59;
   wire [4:0] stage6_60;
   wire [4:0] stage6_61;
   wire [4:0] stage6_62;
   wire [0:0] stage6_63;
   wire [1:0] stage6_64;
   wire [1:0] stage6_65;
   wire [2:0] stage6_66;
   wire [4:0] stage6_67;
   wire [2:0] stage6_68;
   wire [1:0] stage6_69;
   wire [1:0] stage6_70;
   wire [0:0] stage6_71;
   wire [0:0] stage7_0;
   wire [1:0] stage7_1;
   wire [0:0] stage7_2;
   wire [1:0] stage7_3;
   wire [1:0] stage7_4;
   wire [1:0] stage7_5;
   wire [1:0] stage7_6;
   wire [1:0] stage7_7;
   wire [1:0] stage7_8;
   wire [1:0] stage7_9;
   wire [1:0] stage7_10;
   wire [1:0] stage7_11;
   wire [1:0] stage7_12;
   wire [1:0] stage7_13;
   wire [1:0] stage7_14;
   wire [1:0] stage7_15;
   wire [1:0] stage7_16;
   wire [1:0] stage7_17;
   wire [1:0] stage7_18;
   wire [1:0] stage7_19;
   wire [1:0] stage7_20;
   wire [1:0] stage7_21;
   wire [1:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage7_24;
   wire [1:0] stage7_25;
   wire [1:0] stage7_26;
   wire [1:0] stage7_27;
   wire [1:0] stage7_28;
   wire [1:0] stage7_29;
   wire [1:0] stage7_30;
   wire [0:0] stage7_31;
   wire [1:0] stage7_32;
   wire [1:0] stage7_33;
   wire [0:0] stage7_34;
   wire [1:0] stage7_35;
   wire [1:0] stage7_36;
   wire [1:0] stage7_37;
   wire [1:0] stage7_38;
   wire [1:0] stage7_39;
   wire [1:0] stage7_40;
   wire [1:0] stage7_41;
   wire [1:0] stage7_42;
   wire [1:0] stage7_43;
   wire [1:0] stage7_44;
   wire [1:0] stage7_45;
   wire [1:0] stage7_46;
   wire [0:0] stage7_47;
   wire [1:0] stage7_48;
   wire [1:0] stage7_49;
   wire [1:0] stage7_50;
   wire [1:0] stage7_51;
   wire [1:0] stage7_52;
   wire [1:0] stage7_53;
   wire [1:0] stage7_54;
   wire [1:0] stage7_55;
   wire [1:0] stage7_56;
   wire [1:0] stage7_57;
   wire [1:0] stage7_58;
   wire [1:0] stage7_59;
   wire [1:0] stage7_60;
   wire [1:0] stage7_61;
   wire [1:0] stage7_62;
   wire [1:0] stage7_63;
   wire [1:0] stage7_64;
   wire [0:0] stage7_65;
   wire [1:0] stage7_66;
   wire [1:0] stage7_67;
   wire [1:0] stage7_68;
   wire [1:0] stage7_69;
   wire [1:0] stage7_70;
   wire [0:0] stage7_71;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage7_0;
   assign dst1 = stage7_1;
   assign dst2 = stage7_2;
   assign dst3 = stage7_3;
   assign dst4 = stage7_4;
   assign dst5 = stage7_5;
   assign dst6 = stage7_6;
   assign dst7 = stage7_7;
   assign dst8 = stage7_8;
   assign dst9 = stage7_9;
   assign dst10 = stage7_10;
   assign dst11 = stage7_11;
   assign dst12 = stage7_12;
   assign dst13 = stage7_13;
   assign dst14 = stage7_14;
   assign dst15 = stage7_15;
   assign dst16 = stage7_16;
   assign dst17 = stage7_17;
   assign dst18 = stage7_18;
   assign dst19 = stage7_19;
   assign dst20 = stage7_20;
   assign dst21 = stage7_21;
   assign dst22 = stage7_22;
   assign dst23 = stage7_23;
   assign dst24 = stage7_24;
   assign dst25 = stage7_25;
   assign dst26 = stage7_26;
   assign dst27 = stage7_27;
   assign dst28 = stage7_28;
   assign dst29 = stage7_29;
   assign dst30 = stage7_30;
   assign dst31 = stage7_31;
   assign dst32 = stage7_32;
   assign dst33 = stage7_33;
   assign dst34 = stage7_34;
   assign dst35 = stage7_35;
   assign dst36 = stage7_36;
   assign dst37 = stage7_37;
   assign dst38 = stage7_38;
   assign dst39 = stage7_39;
   assign dst40 = stage7_40;
   assign dst41 = stage7_41;
   assign dst42 = stage7_42;
   assign dst43 = stage7_43;
   assign dst44 = stage7_44;
   assign dst45 = stage7_45;
   assign dst46 = stage7_46;
   assign dst47 = stage7_47;
   assign dst48 = stage7_48;
   assign dst49 = stage7_49;
   assign dst50 = stage7_50;
   assign dst51 = stage7_51;
   assign dst52 = stage7_52;
   assign dst53 = stage7_53;
   assign dst54 = stage7_54;
   assign dst55 = stage7_55;
   assign dst56 = stage7_56;
   assign dst57 = stage7_57;
   assign dst58 = stage7_58;
   assign dst59 = stage7_59;
   assign dst60 = stage7_60;
   assign dst61 = stage7_61;
   assign dst62 = stage7_62;
   assign dst63 = stage7_63;
   assign dst64 = stage7_64;
   assign dst65 = stage7_65;
   assign dst66 = stage7_66;
   assign dst67 = stage7_67;
   assign dst68 = stage7_68;
   assign dst69 = stage7_69;
   assign dst70 = stage7_70;
   assign dst71 = stage7_71;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc2135_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44]},
      {stage0_1[24], stage0_1[25], stage0_1[26]},
      {stage0_2[8]},
      {stage0_3[16], stage0_3[17]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc2135_5 gpc9 (
      {stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[9]},
      {stage0_3[18], stage0_3[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[10]},
      {stage0_3[20]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[11]},
      {stage0_3[21]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[12]},
      {stage0_3[22]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[13]},
      {stage0_3[23]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[14]},
      {stage0_3[24]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_2[15]},
      {stage0_3[25]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[68], stage0_0[69], stage0_0[70]},
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_2[16]},
      {stage0_3[26]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[71], stage0_0[72], stage0_0[73]},
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_2[17]},
      {stage0_3[27]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_2[18]},
      {stage0_3[28]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_2[19]},
      {stage0_3[29]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[80], stage0_0[81], stage0_0[82]},
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_2[20]},
      {stage0_3[30]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[83], stage0_0[84], stage0_0[85]},
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_2[21]},
      {stage0_3[31]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[86], stage0_0[87], stage0_0[88]},
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_2[22]},
      {stage0_3[32]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_2[23]},
      {stage0_3[33]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[92], stage0_0[93], stage0_0[94]},
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_2[24]},
      {stage0_3[34]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_2[25]},
      {stage0_3[35]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_2[26]},
      {stage0_3[36]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_2[27]},
      {stage0_3[37]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[104], stage0_0[105], stage0_0[106]},
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_2[28]},
      {stage0_3[38]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_2[29]},
      {stage0_3[39]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_2[30], stage0_2[31], stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_2[36], stage0_2[37], stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41]},
      {stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc606_5 gpc32 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_2[42], stage0_2[43], stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47]},
      {stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc606_5 gpc33 (
      {stage0_0[128], stage0_0[129], stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133]},
      {stage0_2[48], stage0_2[49], stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53]},
      {stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc606_5 gpc34 (
      {stage0_0[134], stage0_0[135], stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139]},
      {stage0_2[54], stage0_2[55], stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59]},
      {stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc606_5 gpc35 (
      {stage0_0[140], stage0_0[141], stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145]},
      {stage0_2[60], stage0_2[61], stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65]},
      {stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc606_5 gpc36 (
      {stage0_0[146], stage0_0[147], stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151]},
      {stage0_2[66], stage0_2[67], stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71]},
      {stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc606_5 gpc37 (
      {stage0_0[152], stage0_0[153], stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157]},
      {stage0_2[72], stage0_2[73], stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77]},
      {stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc606_5 gpc38 (
      {stage0_0[158], stage0_0[159], stage0_0[160], stage0_0[161], stage0_0[162], stage0_0[163]},
      {stage0_2[78], stage0_2[79], stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83]},
      {stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc606_5 gpc39 (
      {stage0_0[164], stage0_0[165], stage0_0[166], stage0_0[167], stage0_0[168], stage0_0[169]},
      {stage0_2[84], stage0_2[85], stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89]},
      {stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc606_5 gpc40 (
      {stage0_0[170], stage0_0[171], stage0_0[172], stage0_0[173], stage0_0[174], stage0_0[175]},
      {stage0_2[90], stage0_2[91], stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95]},
      {stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc606_5 gpc41 (
      {stage0_0[176], stage0_0[177], stage0_0[178], stage0_0[179], stage0_0[180], stage0_0[181]},
      {stage0_2[96], stage0_2[97], stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101]},
      {stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc606_5 gpc42 (
      {stage0_0[182], stage0_0[183], stage0_0[184], stage0_0[185], stage0_0[186], stage0_0[187]},
      {stage0_2[102], stage0_2[103], stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107]},
      {stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc606_5 gpc43 (
      {stage0_0[188], stage0_0[189], stage0_0[190], stage0_0[191], stage0_0[192], stage0_0[193]},
      {stage0_2[108], stage0_2[109], stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113]},
      {stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc606_5 gpc44 (
      {stage0_0[194], stage0_0[195], stage0_0[196], stage0_0[197], stage0_0[198], stage0_0[199]},
      {stage0_2[114], stage0_2[115], stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119]},
      {stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[200], stage0_0[201], stage0_0[202], stage0_0[203], stage0_0[204], stage0_0[205]},
      {stage0_2[120], stage0_2[121], stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125]},
      {stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[206], stage0_0[207], stage0_0[208], stage0_0[209], stage0_0[210], stage0_0[211]},
      {stage0_2[126], stage0_2[127], stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131]},
      {stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[0],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[1],stage1_4[48],stage1_3[48],stage1_2[48],stage1_1[48]}
   );
   gpc606_5 gpc49 (
      {stage0_1[162], stage0_1[163], stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[2],stage1_4[49],stage1_3[49],stage1_2[49],stage1_1[49]}
   );
   gpc606_5 gpc50 (
      {stage0_1[168], stage0_1[169], stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[3],stage1_4[50],stage1_3[50],stage1_2[50],stage1_1[50]}
   );
   gpc606_5 gpc51 (
      {stage0_1[174], stage0_1[175], stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[4],stage1_4[51],stage1_3[51],stage1_2[51],stage1_1[51]}
   );
   gpc606_5 gpc52 (
      {stage0_1[180], stage0_1[181], stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[5],stage1_4[52],stage1_3[52],stage1_2[52],stage1_1[52]}
   );
   gpc606_5 gpc53 (
      {stage0_1[186], stage0_1[187], stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[6],stage1_4[53],stage1_3[53],stage1_2[53],stage1_1[53]}
   );
   gpc606_5 gpc54 (
      {stage0_1[192], stage0_1[193], stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[7],stage1_4[54],stage1_3[54],stage1_2[54],stage1_1[54]}
   );
   gpc606_5 gpc55 (
      {stage0_1[198], stage0_1[199], stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[8],stage1_4[55],stage1_3[55],stage1_2[55],stage1_1[55]}
   );
   gpc606_5 gpc56 (
      {stage0_1[204], stage0_1[205], stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[9],stage1_4[56],stage1_3[56],stage1_2[56],stage1_1[56]}
   );
   gpc606_5 gpc57 (
      {stage0_1[210], stage0_1[211], stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[10],stage1_4[57],stage1_3[57],stage1_2[57],stage1_1[57]}
   );
   gpc606_5 gpc58 (
      {stage0_1[216], stage0_1[217], stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[11],stage1_4[58],stage1_3[58],stage1_2[58],stage1_1[58]}
   );
   gpc606_5 gpc59 (
      {stage0_1[222], stage0_1[223], stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[12],stage1_4[59],stage1_3[59],stage1_2[59],stage1_1[59]}
   );
   gpc606_5 gpc60 (
      {stage0_1[228], stage0_1[229], stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[13],stage1_4[60],stage1_3[60],stage1_2[60],stage1_1[60]}
   );
   gpc606_5 gpc61 (
      {stage0_2[132], stage0_2[133], stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[14],stage1_4[61],stage1_3[61],stage1_2[61]}
   );
   gpc606_5 gpc62 (
      {stage0_2[138], stage0_2[139], stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[15],stage1_4[62],stage1_3[62],stage1_2[62]}
   );
   gpc615_5 gpc63 (
      {stage0_2[144], stage0_2[145], stage0_2[146], stage0_2[147], stage0_2[148]},
      {stage0_3[124]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[16],stage1_4[63],stage1_3[63],stage1_2[63]}
   );
   gpc615_5 gpc64 (
      {stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152], stage0_2[153]},
      {stage0_3[125]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[17],stage1_4[64],stage1_3[64],stage1_2[64]}
   );
   gpc615_5 gpc65 (
      {stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage0_3[126]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[18],stage1_4[65],stage1_3[65],stage1_2[65]}
   );
   gpc615_5 gpc66 (
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163]},
      {stage0_3[127]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[19],stage1_4[66],stage1_3[66],stage1_2[66]}
   );
   gpc615_5 gpc67 (
      {stage0_2[164], stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168]},
      {stage0_3[128]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[20],stage1_4[67],stage1_3[67],stage1_2[67]}
   );
   gpc615_5 gpc68 (
      {stage0_2[169], stage0_2[170], stage0_2[171], stage0_2[172], stage0_2[173]},
      {stage0_3[129]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[21],stage1_4[68],stage1_3[68],stage1_2[68]}
   );
   gpc615_5 gpc69 (
      {stage0_2[174], stage0_2[175], stage0_2[176], stage0_2[177], stage0_2[178]},
      {stage0_3[130]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[22],stage1_4[69],stage1_3[69],stage1_2[69]}
   );
   gpc615_5 gpc70 (
      {stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182], stage0_2[183]},
      {stage0_3[131]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[23],stage1_4[70],stage1_3[70],stage1_2[70]}
   );
   gpc615_5 gpc71 (
      {stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage0_3[132]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[24],stage1_4[71],stage1_3[71],stage1_2[71]}
   );
   gpc615_5 gpc72 (
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193]},
      {stage0_3[133]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[25],stage1_4[72],stage1_3[72],stage1_2[72]}
   );
   gpc615_5 gpc73 (
      {stage0_2[194], stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198]},
      {stage0_3[134]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[26],stage1_4[73],stage1_3[73],stage1_2[73]}
   );
   gpc615_5 gpc74 (
      {stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138], stage0_3[139]},
      {stage0_4[78]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[13],stage1_5[27],stage1_4[74],stage1_3[74]}
   );
   gpc615_5 gpc75 (
      {stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage0_4[79]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[14],stage1_5[28],stage1_4[75],stage1_3[75]}
   );
   gpc615_5 gpc76 (
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149]},
      {stage0_4[80]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[15],stage1_5[29],stage1_4[76],stage1_3[76]}
   );
   gpc615_5 gpc77 (
      {stage0_3[150], stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154]},
      {stage0_4[81]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[16],stage1_5[30],stage1_4[77],stage1_3[77]}
   );
   gpc615_5 gpc78 (
      {stage0_3[155], stage0_3[156], stage0_3[157], stage0_3[158], stage0_3[159]},
      {stage0_4[82]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[17],stage1_5[31],stage1_4[78],stage1_3[78]}
   );
   gpc615_5 gpc79 (
      {stage0_3[160], stage0_3[161], stage0_3[162], stage0_3[163], stage0_3[164]},
      {stage0_4[83]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[18],stage1_5[32],stage1_4[79],stage1_3[79]}
   );
   gpc615_5 gpc80 (
      {stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168], stage0_3[169]},
      {stage0_4[84]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[19],stage1_5[33],stage1_4[80],stage1_3[80]}
   );
   gpc615_5 gpc81 (
      {stage0_3[170], stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174]},
      {stage0_4[85]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[20],stage1_5[34],stage1_4[81],stage1_3[81]}
   );
   gpc615_5 gpc82 (
      {stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178], stage0_3[179]},
      {stage0_4[86]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[21],stage1_5[35],stage1_4[82],stage1_3[82]}
   );
   gpc615_5 gpc83 (
      {stage0_3[180], stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184]},
      {stage0_4[87]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[22],stage1_5[36],stage1_4[83],stage1_3[83]}
   );
   gpc615_5 gpc84 (
      {stage0_3[185], stage0_3[186], stage0_3[187], stage0_3[188], stage0_3[189]},
      {stage0_4[88]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[23],stage1_5[37],stage1_4[84],stage1_3[84]}
   );
   gpc615_5 gpc85 (
      {stage0_3[190], stage0_3[191], stage0_3[192], stage0_3[193], stage0_3[194]},
      {stage0_4[89]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[24],stage1_5[38],stage1_4[85],stage1_3[85]}
   );
   gpc615_5 gpc86 (
      {stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198], stage0_3[199]},
      {stage0_4[90]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[25],stage1_5[39],stage1_4[86],stage1_3[86]}
   );
   gpc615_5 gpc87 (
      {stage0_3[200], stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204]},
      {stage0_4[91]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[26],stage1_5[40],stage1_4[87],stage1_3[87]}
   );
   gpc615_5 gpc88 (
      {stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208], stage0_3[209]},
      {stage0_4[92]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[27],stage1_5[41],stage1_4[88],stage1_3[88]}
   );
   gpc615_5 gpc89 (
      {stage0_3[210], stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214]},
      {stage0_4[93]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[28],stage1_5[42],stage1_4[89],stage1_3[89]}
   );
   gpc615_5 gpc90 (
      {stage0_3[215], stage0_3[216], stage0_3[217], stage0_3[218], stage0_3[219]},
      {stage0_4[94]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[29],stage1_5[43],stage1_4[90],stage1_3[90]}
   );
   gpc615_5 gpc91 (
      {stage0_3[220], stage0_3[221], stage0_3[222], stage0_3[223], stage0_3[224]},
      {stage0_4[95]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[30],stage1_5[44],stage1_4[91],stage1_3[91]}
   );
   gpc615_5 gpc92 (
      {stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228], stage0_3[229]},
      {stage0_4[96]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[31],stage1_5[45],stage1_4[92],stage1_3[92]}
   );
   gpc615_5 gpc93 (
      {stage0_3[230], stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234]},
      {stage0_4[97]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[32],stage1_5[46],stage1_4[93],stage1_3[93]}
   );
   gpc615_5 gpc94 (
      {stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239]},
      {stage0_4[98]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[33],stage1_5[47],stage1_4[94],stage1_3[94]}
   );
   gpc615_5 gpc95 (
      {stage0_3[240], stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244]},
      {stage0_4[99]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[34],stage1_5[48],stage1_4[95],stage1_3[95]}
   );
   gpc606_5 gpc96 (
      {stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[22],stage1_6[35],stage1_5[49],stage1_4[96]}
   );
   gpc606_5 gpc97 (
      {stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[23],stage1_6[36],stage1_5[50],stage1_4[97]}
   );
   gpc606_5 gpc98 (
      {stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[24],stage1_6[37],stage1_5[51],stage1_4[98]}
   );
   gpc606_5 gpc99 (
      {stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[25],stage1_6[38],stage1_5[52],stage1_4[99]}
   );
   gpc606_5 gpc100 (
      {stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[26],stage1_6[39],stage1_5[53],stage1_4[100]}
   );
   gpc606_5 gpc101 (
      {stage0_4[130], stage0_4[131], stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[27],stage1_6[40],stage1_5[54],stage1_4[101]}
   );
   gpc606_5 gpc102 (
      {stage0_4[136], stage0_4[137], stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[28],stage1_6[41],stage1_5[55],stage1_4[102]}
   );
   gpc606_5 gpc103 (
      {stage0_4[142], stage0_4[143], stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[29],stage1_6[42],stage1_5[56],stage1_4[103]}
   );
   gpc606_5 gpc104 (
      {stage0_4[148], stage0_4[149], stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[30],stage1_6[43],stage1_5[57],stage1_4[104]}
   );
   gpc606_5 gpc105 (
      {stage0_4[154], stage0_4[155], stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[31],stage1_6[44],stage1_5[58],stage1_4[105]}
   );
   gpc606_5 gpc106 (
      {stage0_4[160], stage0_4[161], stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[32],stage1_6[45],stage1_5[59],stage1_4[106]}
   );
   gpc606_5 gpc107 (
      {stage0_4[166], stage0_4[167], stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[33],stage1_6[46],stage1_5[60],stage1_4[107]}
   );
   gpc606_5 gpc108 (
      {stage0_4[172], stage0_4[173], stage0_4[174], stage0_4[175], stage0_4[176], stage0_4[177]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[34],stage1_6[47],stage1_5[61],stage1_4[108]}
   );
   gpc606_5 gpc109 (
      {stage0_4[178], stage0_4[179], stage0_4[180], stage0_4[181], stage0_4[182], stage0_4[183]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[35],stage1_6[48],stage1_5[62],stage1_4[109]}
   );
   gpc606_5 gpc110 (
      {stage0_4[184], stage0_4[185], stage0_4[186], stage0_4[187], stage0_4[188], stage0_4[189]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[36],stage1_6[49],stage1_5[63],stage1_4[110]}
   );
   gpc606_5 gpc111 (
      {stage0_4[190], stage0_4[191], stage0_4[192], stage0_4[193], stage0_4[194], stage0_4[195]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[37],stage1_6[50],stage1_5[64],stage1_4[111]}
   );
   gpc606_5 gpc112 (
      {stage0_4[196], stage0_4[197], stage0_4[198], stage0_4[199], stage0_4[200], stage0_4[201]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[38],stage1_6[51],stage1_5[65],stage1_4[112]}
   );
   gpc606_5 gpc113 (
      {stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206], stage0_4[207]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[39],stage1_6[52],stage1_5[66],stage1_4[113]}
   );
   gpc606_5 gpc114 (
      {stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212], stage0_4[213]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[40],stage1_6[53],stage1_5[67],stage1_4[114]}
   );
   gpc606_5 gpc115 (
      {stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218], stage0_4[219]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[41],stage1_6[54],stage1_5[68],stage1_4[115]}
   );
   gpc606_5 gpc116 (
      {stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224], stage0_4[225]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[42],stage1_6[55],stage1_5[69],stage1_4[116]}
   );
   gpc606_5 gpc117 (
      {stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230], stage0_4[231]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[43],stage1_6[56],stage1_5[70],stage1_4[117]}
   );
   gpc606_5 gpc118 (
      {stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236], stage0_4[237]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[44],stage1_6[57],stage1_5[71],stage1_4[118]}
   );
   gpc606_5 gpc119 (
      {stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242], stage0_4[243]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[45],stage1_6[58],stage1_5[72],stage1_4[119]}
   );
   gpc606_5 gpc120 (
      {stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248], stage0_4[249]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[46],stage1_6[59],stage1_5[73],stage1_4[120]}
   );
   gpc606_5 gpc121 (
      {stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254], stage0_4[255]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[47],stage1_6[60],stage1_5[74],stage1_4[121]}
   );
   gpc606_5 gpc122 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[26],stage1_7[48],stage1_6[61],stage1_5[75]}
   );
   gpc606_5 gpc123 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[27],stage1_7[49],stage1_6[62],stage1_5[76]}
   );
   gpc606_5 gpc124 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[28],stage1_7[50],stage1_6[63],stage1_5[77]}
   );
   gpc606_5 gpc125 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[29],stage1_7[51],stage1_6[64],stage1_5[78]}
   );
   gpc606_5 gpc126 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[30],stage1_7[52],stage1_6[65],stage1_5[79]}
   );
   gpc606_5 gpc127 (
      {stage0_5[162], stage0_5[163], stage0_5[164], stage0_5[165], stage0_5[166], stage0_5[167]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[31],stage1_7[53],stage1_6[66],stage1_5[80]}
   );
   gpc606_5 gpc128 (
      {stage0_5[168], stage0_5[169], stage0_5[170], stage0_5[171], stage0_5[172], stage0_5[173]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[32],stage1_7[54],stage1_6[67],stage1_5[81]}
   );
   gpc606_5 gpc129 (
      {stage0_5[174], stage0_5[175], stage0_5[176], stage0_5[177], stage0_5[178], stage0_5[179]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[33],stage1_7[55],stage1_6[68],stage1_5[82]}
   );
   gpc606_5 gpc130 (
      {stage0_5[180], stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[34],stage1_7[56],stage1_6[69],stage1_5[83]}
   );
   gpc606_5 gpc131 (
      {stage0_5[186], stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[35],stage1_7[57],stage1_6[70],stage1_5[84]}
   );
   gpc606_5 gpc132 (
      {stage0_5[192], stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[36],stage1_7[58],stage1_6[71],stage1_5[85]}
   );
   gpc606_5 gpc133 (
      {stage0_5[198], stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[37],stage1_7[59],stage1_6[72],stage1_5[86]}
   );
   gpc606_5 gpc134 (
      {stage0_5[204], stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[38],stage1_7[60],stage1_6[73],stage1_5[87]}
   );
   gpc606_5 gpc135 (
      {stage0_5[210], stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[39],stage1_7[61],stage1_6[74],stage1_5[88]}
   );
   gpc606_5 gpc136 (
      {stage0_5[216], stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[40],stage1_7[62],stage1_6[75],stage1_5[89]}
   );
   gpc606_5 gpc137 (
      {stage0_5[222], stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[41],stage1_7[63],stage1_6[76],stage1_5[90]}
   );
   gpc606_5 gpc138 (
      {stage0_5[228], stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[42],stage1_7[64],stage1_6[77],stage1_5[91]}
   );
   gpc606_5 gpc139 (
      {stage0_5[234], stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[43],stage1_7[65],stage1_6[78],stage1_5[92]}
   );
   gpc606_5 gpc140 (
      {stage0_5[240], stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[44],stage1_7[66],stage1_6[79],stage1_5[93]}
   );
   gpc606_5 gpc141 (
      {stage0_5[246], stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[45],stage1_7[67],stage1_6[80],stage1_5[94]}
   );
   gpc606_5 gpc142 (
      {stage0_5[252], stage0_5[253], stage0_5[254], stage0_5[255], 1'b0, 1'b0},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[46],stage1_7[68],stage1_6[81],stage1_5[95]}
   );
   gpc1415_5 gpc143 (
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160]},
      {stage0_7[126]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3]},
      {stage0_9[0]},
      {stage1_10[0],stage1_9[21],stage1_8[47],stage1_7[69],stage1_6[82]}
   );
   gpc606_5 gpc144 (
      {stage0_6[161], stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166]},
      {stage0_8[4], stage0_8[5], stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9]},
      {stage1_10[1],stage1_9[22],stage1_8[48],stage1_7[70],stage1_6[83]}
   );
   gpc606_5 gpc145 (
      {stage0_6[167], stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172]},
      {stage0_8[10], stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage1_10[2],stage1_9[23],stage1_8[49],stage1_7[71],stage1_6[84]}
   );
   gpc606_5 gpc146 (
      {stage0_6[173], stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178]},
      {stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage1_10[3],stage1_9[24],stage1_8[50],stage1_7[72],stage1_6[85]}
   );
   gpc606_5 gpc147 (
      {stage0_6[179], stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184]},
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage1_10[4],stage1_9[25],stage1_8[51],stage1_7[73],stage1_6[86]}
   );
   gpc606_5 gpc148 (
      {stage0_6[185], stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190]},
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage1_10[5],stage1_9[26],stage1_8[52],stage1_7[74],stage1_6[87]}
   );
   gpc606_5 gpc149 (
      {stage0_6[191], stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196]},
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39]},
      {stage1_10[6],stage1_9[27],stage1_8[53],stage1_7[75],stage1_6[88]}
   );
   gpc606_5 gpc150 (
      {stage0_6[197], stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202]},
      {stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45]},
      {stage1_10[7],stage1_9[28],stage1_8[54],stage1_7[76],stage1_6[89]}
   );
   gpc606_5 gpc151 (
      {stage0_6[203], stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208]},
      {stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51]},
      {stage1_10[8],stage1_9[29],stage1_8[55],stage1_7[77],stage1_6[90]}
   );
   gpc606_5 gpc152 (
      {stage0_6[209], stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214]},
      {stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage1_10[9],stage1_9[30],stage1_8[56],stage1_7[78],stage1_6[91]}
   );
   gpc606_5 gpc153 (
      {stage0_6[215], stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220]},
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage1_10[10],stage1_9[31],stage1_8[57],stage1_7[79],stage1_6[92]}
   );
   gpc615_5 gpc154 (
      {stage0_6[221], stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225]},
      {stage0_7[127]},
      {stage0_8[64], stage0_8[65], stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69]},
      {stage1_10[11],stage1_9[32],stage1_8[58],stage1_7[80],stage1_6[93]}
   );
   gpc615_5 gpc155 (
      {stage0_6[226], stage0_6[227], stage0_6[228], stage0_6[229], stage0_6[230]},
      {stage0_7[128]},
      {stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75]},
      {stage1_10[12],stage1_9[33],stage1_8[59],stage1_7[81],stage1_6[94]}
   );
   gpc615_5 gpc156 (
      {stage0_6[231], stage0_6[232], stage0_6[233], stage0_6[234], stage0_6[235]},
      {stage0_7[129]},
      {stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage1_10[13],stage1_9[34],stage1_8[60],stage1_7[82],stage1_6[95]}
   );
   gpc606_5 gpc157 (
      {stage0_7[130], stage0_7[131], stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135]},
      {stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6]},
      {stage1_11[0],stage1_10[14],stage1_9[35],stage1_8[61],stage1_7[83]}
   );
   gpc606_5 gpc158 (
      {stage0_7[136], stage0_7[137], stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141]},
      {stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12]},
      {stage1_11[1],stage1_10[15],stage1_9[36],stage1_8[62],stage1_7[84]}
   );
   gpc606_5 gpc159 (
      {stage0_7[142], stage0_7[143], stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147]},
      {stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18]},
      {stage1_11[2],stage1_10[16],stage1_9[37],stage1_8[63],stage1_7[85]}
   );
   gpc606_5 gpc160 (
      {stage0_7[148], stage0_7[149], stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153]},
      {stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24]},
      {stage1_11[3],stage1_10[17],stage1_9[38],stage1_8[64],stage1_7[86]}
   );
   gpc606_5 gpc161 (
      {stage0_7[154], stage0_7[155], stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159]},
      {stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30]},
      {stage1_11[4],stage1_10[18],stage1_9[39],stage1_8[65],stage1_7[87]}
   );
   gpc606_5 gpc162 (
      {stage0_7[160], stage0_7[161], stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165]},
      {stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36]},
      {stage1_11[5],stage1_10[19],stage1_9[40],stage1_8[66],stage1_7[88]}
   );
   gpc606_5 gpc163 (
      {stage0_7[166], stage0_7[167], stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171]},
      {stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42]},
      {stage1_11[6],stage1_10[20],stage1_9[41],stage1_8[67],stage1_7[89]}
   );
   gpc606_5 gpc164 (
      {stage0_7[172], stage0_7[173], stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177]},
      {stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48]},
      {stage1_11[7],stage1_10[21],stage1_9[42],stage1_8[68],stage1_7[90]}
   );
   gpc606_5 gpc165 (
      {stage0_7[178], stage0_7[179], stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183]},
      {stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54]},
      {stage1_11[8],stage1_10[22],stage1_9[43],stage1_8[69],stage1_7[91]}
   );
   gpc606_5 gpc166 (
      {stage0_7[184], stage0_7[185], stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189]},
      {stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60]},
      {stage1_11[9],stage1_10[23],stage1_9[44],stage1_8[70],stage1_7[92]}
   );
   gpc606_5 gpc167 (
      {stage0_7[190], stage0_7[191], stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195]},
      {stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66]},
      {stage1_11[10],stage1_10[24],stage1_9[45],stage1_8[71],stage1_7[93]}
   );
   gpc615_5 gpc168 (
      {stage0_7[196], stage0_7[197], stage0_7[198], stage0_7[199], stage0_7[200]},
      {stage0_8[82]},
      {stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72]},
      {stage1_11[11],stage1_10[25],stage1_9[46],stage1_8[72],stage1_7[94]}
   );
   gpc615_5 gpc169 (
      {stage0_7[201], stage0_7[202], stage0_7[203], stage0_7[204], stage0_7[205]},
      {stage0_8[83]},
      {stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78]},
      {stage1_11[12],stage1_10[26],stage1_9[47],stage1_8[73],stage1_7[95]}
   );
   gpc615_5 gpc170 (
      {stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209], stage0_7[210]},
      {stage0_8[84]},
      {stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84]},
      {stage1_11[13],stage1_10[27],stage1_9[48],stage1_8[74],stage1_7[96]}
   );
   gpc615_5 gpc171 (
      {stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage0_8[85]},
      {stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90]},
      {stage1_11[14],stage1_10[28],stage1_9[49],stage1_8[75],stage1_7[97]}
   );
   gpc615_5 gpc172 (
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220]},
      {stage0_8[86]},
      {stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96]},
      {stage1_11[15],stage1_10[29],stage1_9[50],stage1_8[76],stage1_7[98]}
   );
   gpc615_5 gpc173 (
      {stage0_7[221], stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225]},
      {stage0_8[87]},
      {stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102]},
      {stage1_11[16],stage1_10[30],stage1_9[51],stage1_8[77],stage1_7[99]}
   );
   gpc615_5 gpc174 (
      {stage0_7[226], stage0_7[227], stage0_7[228], stage0_7[229], stage0_7[230]},
      {stage0_8[88]},
      {stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108]},
      {stage1_11[17],stage1_10[31],stage1_9[52],stage1_8[78],stage1_7[100]}
   );
   gpc615_5 gpc175 (
      {stage0_7[231], stage0_7[232], stage0_7[233], stage0_7[234], stage0_7[235]},
      {stage0_8[89]},
      {stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114]},
      {stage1_11[18],stage1_10[32],stage1_9[53],stage1_8[79],stage1_7[101]}
   );
   gpc615_5 gpc176 (
      {stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239], stage0_7[240]},
      {stage0_8[90]},
      {stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120]},
      {stage1_11[19],stage1_10[33],stage1_9[54],stage1_8[80],stage1_7[102]}
   );
   gpc615_5 gpc177 (
      {stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage0_8[91]},
      {stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126]},
      {stage1_11[20],stage1_10[34],stage1_9[55],stage1_8[81],stage1_7[103]}
   );
   gpc615_5 gpc178 (
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250]},
      {stage0_8[92]},
      {stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131], stage0_9[132]},
      {stage1_11[21],stage1_10[35],stage1_9[56],stage1_8[82],stage1_7[104]}
   );
   gpc606_5 gpc179 (
      {stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[22],stage1_10[36],stage1_9[57],stage1_8[83]}
   );
   gpc606_5 gpc180 (
      {stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[23],stage1_10[37],stage1_9[58],stage1_8[84]}
   );
   gpc606_5 gpc181 (
      {stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[24],stage1_10[38],stage1_9[59],stage1_8[85]}
   );
   gpc606_5 gpc182 (
      {stage0_8[111], stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[25],stage1_10[39],stage1_9[60],stage1_8[86]}
   );
   gpc606_5 gpc183 (
      {stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[26],stage1_10[40],stage1_9[61],stage1_8[87]}
   );
   gpc606_5 gpc184 (
      {stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127], stage0_8[128]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[27],stage1_10[41],stage1_9[62],stage1_8[88]}
   );
   gpc606_5 gpc185 (
      {stage0_8[129], stage0_8[130], stage0_8[131], stage0_8[132], stage0_8[133], stage0_8[134]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[28],stage1_10[42],stage1_9[63],stage1_8[89]}
   );
   gpc606_5 gpc186 (
      {stage0_8[135], stage0_8[136], stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[29],stage1_10[43],stage1_9[64],stage1_8[90]}
   );
   gpc606_5 gpc187 (
      {stage0_8[141], stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[30],stage1_10[44],stage1_9[65],stage1_8[91]}
   );
   gpc606_5 gpc188 (
      {stage0_8[147], stage0_8[148], stage0_8[149], stage0_8[150], stage0_8[151], stage0_8[152]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[31],stage1_10[45],stage1_9[66],stage1_8[92]}
   );
   gpc615_5 gpc189 (
      {stage0_8[153], stage0_8[154], stage0_8[155], stage0_8[156], stage0_8[157]},
      {stage0_9[133]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[32],stage1_10[46],stage1_9[67],stage1_8[93]}
   );
   gpc615_5 gpc190 (
      {stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161], stage0_8[162]},
      {stage0_9[134]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[33],stage1_10[47],stage1_9[68],stage1_8[94]}
   );
   gpc615_5 gpc191 (
      {stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage0_9[135]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[34],stage1_10[48],stage1_9[69],stage1_8[95]}
   );
   gpc615_5 gpc192 (
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172]},
      {stage0_9[136]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[35],stage1_10[49],stage1_9[70],stage1_8[96]}
   );
   gpc615_5 gpc193 (
      {stage0_8[173], stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177]},
      {stage0_9[137]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[36],stage1_10[50],stage1_9[71],stage1_8[97]}
   );
   gpc615_5 gpc194 (
      {stage0_8[178], stage0_8[179], stage0_8[180], stage0_8[181], stage0_8[182]},
      {stage0_9[138]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[37],stage1_10[51],stage1_9[72],stage1_8[98]}
   );
   gpc615_5 gpc195 (
      {stage0_8[183], stage0_8[184], stage0_8[185], stage0_8[186], stage0_8[187]},
      {stage0_9[139]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[38],stage1_10[52],stage1_9[73],stage1_8[99]}
   );
   gpc615_5 gpc196 (
      {stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191], stage0_8[192]},
      {stage0_9[140]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[39],stage1_10[53],stage1_9[74],stage1_8[100]}
   );
   gpc615_5 gpc197 (
      {stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage0_9[141]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[40],stage1_10[54],stage1_9[75],stage1_8[101]}
   );
   gpc615_5 gpc198 (
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202]},
      {stage0_9[142]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[41],stage1_10[55],stage1_9[76],stage1_8[102]}
   );
   gpc615_5 gpc199 (
      {stage0_8[203], stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207]},
      {stage0_9[143]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[42],stage1_10[56],stage1_9[77],stage1_8[103]}
   );
   gpc615_5 gpc200 (
      {stage0_8[208], stage0_8[209], stage0_8[210], stage0_8[211], stage0_8[212]},
      {stage0_9[144]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[43],stage1_10[57],stage1_9[78],stage1_8[104]}
   );
   gpc615_5 gpc201 (
      {stage0_8[213], stage0_8[214], stage0_8[215], stage0_8[216], stage0_8[217]},
      {stage0_9[145]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[44],stage1_10[58],stage1_9[79],stage1_8[105]}
   );
   gpc615_5 gpc202 (
      {stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222]},
      {stage0_9[146]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[45],stage1_10[59],stage1_9[80],stage1_8[106]}
   );
   gpc615_5 gpc203 (
      {stage0_8[223], stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227]},
      {stage0_9[147]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[46],stage1_10[60],stage1_9[81],stage1_8[107]}
   );
   gpc615_5 gpc204 (
      {stage0_8[228], stage0_8[229], stage0_8[230], stage0_8[231], stage0_8[232]},
      {stage0_9[148]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[47],stage1_10[61],stage1_9[82],stage1_8[108]}
   );
   gpc606_5 gpc205 (
      {stage0_9[149], stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[26],stage1_11[48],stage1_10[62],stage1_9[83]}
   );
   gpc606_5 gpc206 (
      {stage0_9[155], stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[27],stage1_11[49],stage1_10[63],stage1_9[84]}
   );
   gpc606_5 gpc207 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165], stage0_9[166]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[28],stage1_11[50],stage1_10[64],stage1_9[85]}
   );
   gpc606_5 gpc208 (
      {stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170], stage0_9[171], stage0_9[172]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[29],stage1_11[51],stage1_10[65],stage1_9[86]}
   );
   gpc606_5 gpc209 (
      {stage0_9[173], stage0_9[174], stage0_9[175], stage0_9[176], stage0_9[177], stage0_9[178]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[30],stage1_11[52],stage1_10[66],stage1_9[87]}
   );
   gpc606_5 gpc210 (
      {stage0_9[179], stage0_9[180], stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[31],stage1_11[53],stage1_10[67],stage1_9[88]}
   );
   gpc615_5 gpc211 (
      {stage0_9[185], stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189]},
      {stage0_10[156]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[32],stage1_11[54],stage1_10[68],stage1_9[89]}
   );
   gpc615_5 gpc212 (
      {stage0_9[190], stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194]},
      {stage0_10[157]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[33],stage1_11[55],stage1_10[69],stage1_9[90]}
   );
   gpc615_5 gpc213 (
      {stage0_9[195], stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199]},
      {stage0_10[158]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[34],stage1_11[56],stage1_10[70],stage1_9[91]}
   );
   gpc615_5 gpc214 (
      {stage0_9[200], stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204]},
      {stage0_10[159]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[35],stage1_11[57],stage1_10[71],stage1_9[92]}
   );
   gpc615_5 gpc215 (
      {stage0_9[205], stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209]},
      {stage0_10[160]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[36],stage1_11[58],stage1_10[72],stage1_9[93]}
   );
   gpc615_5 gpc216 (
      {stage0_9[210], stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214]},
      {stage0_10[161]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[37],stage1_11[59],stage1_10[73],stage1_9[94]}
   );
   gpc615_5 gpc217 (
      {stage0_9[215], stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219]},
      {stage0_10[162]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[38],stage1_11[60],stage1_10[74],stage1_9[95]}
   );
   gpc615_5 gpc218 (
      {stage0_9[220], stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224]},
      {stage0_10[163]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[39],stage1_11[61],stage1_10[75],stage1_9[96]}
   );
   gpc615_5 gpc219 (
      {stage0_9[225], stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229]},
      {stage0_10[164]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[40],stage1_11[62],stage1_10[76],stage1_9[97]}
   );
   gpc615_5 gpc220 (
      {stage0_9[230], stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234]},
      {stage0_10[165]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[41],stage1_11[63],stage1_10[77],stage1_9[98]}
   );
   gpc615_5 gpc221 (
      {stage0_10[166], stage0_10[167], stage0_10[168], stage0_10[169], stage0_10[170]},
      {stage0_11[96]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[16],stage1_12[42],stage1_11[64],stage1_10[78]}
   );
   gpc615_5 gpc222 (
      {stage0_10[171], stage0_10[172], stage0_10[173], stage0_10[174], stage0_10[175]},
      {stage0_11[97]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[17],stage1_12[43],stage1_11[65],stage1_10[79]}
   );
   gpc615_5 gpc223 (
      {stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179], stage0_10[180]},
      {stage0_11[98]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[18],stage1_12[44],stage1_11[66],stage1_10[80]}
   );
   gpc606_5 gpc224 (
      {stage0_11[99], stage0_11[100], stage0_11[101], stage0_11[102], stage0_11[103], stage0_11[104]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[3],stage1_13[19],stage1_12[45],stage1_11[67]}
   );
   gpc606_5 gpc225 (
      {stage0_11[105], stage0_11[106], stage0_11[107], stage0_11[108], stage0_11[109], stage0_11[110]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[4],stage1_13[20],stage1_12[46],stage1_11[68]}
   );
   gpc606_5 gpc226 (
      {stage0_11[111], stage0_11[112], stage0_11[113], stage0_11[114], stage0_11[115], stage0_11[116]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[5],stage1_13[21],stage1_12[47],stage1_11[69]}
   );
   gpc606_5 gpc227 (
      {stage0_11[117], stage0_11[118], stage0_11[119], stage0_11[120], stage0_11[121], stage0_11[122]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[6],stage1_13[22],stage1_12[48],stage1_11[70]}
   );
   gpc606_5 gpc228 (
      {stage0_11[123], stage0_11[124], stage0_11[125], stage0_11[126], stage0_11[127], stage0_11[128]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[7],stage1_13[23],stage1_12[49],stage1_11[71]}
   );
   gpc606_5 gpc229 (
      {stage0_11[129], stage0_11[130], stage0_11[131], stage0_11[132], stage0_11[133], stage0_11[134]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[8],stage1_13[24],stage1_12[50],stage1_11[72]}
   );
   gpc606_5 gpc230 (
      {stage0_11[135], stage0_11[136], stage0_11[137], stage0_11[138], stage0_11[139], stage0_11[140]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[9],stage1_13[25],stage1_12[51],stage1_11[73]}
   );
   gpc606_5 gpc231 (
      {stage0_11[141], stage0_11[142], stage0_11[143], stage0_11[144], stage0_11[145], stage0_11[146]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[10],stage1_13[26],stage1_12[52],stage1_11[74]}
   );
   gpc606_5 gpc232 (
      {stage0_11[147], stage0_11[148], stage0_11[149], stage0_11[150], stage0_11[151], stage0_11[152]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[11],stage1_13[27],stage1_12[53],stage1_11[75]}
   );
   gpc606_5 gpc233 (
      {stage0_11[153], stage0_11[154], stage0_11[155], stage0_11[156], stage0_11[157], stage0_11[158]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[12],stage1_13[28],stage1_12[54],stage1_11[76]}
   );
   gpc606_5 gpc234 (
      {stage0_11[159], stage0_11[160], stage0_11[161], stage0_11[162], stage0_11[163], stage0_11[164]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[13],stage1_13[29],stage1_12[55],stage1_11[77]}
   );
   gpc606_5 gpc235 (
      {stage0_11[165], stage0_11[166], stage0_11[167], stage0_11[168], stage0_11[169], stage0_11[170]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[14],stage1_13[30],stage1_12[56],stage1_11[78]}
   );
   gpc606_5 gpc236 (
      {stage0_11[171], stage0_11[172], stage0_11[173], stage0_11[174], stage0_11[175], stage0_11[176]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[15],stage1_13[31],stage1_12[57],stage1_11[79]}
   );
   gpc606_5 gpc237 (
      {stage0_11[177], stage0_11[178], stage0_11[179], stage0_11[180], stage0_11[181], stage0_11[182]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[16],stage1_13[32],stage1_12[58],stage1_11[80]}
   );
   gpc606_5 gpc238 (
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[14],stage1_14[17],stage1_13[33],stage1_12[59]}
   );
   gpc606_5 gpc239 (
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[15],stage1_14[18],stage1_13[34],stage1_12[60]}
   );
   gpc606_5 gpc240 (
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[16],stage1_14[19],stage1_13[35],stage1_12[61]}
   );
   gpc606_5 gpc241 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[17],stage1_14[20],stage1_13[36],stage1_12[62]}
   );
   gpc606_5 gpc242 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[18],stage1_14[21],stage1_13[37],stage1_12[63]}
   );
   gpc606_5 gpc243 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[19],stage1_14[22],stage1_13[38],stage1_12[64]}
   );
   gpc606_5 gpc244 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[20],stage1_14[23],stage1_13[39],stage1_12[65]}
   );
   gpc606_5 gpc245 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[21],stage1_14[24],stage1_13[40],stage1_12[66]}
   );
   gpc606_5 gpc246 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[22],stage1_14[25],stage1_13[41],stage1_12[67]}
   );
   gpc606_5 gpc247 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[23],stage1_14[26],stage1_13[42],stage1_12[68]}
   );
   gpc606_5 gpc248 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[24],stage1_14[27],stage1_13[43],stage1_12[69]}
   );
   gpc606_5 gpc249 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[25],stage1_14[28],stage1_13[44],stage1_12[70]}
   );
   gpc615_5 gpc250 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94]},
      {stage0_13[84]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[26],stage1_14[29],stage1_13[45],stage1_12[71]}
   );
   gpc615_5 gpc251 (
      {stage0_12[95], stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99]},
      {stage0_13[85]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[27],stage1_14[30],stage1_13[46],stage1_12[72]}
   );
   gpc615_5 gpc252 (
      {stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103], stage0_12[104]},
      {stage0_13[86]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[28],stage1_14[31],stage1_13[47],stage1_12[73]}
   );
   gpc615_5 gpc253 (
      {stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109]},
      {stage0_13[87]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[29],stage1_14[32],stage1_13[48],stage1_12[74]}
   );
   gpc615_5 gpc254 (
      {stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114]},
      {stage0_13[88]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[30],stage1_14[33],stage1_13[49],stage1_12[75]}
   );
   gpc615_5 gpc255 (
      {stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_13[89]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[31],stage1_14[34],stage1_13[50],stage1_12[76]}
   );
   gpc615_5 gpc256 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124]},
      {stage0_13[90]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[32],stage1_14[35],stage1_13[51],stage1_12[77]}
   );
   gpc615_5 gpc257 (
      {stage0_12[125], stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129]},
      {stage0_13[91]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[33],stage1_14[36],stage1_13[52],stage1_12[78]}
   );
   gpc615_5 gpc258 (
      {stage0_12[130], stage0_12[131], stage0_12[132], stage0_12[133], stage0_12[134]},
      {stage0_13[92]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[34],stage1_14[37],stage1_13[53],stage1_12[79]}
   );
   gpc615_5 gpc259 (
      {stage0_12[135], stage0_12[136], stage0_12[137], stage0_12[138], stage0_12[139]},
      {stage0_13[93]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[35],stage1_14[38],stage1_13[54],stage1_12[80]}
   );
   gpc615_5 gpc260 (
      {stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143], stage0_12[144]},
      {stage0_13[94]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[36],stage1_14[39],stage1_13[55],stage1_12[81]}
   );
   gpc615_5 gpc261 (
      {stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage0_13[95]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[37],stage1_14[40],stage1_13[56],stage1_12[82]}
   );
   gpc615_5 gpc262 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154]},
      {stage0_13[96]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[38],stage1_14[41],stage1_13[57],stage1_12[83]}
   );
   gpc615_5 gpc263 (
      {stage0_12[155], stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159]},
      {stage0_13[97]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[39],stage1_14[42],stage1_13[58],stage1_12[84]}
   );
   gpc615_5 gpc264 (
      {stage0_12[160], stage0_12[161], stage0_12[162], stage0_12[163], stage0_12[164]},
      {stage0_13[98]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[40],stage1_14[43],stage1_13[59],stage1_12[85]}
   );
   gpc615_5 gpc265 (
      {stage0_12[165], stage0_12[166], stage0_12[167], stage0_12[168], stage0_12[169]},
      {stage0_13[99]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[41],stage1_14[44],stage1_13[60],stage1_12[86]}
   );
   gpc615_5 gpc266 (
      {stage0_12[170], stage0_12[171], stage0_12[172], stage0_12[173], stage0_12[174]},
      {stage0_13[100]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[42],stage1_14[45],stage1_13[61],stage1_12[87]}
   );
   gpc615_5 gpc267 (
      {stage0_12[175], stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179]},
      {stage0_13[101]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[43],stage1_14[46],stage1_13[62],stage1_12[88]}
   );
   gpc615_5 gpc268 (
      {stage0_12[180], stage0_12[181], stage0_12[182], stage0_12[183], stage0_12[184]},
      {stage0_13[102]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[44],stage1_14[47],stage1_13[63],stage1_12[89]}
   );
   gpc615_5 gpc269 (
      {stage0_12[185], stage0_12[186], stage0_12[187], stage0_12[188], stage0_12[189]},
      {stage0_13[103]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[45],stage1_14[48],stage1_13[64],stage1_12[90]}
   );
   gpc615_5 gpc270 (
      {stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193], stage0_12[194]},
      {stage0_13[104]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[46],stage1_14[49],stage1_13[65],stage1_12[91]}
   );
   gpc615_5 gpc271 (
      {stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199]},
      {stage0_13[105]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[47],stage1_14[50],stage1_13[66],stage1_12[92]}
   );
   gpc615_5 gpc272 (
      {stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203], stage0_12[204]},
      {stage0_13[106]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[48],stage1_14[51],stage1_13[67],stage1_12[93]}
   );
   gpc615_5 gpc273 (
      {stage0_12[205], stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209]},
      {stage0_13[107]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[49],stage1_14[52],stage1_13[68],stage1_12[94]}
   );
   gpc615_5 gpc274 (
      {stage0_12[210], stage0_12[211], stage0_12[212], stage0_12[213], stage0_12[214]},
      {stage0_13[108]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[50],stage1_14[53],stage1_13[69],stage1_12[95]}
   );
   gpc615_5 gpc275 (
      {stage0_12[215], stage0_12[216], stage0_12[217], stage0_12[218], stage0_12[219]},
      {stage0_13[109]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[51],stage1_14[54],stage1_13[70],stage1_12[96]}
   );
   gpc606_5 gpc276 (
      {stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113], stage0_13[114], stage0_13[115]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[38],stage1_15[52],stage1_14[55],stage1_13[71]}
   );
   gpc606_5 gpc277 (
      {stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119], stage0_13[120], stage0_13[121]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[39],stage1_15[53],stage1_14[56],stage1_13[72]}
   );
   gpc606_5 gpc278 (
      {stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125], stage0_13[126], stage0_13[127]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[40],stage1_15[54],stage1_14[57],stage1_13[73]}
   );
   gpc606_5 gpc279 (
      {stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131], stage0_13[132], stage0_13[133]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[41],stage1_15[55],stage1_14[58],stage1_13[74]}
   );
   gpc606_5 gpc280 (
      {stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137], stage0_13[138], stage0_13[139]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[42],stage1_15[56],stage1_14[59],stage1_13[75]}
   );
   gpc606_5 gpc281 (
      {stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143], stage0_13[144], stage0_13[145]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[43],stage1_15[57],stage1_14[60],stage1_13[76]}
   );
   gpc606_5 gpc282 (
      {stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149], stage0_13[150], stage0_13[151]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[44],stage1_15[58],stage1_14[61],stage1_13[77]}
   );
   gpc606_5 gpc283 (
      {stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155], stage0_13[156], stage0_13[157]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[45],stage1_15[59],stage1_14[62],stage1_13[78]}
   );
   gpc606_5 gpc284 (
      {stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161], stage0_13[162], stage0_13[163]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[46],stage1_15[60],stage1_14[63],stage1_13[79]}
   );
   gpc606_5 gpc285 (
      {stage0_13[164], stage0_13[165], stage0_13[166], stage0_13[167], stage0_13[168], stage0_13[169]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[47],stage1_15[61],stage1_14[64],stage1_13[80]}
   );
   gpc606_5 gpc286 (
      {stage0_13[170], stage0_13[171], stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[48],stage1_15[62],stage1_14[65],stage1_13[81]}
   );
   gpc606_5 gpc287 (
      {stage0_13[176], stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[49],stage1_15[63],stage1_14[66],stage1_13[82]}
   );
   gpc606_5 gpc288 (
      {stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186], stage0_13[187]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[50],stage1_15[64],stage1_14[67],stage1_13[83]}
   );
   gpc606_5 gpc289 (
      {stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191], stage0_13[192], stage0_13[193]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[51],stage1_15[65],stage1_14[68],stage1_13[84]}
   );
   gpc606_5 gpc290 (
      {stage0_13[194], stage0_13[195], stage0_13[196], stage0_13[197], stage0_13[198], stage0_13[199]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[52],stage1_15[66],stage1_14[69],stage1_13[85]}
   );
   gpc606_5 gpc291 (
      {stage0_13[200], stage0_13[201], stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[53],stage1_15[67],stage1_14[70],stage1_13[86]}
   );
   gpc606_5 gpc292 (
      {stage0_13[206], stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[54],stage1_15[68],stage1_14[71],stage1_13[87]}
   );
   gpc606_5 gpc293 (
      {stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215], stage0_13[216], stage0_13[217]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[55],stage1_15[69],stage1_14[72],stage1_13[88]}
   );
   gpc606_5 gpc294 (
      {stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221], stage0_13[222], stage0_13[223]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[56],stage1_15[70],stage1_14[73],stage1_13[89]}
   );
   gpc606_5 gpc295 (
      {stage0_13[224], stage0_13[225], stage0_13[226], stage0_13[227], stage0_13[228], stage0_13[229]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[57],stage1_15[71],stage1_14[74],stage1_13[90]}
   );
   gpc606_5 gpc296 (
      {stage0_13[230], stage0_13[231], stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[58],stage1_15[72],stage1_14[75],stage1_13[91]}
   );
   gpc606_5 gpc297 (
      {stage0_13[236], stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240], stage0_13[241]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[59],stage1_15[73],stage1_14[76],stage1_13[92]}
   );
   gpc606_5 gpc298 (
      {stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245], stage0_13[246], stage0_13[247]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[60],stage1_15[74],stage1_14[77],stage1_13[93]}
   );
   gpc606_5 gpc299 (
      {stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251], stage0_13[252], stage0_13[253]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[61],stage1_15[75],stage1_14[78],stage1_13[94]}
   );
   gpc615_5 gpc300 (
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232]},
      {stage0_15[144]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[24],stage1_16[62],stage1_15[76],stage1_14[79]}
   );
   gpc615_5 gpc301 (
      {stage0_14[233], stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237]},
      {stage0_15[145]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[25],stage1_16[63],stage1_15[77],stage1_14[80]}
   );
   gpc615_5 gpc302 (
      {stage0_14[238], stage0_14[239], stage0_14[240], stage0_14[241], stage0_14[242]},
      {stage0_15[146]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[26],stage1_16[64],stage1_15[78],stage1_14[81]}
   );
   gpc615_5 gpc303 (
      {stage0_14[243], stage0_14[244], stage0_14[245], stage0_14[246], stage0_14[247]},
      {stage0_15[147]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[27],stage1_16[65],stage1_15[79],stage1_14[82]}
   );
   gpc615_5 gpc304 (
      {stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251], stage0_14[252]},
      {stage0_15[148]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[28],stage1_16[66],stage1_15[80],stage1_14[83]}
   );
   gpc615_5 gpc305 (
      {stage0_14[253], stage0_14[254], stage0_14[255], 1'b0, 1'b0},
      {stage0_15[149]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[29],stage1_16[67],stage1_15[81],stage1_14[84]}
   );
   gpc615_5 gpc306 (
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154]},
      {stage0_16[36]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[6],stage1_17[30],stage1_16[68],stage1_15[82]}
   );
   gpc615_5 gpc307 (
      {stage0_15[155], stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159]},
      {stage0_16[37]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[7],stage1_17[31],stage1_16[69],stage1_15[83]}
   );
   gpc615_5 gpc308 (
      {stage0_15[160], stage0_15[161], stage0_15[162], stage0_15[163], stage0_15[164]},
      {stage0_16[38]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[8],stage1_17[32],stage1_16[70],stage1_15[84]}
   );
   gpc615_5 gpc309 (
      {stage0_15[165], stage0_15[166], stage0_15[167], stage0_15[168], stage0_15[169]},
      {stage0_16[39]},
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage1_19[3],stage1_18[9],stage1_17[33],stage1_16[71],stage1_15[85]}
   );
   gpc615_5 gpc310 (
      {stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173], stage0_15[174]},
      {stage0_16[40]},
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage1_19[4],stage1_18[10],stage1_17[34],stage1_16[72],stage1_15[86]}
   );
   gpc615_5 gpc311 (
      {stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage0_16[41]},
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage1_19[5],stage1_18[11],stage1_17[35],stage1_16[73],stage1_15[87]}
   );
   gpc615_5 gpc312 (
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184]},
      {stage0_16[42]},
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage1_19[6],stage1_18[12],stage1_17[36],stage1_16[74],stage1_15[88]}
   );
   gpc615_5 gpc313 (
      {stage0_15[185], stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189]},
      {stage0_16[43]},
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage1_19[7],stage1_18[13],stage1_17[37],stage1_16[75],stage1_15[89]}
   );
   gpc615_5 gpc314 (
      {stage0_15[190], stage0_15[191], stage0_15[192], stage0_15[193], stage0_15[194]},
      {stage0_16[44]},
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage1_19[8],stage1_18[14],stage1_17[38],stage1_16[76],stage1_15[90]}
   );
   gpc615_5 gpc315 (
      {stage0_15[195], stage0_15[196], stage0_15[197], stage0_15[198], stage0_15[199]},
      {stage0_16[45]},
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage1_19[9],stage1_18[15],stage1_17[39],stage1_16[77],stage1_15[91]}
   );
   gpc615_5 gpc316 (
      {stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203], stage0_15[204]},
      {stage0_16[46]},
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage1_19[10],stage1_18[16],stage1_17[40],stage1_16[78],stage1_15[92]}
   );
   gpc615_5 gpc317 (
      {stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage0_16[47]},
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage1_19[11],stage1_18[17],stage1_17[41],stage1_16[79],stage1_15[93]}
   );
   gpc615_5 gpc318 (
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214]},
      {stage0_16[48]},
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage1_19[12],stage1_18[18],stage1_17[42],stage1_16[80],stage1_15[94]}
   );
   gpc615_5 gpc319 (
      {stage0_15[215], stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219]},
      {stage0_16[49]},
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage1_19[13],stage1_18[19],stage1_17[43],stage1_16[81],stage1_15[95]}
   );
   gpc606_5 gpc320 (
      {stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53], stage0_16[54], stage0_16[55]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[14],stage1_18[20],stage1_17[44],stage1_16[82]}
   );
   gpc606_5 gpc321 (
      {stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59], stage0_16[60], stage0_16[61]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[15],stage1_18[21],stage1_17[45],stage1_16[83]}
   );
   gpc606_5 gpc322 (
      {stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65], stage0_16[66], stage0_16[67]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[16],stage1_18[22],stage1_17[46],stage1_16[84]}
   );
   gpc606_5 gpc323 (
      {stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71], stage0_16[72], stage0_16[73]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[17],stage1_18[23],stage1_17[47],stage1_16[85]}
   );
   gpc606_5 gpc324 (
      {stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78], stage0_16[79]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[18],stage1_18[24],stage1_17[48],stage1_16[86]}
   );
   gpc606_5 gpc325 (
      {stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84], stage0_16[85]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[19],stage1_18[25],stage1_17[49],stage1_16[87]}
   );
   gpc606_5 gpc326 (
      {stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[20],stage1_18[26],stage1_17[50],stage1_16[88]}
   );
   gpc606_5 gpc327 (
      {stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[21],stage1_18[27],stage1_17[51],stage1_16[89]}
   );
   gpc606_5 gpc328 (
      {stage0_16[98], stage0_16[99], stage0_16[100], stage0_16[101], stage0_16[102], stage0_16[103]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[22],stage1_18[28],stage1_17[52],stage1_16[90]}
   );
   gpc606_5 gpc329 (
      {stage0_16[104], stage0_16[105], stage0_16[106], stage0_16[107], stage0_16[108], stage0_16[109]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[23],stage1_18[29],stage1_17[53],stage1_16[91]}
   );
   gpc606_5 gpc330 (
      {stage0_16[110], stage0_16[111], stage0_16[112], stage0_16[113], stage0_16[114], stage0_16[115]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[24],stage1_18[30],stage1_17[54],stage1_16[92]}
   );
   gpc606_5 gpc331 (
      {stage0_16[116], stage0_16[117], stage0_16[118], stage0_16[119], stage0_16[120], stage0_16[121]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[25],stage1_18[31],stage1_17[55],stage1_16[93]}
   );
   gpc606_5 gpc332 (
      {stage0_16[122], stage0_16[123], stage0_16[124], stage0_16[125], stage0_16[126], stage0_16[127]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[26],stage1_18[32],stage1_17[56],stage1_16[94]}
   );
   gpc606_5 gpc333 (
      {stage0_16[128], stage0_16[129], stage0_16[130], stage0_16[131], stage0_16[132], stage0_16[133]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[27],stage1_18[33],stage1_17[57],stage1_16[95]}
   );
   gpc606_5 gpc334 (
      {stage0_16[134], stage0_16[135], stage0_16[136], stage0_16[137], stage0_16[138], stage0_16[139]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[28],stage1_18[34],stage1_17[58],stage1_16[96]}
   );
   gpc606_5 gpc335 (
      {stage0_16[140], stage0_16[141], stage0_16[142], stage0_16[143], stage0_16[144], stage0_16[145]},
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94], stage0_18[95]},
      {stage1_20[15],stage1_19[29],stage1_18[35],stage1_17[59],stage1_16[97]}
   );
   gpc606_5 gpc336 (
      {stage0_16[146], stage0_16[147], stage0_16[148], stage0_16[149], stage0_16[150], stage0_16[151]},
      {stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99], stage0_18[100], stage0_18[101]},
      {stage1_20[16],stage1_19[30],stage1_18[36],stage1_17[60],stage1_16[98]}
   );
   gpc606_5 gpc337 (
      {stage0_16[152], stage0_16[153], stage0_16[154], stage0_16[155], stage0_16[156], stage0_16[157]},
      {stage0_18[102], stage0_18[103], stage0_18[104], stage0_18[105], stage0_18[106], stage0_18[107]},
      {stage1_20[17],stage1_19[31],stage1_18[37],stage1_17[61],stage1_16[99]}
   );
   gpc606_5 gpc338 (
      {stage0_16[158], stage0_16[159], stage0_16[160], stage0_16[161], stage0_16[162], stage0_16[163]},
      {stage0_18[108], stage0_18[109], stage0_18[110], stage0_18[111], stage0_18[112], stage0_18[113]},
      {stage1_20[18],stage1_19[32],stage1_18[38],stage1_17[62],stage1_16[100]}
   );
   gpc606_5 gpc339 (
      {stage0_16[164], stage0_16[165], stage0_16[166], stage0_16[167], stage0_16[168], stage0_16[169]},
      {stage0_18[114], stage0_18[115], stage0_18[116], stage0_18[117], stage0_18[118], stage0_18[119]},
      {stage1_20[19],stage1_19[33],stage1_18[39],stage1_17[63],stage1_16[101]}
   );
   gpc615_5 gpc340 (
      {stage0_16[170], stage0_16[171], stage0_16[172], stage0_16[173], stage0_16[174]},
      {stage0_17[84]},
      {stage0_18[120], stage0_18[121], stage0_18[122], stage0_18[123], stage0_18[124], stage0_18[125]},
      {stage1_20[20],stage1_19[34],stage1_18[40],stage1_17[64],stage1_16[102]}
   );
   gpc615_5 gpc341 (
      {stage0_16[175], stage0_16[176], stage0_16[177], stage0_16[178], stage0_16[179]},
      {stage0_17[85]},
      {stage0_18[126], stage0_18[127], stage0_18[128], stage0_18[129], stage0_18[130], stage0_18[131]},
      {stage1_20[21],stage1_19[35],stage1_18[41],stage1_17[65],stage1_16[103]}
   );
   gpc615_5 gpc342 (
      {stage0_16[180], stage0_16[181], stage0_16[182], stage0_16[183], stage0_16[184]},
      {stage0_17[86]},
      {stage0_18[132], stage0_18[133], stage0_18[134], stage0_18[135], stage0_18[136], stage0_18[137]},
      {stage1_20[22],stage1_19[36],stage1_18[42],stage1_17[66],stage1_16[104]}
   );
   gpc615_5 gpc343 (
      {stage0_16[185], stage0_16[186], stage0_16[187], stage0_16[188], stage0_16[189]},
      {stage0_17[87]},
      {stage0_18[138], stage0_18[139], stage0_18[140], stage0_18[141], stage0_18[142], stage0_18[143]},
      {stage1_20[23],stage1_19[37],stage1_18[43],stage1_17[67],stage1_16[105]}
   );
   gpc615_5 gpc344 (
      {stage0_16[190], stage0_16[191], stage0_16[192], stage0_16[193], stage0_16[194]},
      {stage0_17[88]},
      {stage0_18[144], stage0_18[145], stage0_18[146], stage0_18[147], stage0_18[148], stage0_18[149]},
      {stage1_20[24],stage1_19[38],stage1_18[44],stage1_17[68],stage1_16[106]}
   );
   gpc615_5 gpc345 (
      {stage0_16[195], stage0_16[196], stage0_16[197], stage0_16[198], stage0_16[199]},
      {stage0_17[89]},
      {stage0_18[150], stage0_18[151], stage0_18[152], stage0_18[153], stage0_18[154], stage0_18[155]},
      {stage1_20[25],stage1_19[39],stage1_18[45],stage1_17[69],stage1_16[107]}
   );
   gpc615_5 gpc346 (
      {stage0_16[200], stage0_16[201], stage0_16[202], stage0_16[203], stage0_16[204]},
      {stage0_17[90]},
      {stage0_18[156], stage0_18[157], stage0_18[158], stage0_18[159], stage0_18[160], stage0_18[161]},
      {stage1_20[26],stage1_19[40],stage1_18[46],stage1_17[70],stage1_16[108]}
   );
   gpc615_5 gpc347 (
      {stage0_16[205], stage0_16[206], stage0_16[207], stage0_16[208], stage0_16[209]},
      {stage0_17[91]},
      {stage0_18[162], stage0_18[163], stage0_18[164], stage0_18[165], stage0_18[166], stage0_18[167]},
      {stage1_20[27],stage1_19[41],stage1_18[47],stage1_17[71],stage1_16[109]}
   );
   gpc615_5 gpc348 (
      {stage0_16[210], stage0_16[211], stage0_16[212], stage0_16[213], stage0_16[214]},
      {stage0_17[92]},
      {stage0_18[168], stage0_18[169], stage0_18[170], stage0_18[171], stage0_18[172], stage0_18[173]},
      {stage1_20[28],stage1_19[42],stage1_18[48],stage1_17[72],stage1_16[110]}
   );
   gpc615_5 gpc349 (
      {stage0_16[215], stage0_16[216], stage0_16[217], stage0_16[218], stage0_16[219]},
      {stage0_17[93]},
      {stage0_18[174], stage0_18[175], stage0_18[176], stage0_18[177], stage0_18[178], stage0_18[179]},
      {stage1_20[29],stage1_19[43],stage1_18[49],stage1_17[73],stage1_16[111]}
   );
   gpc615_5 gpc350 (
      {stage0_16[220], stage0_16[221], stage0_16[222], stage0_16[223], stage0_16[224]},
      {stage0_17[94]},
      {stage0_18[180], stage0_18[181], stage0_18[182], stage0_18[183], stage0_18[184], stage0_18[185]},
      {stage1_20[30],stage1_19[44],stage1_18[50],stage1_17[74],stage1_16[112]}
   );
   gpc615_5 gpc351 (
      {stage0_16[225], stage0_16[226], stage0_16[227], stage0_16[228], stage0_16[229]},
      {stage0_17[95]},
      {stage0_18[186], stage0_18[187], stage0_18[188], stage0_18[189], stage0_18[190], stage0_18[191]},
      {stage1_20[31],stage1_19[45],stage1_18[51],stage1_17[75],stage1_16[113]}
   );
   gpc615_5 gpc352 (
      {stage0_16[230], stage0_16[231], stage0_16[232], stage0_16[233], stage0_16[234]},
      {stage0_17[96]},
      {stage0_18[192], stage0_18[193], stage0_18[194], stage0_18[195], stage0_18[196], stage0_18[197]},
      {stage1_20[32],stage1_19[46],stage1_18[52],stage1_17[76],stage1_16[114]}
   );
   gpc615_5 gpc353 (
      {stage0_16[235], stage0_16[236], stage0_16[237], stage0_16[238], stage0_16[239]},
      {stage0_17[97]},
      {stage0_18[198], stage0_18[199], stage0_18[200], stage0_18[201], stage0_18[202], stage0_18[203]},
      {stage1_20[33],stage1_19[47],stage1_18[53],stage1_17[77],stage1_16[115]}
   );
   gpc615_5 gpc354 (
      {stage0_16[240], stage0_16[241], stage0_16[242], stage0_16[243], stage0_16[244]},
      {stage0_17[98]},
      {stage0_18[204], stage0_18[205], stage0_18[206], stage0_18[207], stage0_18[208], stage0_18[209]},
      {stage1_20[34],stage1_19[48],stage1_18[54],stage1_17[78],stage1_16[116]}
   );
   gpc615_5 gpc355 (
      {stage0_16[245], stage0_16[246], stage0_16[247], stage0_16[248], stage0_16[249]},
      {stage0_17[99]},
      {stage0_18[210], stage0_18[211], stage0_18[212], stage0_18[213], stage0_18[214], stage0_18[215]},
      {stage1_20[35],stage1_19[49],stage1_18[55],stage1_17[79],stage1_16[117]}
   );
   gpc615_5 gpc356 (
      {stage0_16[250], stage0_16[251], stage0_16[252], stage0_16[253], stage0_16[254]},
      {stage0_17[100]},
      {stage0_18[216], stage0_18[217], stage0_18[218], stage0_18[219], stage0_18[220], stage0_18[221]},
      {stage1_20[36],stage1_19[50],stage1_18[56],stage1_17[80],stage1_16[118]}
   );
   gpc606_5 gpc357 (
      {stage0_17[101], stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[37],stage1_19[51],stage1_18[57],stage1_17[81]}
   );
   gpc606_5 gpc358 (
      {stage0_17[107], stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[38],stage1_19[52],stage1_18[58],stage1_17[82]}
   );
   gpc606_5 gpc359 (
      {stage0_17[113], stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[39],stage1_19[53],stage1_18[59],stage1_17[83]}
   );
   gpc606_5 gpc360 (
      {stage0_17[119], stage0_17[120], stage0_17[121], stage0_17[122], stage0_17[123], stage0_17[124]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[40],stage1_19[54],stage1_18[60],stage1_17[84]}
   );
   gpc606_5 gpc361 (
      {stage0_17[125], stage0_17[126], stage0_17[127], stage0_17[128], stage0_17[129], stage0_17[130]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[41],stage1_19[55],stage1_18[61],stage1_17[85]}
   );
   gpc606_5 gpc362 (
      {stage0_17[131], stage0_17[132], stage0_17[133], stage0_17[134], stage0_17[135], stage0_17[136]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[42],stage1_19[56],stage1_18[62],stage1_17[86]}
   );
   gpc606_5 gpc363 (
      {stage0_17[137], stage0_17[138], stage0_17[139], stage0_17[140], stage0_17[141], stage0_17[142]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[43],stage1_19[57],stage1_18[63],stage1_17[87]}
   );
   gpc606_5 gpc364 (
      {stage0_17[143], stage0_17[144], stage0_17[145], stage0_17[146], stage0_17[147], stage0_17[148]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[44],stage1_19[58],stage1_18[64],stage1_17[88]}
   );
   gpc606_5 gpc365 (
      {stage0_17[149], stage0_17[150], stage0_17[151], stage0_17[152], stage0_17[153], stage0_17[154]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[45],stage1_19[59],stage1_18[65],stage1_17[89]}
   );
   gpc606_5 gpc366 (
      {stage0_17[155], stage0_17[156], stage0_17[157], stage0_17[158], stage0_17[159], stage0_17[160]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[46],stage1_19[60],stage1_18[66],stage1_17[90]}
   );
   gpc606_5 gpc367 (
      {stage0_17[161], stage0_17[162], stage0_17[163], stage0_17[164], stage0_17[165], stage0_17[166]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[47],stage1_19[61],stage1_18[67],stage1_17[91]}
   );
   gpc606_5 gpc368 (
      {stage0_17[167], stage0_17[168], stage0_17[169], stage0_17[170], stage0_17[171], stage0_17[172]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[48],stage1_19[62],stage1_18[68],stage1_17[92]}
   );
   gpc606_5 gpc369 (
      {stage0_17[173], stage0_17[174], stage0_17[175], stage0_17[176], stage0_17[177], stage0_17[178]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[49],stage1_19[63],stage1_18[69],stage1_17[93]}
   );
   gpc606_5 gpc370 (
      {stage0_17[179], stage0_17[180], stage0_17[181], stage0_17[182], stage0_17[183], stage0_17[184]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[50],stage1_19[64],stage1_18[70],stage1_17[94]}
   );
   gpc606_5 gpc371 (
      {stage0_17[185], stage0_17[186], stage0_17[187], stage0_17[188], stage0_17[189], stage0_17[190]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[51],stage1_19[65],stage1_18[71],stage1_17[95]}
   );
   gpc606_5 gpc372 (
      {stage0_17[191], stage0_17[192], stage0_17[193], stage0_17[194], stage0_17[195], stage0_17[196]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[52],stage1_19[66],stage1_18[72],stage1_17[96]}
   );
   gpc606_5 gpc373 (
      {stage0_17[197], stage0_17[198], stage0_17[199], stage0_17[200], stage0_17[201], stage0_17[202]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[53],stage1_19[67],stage1_18[73],stage1_17[97]}
   );
   gpc606_5 gpc374 (
      {stage0_17[203], stage0_17[204], stage0_17[205], stage0_17[206], stage0_17[207], stage0_17[208]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[54],stage1_19[68],stage1_18[74],stage1_17[98]}
   );
   gpc606_5 gpc375 (
      {stage0_17[209], stage0_17[210], stage0_17[211], stage0_17[212], stage0_17[213], stage0_17[214]},
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113]},
      {stage1_21[18],stage1_20[55],stage1_19[69],stage1_18[75],stage1_17[99]}
   );
   gpc606_5 gpc376 (
      {stage0_17[215], stage0_17[216], stage0_17[217], stage0_17[218], stage0_17[219], stage0_17[220]},
      {stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage1_21[19],stage1_20[56],stage1_19[70],stage1_18[76],stage1_17[100]}
   );
   gpc606_5 gpc377 (
      {stage0_17[221], stage0_17[222], stage0_17[223], stage0_17[224], stage0_17[225], stage0_17[226]},
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124], stage0_19[125]},
      {stage1_21[20],stage1_20[57],stage1_19[71],stage1_18[77],stage1_17[101]}
   );
   gpc606_5 gpc378 (
      {stage0_17[227], stage0_17[228], stage0_17[229], stage0_17[230], stage0_17[231], stage0_17[232]},
      {stage0_19[126], stage0_19[127], stage0_19[128], stage0_19[129], stage0_19[130], stage0_19[131]},
      {stage1_21[21],stage1_20[58],stage1_19[72],stage1_18[78],stage1_17[102]}
   );
   gpc606_5 gpc379 (
      {stage0_17[233], stage0_17[234], stage0_17[235], stage0_17[236], stage0_17[237], stage0_17[238]},
      {stage0_19[132], stage0_19[133], stage0_19[134], stage0_19[135], stage0_19[136], stage0_19[137]},
      {stage1_21[22],stage1_20[59],stage1_19[73],stage1_18[79],stage1_17[103]}
   );
   gpc606_5 gpc380 (
      {stage0_17[239], stage0_17[240], stage0_17[241], stage0_17[242], stage0_17[243], stage0_17[244]},
      {stage0_19[138], stage0_19[139], stage0_19[140], stage0_19[141], stage0_19[142], stage0_19[143]},
      {stage1_21[23],stage1_20[60],stage1_19[74],stage1_18[80],stage1_17[104]}
   );
   gpc606_5 gpc381 (
      {stage0_17[245], stage0_17[246], stage0_17[247], stage0_17[248], stage0_17[249], stage0_17[250]},
      {stage0_19[144], stage0_19[145], stage0_19[146], stage0_19[147], stage0_19[148], stage0_19[149]},
      {stage1_21[24],stage1_20[61],stage1_19[75],stage1_18[81],stage1_17[105]}
   );
   gpc615_5 gpc382 (
      {stage0_18[222], stage0_18[223], stage0_18[224], stage0_18[225], stage0_18[226]},
      {stage0_19[150]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[25],stage1_20[62],stage1_19[76],stage1_18[82]}
   );
   gpc615_5 gpc383 (
      {stage0_18[227], stage0_18[228], stage0_18[229], stage0_18[230], stage0_18[231]},
      {stage0_19[151]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[26],stage1_20[63],stage1_19[77],stage1_18[83]}
   );
   gpc615_5 gpc384 (
      {stage0_18[232], stage0_18[233], stage0_18[234], stage0_18[235], stage0_18[236]},
      {stage0_19[152]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[27],stage1_20[64],stage1_19[78],stage1_18[84]}
   );
   gpc615_5 gpc385 (
      {stage0_18[237], stage0_18[238], stage0_18[239], stage0_18[240], stage0_18[241]},
      {stage0_19[153]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[28],stage1_20[65],stage1_19[79],stage1_18[85]}
   );
   gpc615_5 gpc386 (
      {stage0_19[154], stage0_19[155], stage0_19[156], stage0_19[157], stage0_19[158]},
      {stage0_20[24]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[4],stage1_21[29],stage1_20[66],stage1_19[80]}
   );
   gpc615_5 gpc387 (
      {stage0_19[159], stage0_19[160], stage0_19[161], stage0_19[162], stage0_19[163]},
      {stage0_20[25]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[5],stage1_21[30],stage1_20[67],stage1_19[81]}
   );
   gpc615_5 gpc388 (
      {stage0_19[164], stage0_19[165], stage0_19[166], stage0_19[167], stage0_19[168]},
      {stage0_20[26]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[6],stage1_21[31],stage1_20[68],stage1_19[82]}
   );
   gpc615_5 gpc389 (
      {stage0_19[169], stage0_19[170], stage0_19[171], stage0_19[172], stage0_19[173]},
      {stage0_20[27]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[7],stage1_21[32],stage1_20[69],stage1_19[83]}
   );
   gpc615_5 gpc390 (
      {stage0_19[174], stage0_19[175], stage0_19[176], stage0_19[177], stage0_19[178]},
      {stage0_20[28]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[8],stage1_21[33],stage1_20[70],stage1_19[84]}
   );
   gpc615_5 gpc391 (
      {stage0_19[179], stage0_19[180], stage0_19[181], stage0_19[182], stage0_19[183]},
      {stage0_20[29]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[9],stage1_21[34],stage1_20[71],stage1_19[85]}
   );
   gpc615_5 gpc392 (
      {stage0_19[184], stage0_19[185], stage0_19[186], stage0_19[187], stage0_19[188]},
      {stage0_20[30]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[10],stage1_21[35],stage1_20[72],stage1_19[86]}
   );
   gpc615_5 gpc393 (
      {stage0_19[189], stage0_19[190], stage0_19[191], stage0_19[192], stage0_19[193]},
      {stage0_20[31]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[11],stage1_21[36],stage1_20[73],stage1_19[87]}
   );
   gpc615_5 gpc394 (
      {stage0_19[194], stage0_19[195], stage0_19[196], stage0_19[197], stage0_19[198]},
      {stage0_20[32]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[12],stage1_21[37],stage1_20[74],stage1_19[88]}
   );
   gpc615_5 gpc395 (
      {stage0_19[199], stage0_19[200], stage0_19[201], stage0_19[202], stage0_19[203]},
      {stage0_20[33]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[13],stage1_21[38],stage1_20[75],stage1_19[89]}
   );
   gpc615_5 gpc396 (
      {stage0_19[204], stage0_19[205], stage0_19[206], stage0_19[207], stage0_19[208]},
      {stage0_20[34]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[14],stage1_21[39],stage1_20[76],stage1_19[90]}
   );
   gpc615_5 gpc397 (
      {stage0_19[209], stage0_19[210], stage0_19[211], stage0_19[212], stage0_19[213]},
      {stage0_20[35]},
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage1_23[11],stage1_22[15],stage1_21[40],stage1_20[77],stage1_19[91]}
   );
   gpc615_5 gpc398 (
      {stage0_19[214], stage0_19[215], stage0_19[216], stage0_19[217], stage0_19[218]},
      {stage0_20[36]},
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage1_23[12],stage1_22[16],stage1_21[41],stage1_20[78],stage1_19[92]}
   );
   gpc615_5 gpc399 (
      {stage0_19[219], stage0_19[220], stage0_19[221], stage0_19[222], stage0_19[223]},
      {stage0_20[37]},
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage1_23[13],stage1_22[17],stage1_21[42],stage1_20[79],stage1_19[93]}
   );
   gpc1343_5 gpc400 (
      {stage0_20[38], stage0_20[39], stage0_20[40]},
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87]},
      {stage0_22[0], stage0_22[1], stage0_22[2]},
      {stage0_23[0]},
      {stage1_24[0],stage1_23[14],stage1_22[18],stage1_21[43],stage1_20[80]}
   );
   gpc1343_5 gpc401 (
      {stage0_20[41], stage0_20[42], stage0_20[43]},
      {stage0_21[88], stage0_21[89], stage0_21[90], stage0_21[91]},
      {stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage0_23[1]},
      {stage1_24[1],stage1_23[15],stage1_22[19],stage1_21[44],stage1_20[81]}
   );
   gpc1343_5 gpc402 (
      {stage0_20[44], stage0_20[45], stage0_20[46]},
      {stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_22[6], stage0_22[7], stage0_22[8]},
      {stage0_23[2]},
      {stage1_24[2],stage1_23[16],stage1_22[20],stage1_21[45],stage1_20[82]}
   );
   gpc1343_5 gpc403 (
      {stage0_20[47], stage0_20[48], stage0_20[49]},
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99]},
      {stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage0_23[3]},
      {stage1_24[3],stage1_23[17],stage1_22[21],stage1_21[46],stage1_20[83]}
   );
   gpc1343_5 gpc404 (
      {stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[100], stage0_21[101], stage0_21[102], stage0_21[103]},
      {stage0_22[12], stage0_22[13], stage0_22[14]},
      {stage0_23[4]},
      {stage1_24[4],stage1_23[18],stage1_22[22],stage1_21[47],stage1_20[84]}
   );
   gpc1343_5 gpc405 (
      {stage0_20[53], stage0_20[54], stage0_20[55]},
      {stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage0_23[5]},
      {stage1_24[5],stage1_23[19],stage1_22[23],stage1_21[48],stage1_20[85]}
   );
   gpc1343_5 gpc406 (
      {stage0_20[56], stage0_20[57], stage0_20[58]},
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111]},
      {stage0_22[18], stage0_22[19], stage0_22[20]},
      {stage0_23[6]},
      {stage1_24[6],stage1_23[20],stage1_22[24],stage1_21[49],stage1_20[86]}
   );
   gpc1343_5 gpc407 (
      {stage0_20[59], stage0_20[60], stage0_20[61]},
      {stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115]},
      {stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage0_23[7]},
      {stage1_24[7],stage1_23[21],stage1_22[25],stage1_21[50],stage1_20[87]}
   );
   gpc1343_5 gpc408 (
      {stage0_20[62], stage0_20[63], stage0_20[64]},
      {stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_22[24], stage0_22[25], stage0_22[26]},
      {stage0_23[8]},
      {stage1_24[8],stage1_23[22],stage1_22[26],stage1_21[51],stage1_20[88]}
   );
   gpc606_5 gpc409 (
      {stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68], stage0_20[69], stage0_20[70]},
      {stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30], stage0_22[31], stage0_22[32]},
      {stage1_24[9],stage1_23[23],stage1_22[27],stage1_21[52],stage1_20[89]}
   );
   gpc606_5 gpc410 (
      {stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74], stage0_20[75], stage0_20[76]},
      {stage0_22[33], stage0_22[34], stage0_22[35], stage0_22[36], stage0_22[37], stage0_22[38]},
      {stage1_24[10],stage1_23[24],stage1_22[28],stage1_21[53],stage1_20[90]}
   );
   gpc606_5 gpc411 (
      {stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81], stage0_20[82]},
      {stage0_22[39], stage0_22[40], stage0_22[41], stage0_22[42], stage0_22[43], stage0_22[44]},
      {stage1_24[11],stage1_23[25],stage1_22[29],stage1_21[54],stage1_20[91]}
   );
   gpc606_5 gpc412 (
      {stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87], stage0_20[88]},
      {stage0_22[45], stage0_22[46], stage0_22[47], stage0_22[48], stage0_22[49], stage0_22[50]},
      {stage1_24[12],stage1_23[26],stage1_22[30],stage1_21[55],stage1_20[92]}
   );
   gpc606_5 gpc413 (
      {stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93], stage0_20[94]},
      {stage0_22[51], stage0_22[52], stage0_22[53], stage0_22[54], stage0_22[55], stage0_22[56]},
      {stage1_24[13],stage1_23[27],stage1_22[31],stage1_21[56],stage1_20[93]}
   );
   gpc606_5 gpc414 (
      {stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98], stage0_20[99], stage0_20[100]},
      {stage0_22[57], stage0_22[58], stage0_22[59], stage0_22[60], stage0_22[61], stage0_22[62]},
      {stage1_24[14],stage1_23[28],stage1_22[32],stage1_21[57],stage1_20[94]}
   );
   gpc606_5 gpc415 (
      {stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104], stage0_20[105], stage0_20[106]},
      {stage0_22[63], stage0_22[64], stage0_22[65], stage0_22[66], stage0_22[67], stage0_22[68]},
      {stage1_24[15],stage1_23[29],stage1_22[33],stage1_21[58],stage1_20[95]}
   );
   gpc606_5 gpc416 (
      {stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110], stage0_20[111], stage0_20[112]},
      {stage0_22[69], stage0_22[70], stage0_22[71], stage0_22[72], stage0_22[73], stage0_22[74]},
      {stage1_24[16],stage1_23[30],stage1_22[34],stage1_21[59],stage1_20[96]}
   );
   gpc606_5 gpc417 (
      {stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116], stage0_20[117], stage0_20[118]},
      {stage0_22[75], stage0_22[76], stage0_22[77], stage0_22[78], stage0_22[79], stage0_22[80]},
      {stage1_24[17],stage1_23[31],stage1_22[35],stage1_21[60],stage1_20[97]}
   );
   gpc606_5 gpc418 (
      {stage0_20[119], stage0_20[120], stage0_20[121], stage0_20[122], stage0_20[123], stage0_20[124]},
      {stage0_22[81], stage0_22[82], stage0_22[83], stage0_22[84], stage0_22[85], stage0_22[86]},
      {stage1_24[18],stage1_23[32],stage1_22[36],stage1_21[61],stage1_20[98]}
   );
   gpc606_5 gpc419 (
      {stage0_20[125], stage0_20[126], stage0_20[127], stage0_20[128], stage0_20[129], stage0_20[130]},
      {stage0_22[87], stage0_22[88], stage0_22[89], stage0_22[90], stage0_22[91], stage0_22[92]},
      {stage1_24[19],stage1_23[33],stage1_22[37],stage1_21[62],stage1_20[99]}
   );
   gpc606_5 gpc420 (
      {stage0_20[131], stage0_20[132], stage0_20[133], stage0_20[134], stage0_20[135], stage0_20[136]},
      {stage0_22[93], stage0_22[94], stage0_22[95], stage0_22[96], stage0_22[97], stage0_22[98]},
      {stage1_24[20],stage1_23[34],stage1_22[38],stage1_21[63],stage1_20[100]}
   );
   gpc606_5 gpc421 (
      {stage0_20[137], stage0_20[138], stage0_20[139], stage0_20[140], stage0_20[141], stage0_20[142]},
      {stage0_22[99], stage0_22[100], stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104]},
      {stage1_24[21],stage1_23[35],stage1_22[39],stage1_21[64],stage1_20[101]}
   );
   gpc606_5 gpc422 (
      {stage0_20[143], stage0_20[144], stage0_20[145], stage0_20[146], stage0_20[147], stage0_20[148]},
      {stage0_22[105], stage0_22[106], stage0_22[107], stage0_22[108], stage0_22[109], stage0_22[110]},
      {stage1_24[22],stage1_23[36],stage1_22[40],stage1_21[65],stage1_20[102]}
   );
   gpc606_5 gpc423 (
      {stage0_20[149], stage0_20[150], stage0_20[151], stage0_20[152], stage0_20[153], stage0_20[154]},
      {stage0_22[111], stage0_22[112], stage0_22[113], stage0_22[114], stage0_22[115], stage0_22[116]},
      {stage1_24[23],stage1_23[37],stage1_22[41],stage1_21[66],stage1_20[103]}
   );
   gpc606_5 gpc424 (
      {stage0_20[155], stage0_20[156], stage0_20[157], stage0_20[158], stage0_20[159], stage0_20[160]},
      {stage0_22[117], stage0_22[118], stage0_22[119], stage0_22[120], stage0_22[121], stage0_22[122]},
      {stage1_24[24],stage1_23[38],stage1_22[42],stage1_21[67],stage1_20[104]}
   );
   gpc606_5 gpc425 (
      {stage0_20[161], stage0_20[162], stage0_20[163], stage0_20[164], stage0_20[165], stage0_20[166]},
      {stage0_22[123], stage0_22[124], stage0_22[125], stage0_22[126], stage0_22[127], stage0_22[128]},
      {stage1_24[25],stage1_23[39],stage1_22[43],stage1_21[68],stage1_20[105]}
   );
   gpc606_5 gpc426 (
      {stage0_20[167], stage0_20[168], stage0_20[169], stage0_20[170], stage0_20[171], stage0_20[172]},
      {stage0_22[129], stage0_22[130], stage0_22[131], stage0_22[132], stage0_22[133], stage0_22[134]},
      {stage1_24[26],stage1_23[40],stage1_22[44],stage1_21[69],stage1_20[106]}
   );
   gpc606_5 gpc427 (
      {stage0_20[173], stage0_20[174], stage0_20[175], stage0_20[176], stage0_20[177], stage0_20[178]},
      {stage0_22[135], stage0_22[136], stage0_22[137], stage0_22[138], stage0_22[139], stage0_22[140]},
      {stage1_24[27],stage1_23[41],stage1_22[45],stage1_21[70],stage1_20[107]}
   );
   gpc606_5 gpc428 (
      {stage0_20[179], stage0_20[180], stage0_20[181], stage0_20[182], stage0_20[183], stage0_20[184]},
      {stage0_22[141], stage0_22[142], stage0_22[143], stage0_22[144], stage0_22[145], stage0_22[146]},
      {stage1_24[28],stage1_23[42],stage1_22[46],stage1_21[71],stage1_20[108]}
   );
   gpc606_5 gpc429 (
      {stage0_20[185], stage0_20[186], stage0_20[187], stage0_20[188], stage0_20[189], stage0_20[190]},
      {stage0_22[147], stage0_22[148], stage0_22[149], stage0_22[150], stage0_22[151], stage0_22[152]},
      {stage1_24[29],stage1_23[43],stage1_22[47],stage1_21[72],stage1_20[109]}
   );
   gpc606_5 gpc430 (
      {stage0_20[191], stage0_20[192], stage0_20[193], stage0_20[194], stage0_20[195], stage0_20[196]},
      {stage0_22[153], stage0_22[154], stage0_22[155], stage0_22[156], stage0_22[157], stage0_22[158]},
      {stage1_24[30],stage1_23[44],stage1_22[48],stage1_21[73],stage1_20[110]}
   );
   gpc606_5 gpc431 (
      {stage0_20[197], stage0_20[198], stage0_20[199], stage0_20[200], stage0_20[201], stage0_20[202]},
      {stage0_22[159], stage0_22[160], stage0_22[161], stage0_22[162], stage0_22[163], stage0_22[164]},
      {stage1_24[31],stage1_23[45],stage1_22[49],stage1_21[74],stage1_20[111]}
   );
   gpc606_5 gpc432 (
      {stage0_20[203], stage0_20[204], stage0_20[205], stage0_20[206], stage0_20[207], stage0_20[208]},
      {stage0_22[165], stage0_22[166], stage0_22[167], stage0_22[168], stage0_22[169], stage0_22[170]},
      {stage1_24[32],stage1_23[46],stage1_22[50],stage1_21[75],stage1_20[112]}
   );
   gpc606_5 gpc433 (
      {stage0_20[209], stage0_20[210], stage0_20[211], stage0_20[212], stage0_20[213], stage0_20[214]},
      {stage0_22[171], stage0_22[172], stage0_22[173], stage0_22[174], stage0_22[175], stage0_22[176]},
      {stage1_24[33],stage1_23[47],stage1_22[51],stage1_21[76],stage1_20[113]}
   );
   gpc606_5 gpc434 (
      {stage0_20[215], stage0_20[216], stage0_20[217], stage0_20[218], stage0_20[219], stage0_20[220]},
      {stage0_22[177], stage0_22[178], stage0_22[179], stage0_22[180], stage0_22[181], stage0_22[182]},
      {stage1_24[34],stage1_23[48],stage1_22[52],stage1_21[77],stage1_20[114]}
   );
   gpc606_5 gpc435 (
      {stage0_20[221], stage0_20[222], stage0_20[223], stage0_20[224], stage0_20[225], stage0_20[226]},
      {stage0_22[183], stage0_22[184], stage0_22[185], stage0_22[186], stage0_22[187], stage0_22[188]},
      {stage1_24[35],stage1_23[49],stage1_22[53],stage1_21[78],stage1_20[115]}
   );
   gpc606_5 gpc436 (
      {stage0_20[227], stage0_20[228], stage0_20[229], stage0_20[230], stage0_20[231], stage0_20[232]},
      {stage0_22[189], stage0_22[190], stage0_22[191], stage0_22[192], stage0_22[193], stage0_22[194]},
      {stage1_24[36],stage1_23[50],stage1_22[54],stage1_21[79],stage1_20[116]}
   );
   gpc606_5 gpc437 (
      {stage0_20[233], stage0_20[234], stage0_20[235], stage0_20[236], stage0_20[237], stage0_20[238]},
      {stage0_22[195], stage0_22[196], stage0_22[197], stage0_22[198], stage0_22[199], stage0_22[200]},
      {stage1_24[37],stage1_23[51],stage1_22[55],stage1_21[80],stage1_20[117]}
   );
   gpc606_5 gpc438 (
      {stage0_20[239], stage0_20[240], stage0_20[241], stage0_20[242], stage0_20[243], stage0_20[244]},
      {stage0_22[201], stage0_22[202], stage0_22[203], stage0_22[204], stage0_22[205], stage0_22[206]},
      {stage1_24[38],stage1_23[52],stage1_22[56],stage1_21[81],stage1_20[118]}
   );
   gpc606_5 gpc439 (
      {stage0_21[120], stage0_21[121], stage0_21[122], stage0_21[123], stage0_21[124], stage0_21[125]},
      {stage0_23[9], stage0_23[10], stage0_23[11], stage0_23[12], stage0_23[13], stage0_23[14]},
      {stage1_25[0],stage1_24[39],stage1_23[53],stage1_22[57],stage1_21[82]}
   );
   gpc606_5 gpc440 (
      {stage0_21[126], stage0_21[127], stage0_21[128], stage0_21[129], stage0_21[130], stage0_21[131]},
      {stage0_23[15], stage0_23[16], stage0_23[17], stage0_23[18], stage0_23[19], stage0_23[20]},
      {stage1_25[1],stage1_24[40],stage1_23[54],stage1_22[58],stage1_21[83]}
   );
   gpc606_5 gpc441 (
      {stage0_21[132], stage0_21[133], stage0_21[134], stage0_21[135], stage0_21[136], stage0_21[137]},
      {stage0_23[21], stage0_23[22], stage0_23[23], stage0_23[24], stage0_23[25], stage0_23[26]},
      {stage1_25[2],stage1_24[41],stage1_23[55],stage1_22[59],stage1_21[84]}
   );
   gpc606_5 gpc442 (
      {stage0_21[138], stage0_21[139], stage0_21[140], stage0_21[141], stage0_21[142], stage0_21[143]},
      {stage0_23[27], stage0_23[28], stage0_23[29], stage0_23[30], stage0_23[31], stage0_23[32]},
      {stage1_25[3],stage1_24[42],stage1_23[56],stage1_22[60],stage1_21[85]}
   );
   gpc606_5 gpc443 (
      {stage0_21[144], stage0_21[145], stage0_21[146], stage0_21[147], stage0_21[148], stage0_21[149]},
      {stage0_23[33], stage0_23[34], stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38]},
      {stage1_25[4],stage1_24[43],stage1_23[57],stage1_22[61],stage1_21[86]}
   );
   gpc606_5 gpc444 (
      {stage0_21[150], stage0_21[151], stage0_21[152], stage0_21[153], stage0_21[154], stage0_21[155]},
      {stage0_23[39], stage0_23[40], stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44]},
      {stage1_25[5],stage1_24[44],stage1_23[58],stage1_22[62],stage1_21[87]}
   );
   gpc606_5 gpc445 (
      {stage0_21[156], stage0_21[157], stage0_21[158], stage0_21[159], stage0_21[160], stage0_21[161]},
      {stage0_23[45], stage0_23[46], stage0_23[47], stage0_23[48], stage0_23[49], stage0_23[50]},
      {stage1_25[6],stage1_24[45],stage1_23[59],stage1_22[63],stage1_21[88]}
   );
   gpc606_5 gpc446 (
      {stage0_21[162], stage0_21[163], stage0_21[164], stage0_21[165], stage0_21[166], stage0_21[167]},
      {stage0_23[51], stage0_23[52], stage0_23[53], stage0_23[54], stage0_23[55], stage0_23[56]},
      {stage1_25[7],stage1_24[46],stage1_23[60],stage1_22[64],stage1_21[89]}
   );
   gpc606_5 gpc447 (
      {stage0_21[168], stage0_21[169], stage0_21[170], stage0_21[171], stage0_21[172], stage0_21[173]},
      {stage0_23[57], stage0_23[58], stage0_23[59], stage0_23[60], stage0_23[61], stage0_23[62]},
      {stage1_25[8],stage1_24[47],stage1_23[61],stage1_22[65],stage1_21[90]}
   );
   gpc606_5 gpc448 (
      {stage0_21[174], stage0_21[175], stage0_21[176], stage0_21[177], stage0_21[178], stage0_21[179]},
      {stage0_23[63], stage0_23[64], stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68]},
      {stage1_25[9],stage1_24[48],stage1_23[62],stage1_22[66],stage1_21[91]}
   );
   gpc606_5 gpc449 (
      {stage0_21[180], stage0_21[181], stage0_21[182], stage0_21[183], stage0_21[184], stage0_21[185]},
      {stage0_23[69], stage0_23[70], stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74]},
      {stage1_25[10],stage1_24[49],stage1_23[63],stage1_22[67],stage1_21[92]}
   );
   gpc606_5 gpc450 (
      {stage0_21[186], stage0_21[187], stage0_21[188], stage0_21[189], stage0_21[190], stage0_21[191]},
      {stage0_23[75], stage0_23[76], stage0_23[77], stage0_23[78], stage0_23[79], stage0_23[80]},
      {stage1_25[11],stage1_24[50],stage1_23[64],stage1_22[68],stage1_21[93]}
   );
   gpc606_5 gpc451 (
      {stage0_21[192], stage0_21[193], stage0_21[194], stage0_21[195], stage0_21[196], stage0_21[197]},
      {stage0_23[81], stage0_23[82], stage0_23[83], stage0_23[84], stage0_23[85], stage0_23[86]},
      {stage1_25[12],stage1_24[51],stage1_23[65],stage1_22[69],stage1_21[94]}
   );
   gpc606_5 gpc452 (
      {stage0_21[198], stage0_21[199], stage0_21[200], stage0_21[201], stage0_21[202], stage0_21[203]},
      {stage0_23[87], stage0_23[88], stage0_23[89], stage0_23[90], stage0_23[91], stage0_23[92]},
      {stage1_25[13],stage1_24[52],stage1_23[66],stage1_22[70],stage1_21[95]}
   );
   gpc606_5 gpc453 (
      {stage0_21[204], stage0_21[205], stage0_21[206], stage0_21[207], stage0_21[208], stage0_21[209]},
      {stage0_23[93], stage0_23[94], stage0_23[95], stage0_23[96], stage0_23[97], stage0_23[98]},
      {stage1_25[14],stage1_24[53],stage1_23[67],stage1_22[71],stage1_21[96]}
   );
   gpc606_5 gpc454 (
      {stage0_21[210], stage0_21[211], stage0_21[212], stage0_21[213], stage0_21[214], stage0_21[215]},
      {stage0_23[99], stage0_23[100], stage0_23[101], stage0_23[102], stage0_23[103], stage0_23[104]},
      {stage1_25[15],stage1_24[54],stage1_23[68],stage1_22[72],stage1_21[97]}
   );
   gpc606_5 gpc455 (
      {stage0_21[216], stage0_21[217], stage0_21[218], stage0_21[219], stage0_21[220], stage0_21[221]},
      {stage0_23[105], stage0_23[106], stage0_23[107], stage0_23[108], stage0_23[109], stage0_23[110]},
      {stage1_25[16],stage1_24[55],stage1_23[69],stage1_22[73],stage1_21[98]}
   );
   gpc606_5 gpc456 (
      {stage0_21[222], stage0_21[223], stage0_21[224], stage0_21[225], stage0_21[226], stage0_21[227]},
      {stage0_23[111], stage0_23[112], stage0_23[113], stage0_23[114], stage0_23[115], stage0_23[116]},
      {stage1_25[17],stage1_24[56],stage1_23[70],stage1_22[74],stage1_21[99]}
   );
   gpc606_5 gpc457 (
      {stage0_21[228], stage0_21[229], stage0_21[230], stage0_21[231], stage0_21[232], stage0_21[233]},
      {stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120], stage0_23[121], stage0_23[122]},
      {stage1_25[18],stage1_24[57],stage1_23[71],stage1_22[75],stage1_21[100]}
   );
   gpc606_5 gpc458 (
      {stage0_21[234], stage0_21[235], stage0_21[236], stage0_21[237], stage0_21[238], stage0_21[239]},
      {stage0_23[123], stage0_23[124], stage0_23[125], stage0_23[126], stage0_23[127], stage0_23[128]},
      {stage1_25[19],stage1_24[58],stage1_23[72],stage1_22[76],stage1_21[101]}
   );
   gpc606_5 gpc459 (
      {stage0_21[240], stage0_21[241], stage0_21[242], stage0_21[243], stage0_21[244], stage0_21[245]},
      {stage0_23[129], stage0_23[130], stage0_23[131], stage0_23[132], stage0_23[133], stage0_23[134]},
      {stage1_25[20],stage1_24[59],stage1_23[73],stage1_22[77],stage1_21[102]}
   );
   gpc606_5 gpc460 (
      {stage0_21[246], stage0_21[247], stage0_21[248], stage0_21[249], stage0_21[250], stage0_21[251]},
      {stage0_23[135], stage0_23[136], stage0_23[137], stage0_23[138], stage0_23[139], stage0_23[140]},
      {stage1_25[21],stage1_24[60],stage1_23[74],stage1_22[78],stage1_21[103]}
   );
   gpc615_5 gpc461 (
      {stage0_22[207], stage0_22[208], stage0_22[209], stage0_22[210], stage0_22[211]},
      {stage0_23[141]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[22],stage1_24[61],stage1_23[75],stage1_22[79]}
   );
   gpc615_5 gpc462 (
      {stage0_22[212], stage0_22[213], stage0_22[214], stage0_22[215], stage0_22[216]},
      {stage0_23[142]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[23],stage1_24[62],stage1_23[76],stage1_22[80]}
   );
   gpc615_5 gpc463 (
      {stage0_22[217], stage0_22[218], stage0_22[219], stage0_22[220], stage0_22[221]},
      {stage0_23[143]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[24],stage1_24[63],stage1_23[77],stage1_22[81]}
   );
   gpc615_5 gpc464 (
      {stage0_22[222], stage0_22[223], stage0_22[224], stage0_22[225], stage0_22[226]},
      {stage0_23[144]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[25],stage1_24[64],stage1_23[78],stage1_22[82]}
   );
   gpc615_5 gpc465 (
      {stage0_22[227], stage0_22[228], stage0_22[229], stage0_22[230], stage0_22[231]},
      {stage0_23[145]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[26],stage1_24[65],stage1_23[79],stage1_22[83]}
   );
   gpc615_5 gpc466 (
      {stage0_22[232], stage0_22[233], stage0_22[234], stage0_22[235], stage0_22[236]},
      {stage0_23[146]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[27],stage1_24[66],stage1_23[80],stage1_22[84]}
   );
   gpc615_5 gpc467 (
      {stage0_22[237], stage0_22[238], stage0_22[239], stage0_22[240], stage0_22[241]},
      {stage0_23[147]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[28],stage1_24[67],stage1_23[81],stage1_22[85]}
   );
   gpc615_5 gpc468 (
      {stage0_22[242], stage0_22[243], stage0_22[244], stage0_22[245], stage0_22[246]},
      {stage0_23[148]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[29],stage1_24[68],stage1_23[82],stage1_22[86]}
   );
   gpc615_5 gpc469 (
      {stage0_22[247], stage0_22[248], stage0_22[249], stage0_22[250], stage0_22[251]},
      {stage0_23[149]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[30],stage1_24[69],stage1_23[83],stage1_22[87]}
   );
   gpc606_5 gpc470 (
      {stage0_23[150], stage0_23[151], stage0_23[152], stage0_23[153], stage0_23[154], stage0_23[155]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[9],stage1_25[31],stage1_24[70],stage1_23[84]}
   );
   gpc615_5 gpc471 (
      {stage0_23[156], stage0_23[157], stage0_23[158], stage0_23[159], stage0_23[160]},
      {stage0_24[54]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[10],stage1_25[32],stage1_24[71],stage1_23[85]}
   );
   gpc615_5 gpc472 (
      {stage0_23[161], stage0_23[162], stage0_23[163], stage0_23[164], stage0_23[165]},
      {stage0_24[55]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[11],stage1_25[33],stage1_24[72],stage1_23[86]}
   );
   gpc615_5 gpc473 (
      {stage0_23[166], stage0_23[167], stage0_23[168], stage0_23[169], stage0_23[170]},
      {stage0_24[56]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[12],stage1_25[34],stage1_24[73],stage1_23[87]}
   );
   gpc615_5 gpc474 (
      {stage0_23[171], stage0_23[172], stage0_23[173], stage0_23[174], stage0_23[175]},
      {stage0_24[57]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[13],stage1_25[35],stage1_24[74],stage1_23[88]}
   );
   gpc615_5 gpc475 (
      {stage0_23[176], stage0_23[177], stage0_23[178], stage0_23[179], stage0_23[180]},
      {stage0_24[58]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[14],stage1_25[36],stage1_24[75],stage1_23[89]}
   );
   gpc615_5 gpc476 (
      {stage0_23[181], stage0_23[182], stage0_23[183], stage0_23[184], stage0_23[185]},
      {stage0_24[59]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[15],stage1_25[37],stage1_24[76],stage1_23[90]}
   );
   gpc615_5 gpc477 (
      {stage0_23[186], stage0_23[187], stage0_23[188], stage0_23[189], stage0_23[190]},
      {stage0_24[60]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[16],stage1_25[38],stage1_24[77],stage1_23[91]}
   );
   gpc615_5 gpc478 (
      {stage0_23[191], stage0_23[192], stage0_23[193], stage0_23[194], stage0_23[195]},
      {stage0_24[61]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[17],stage1_25[39],stage1_24[78],stage1_23[92]}
   );
   gpc615_5 gpc479 (
      {stage0_23[196], stage0_23[197], stage0_23[198], stage0_23[199], stage0_23[200]},
      {stage0_24[62]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[18],stage1_25[40],stage1_24[79],stage1_23[93]}
   );
   gpc615_5 gpc480 (
      {stage0_23[201], stage0_23[202], stage0_23[203], stage0_23[204], stage0_23[205]},
      {stage0_24[63]},
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage1_27[10],stage1_26[19],stage1_25[41],stage1_24[80],stage1_23[94]}
   );
   gpc615_5 gpc481 (
      {stage0_23[206], stage0_23[207], stage0_23[208], stage0_23[209], stage0_23[210]},
      {stage0_24[64]},
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage1_27[11],stage1_26[20],stage1_25[42],stage1_24[81],stage1_23[95]}
   );
   gpc615_5 gpc482 (
      {stage0_23[211], stage0_23[212], stage0_23[213], stage0_23[214], stage0_23[215]},
      {stage0_24[65]},
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage1_27[12],stage1_26[21],stage1_25[43],stage1_24[82],stage1_23[96]}
   );
   gpc615_5 gpc483 (
      {stage0_23[216], stage0_23[217], stage0_23[218], stage0_23[219], stage0_23[220]},
      {stage0_24[66]},
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage1_27[13],stage1_26[22],stage1_25[44],stage1_24[83],stage1_23[97]}
   );
   gpc615_5 gpc484 (
      {stage0_23[221], stage0_23[222], stage0_23[223], stage0_23[224], stage0_23[225]},
      {stage0_24[67]},
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage1_27[14],stage1_26[23],stage1_25[45],stage1_24[84],stage1_23[98]}
   );
   gpc606_5 gpc485 (
      {stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71], stage0_24[72], stage0_24[73]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[15],stage1_26[24],stage1_25[46],stage1_24[85]}
   );
   gpc606_5 gpc486 (
      {stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77], stage0_24[78], stage0_24[79]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[16],stage1_26[25],stage1_25[47],stage1_24[86]}
   );
   gpc606_5 gpc487 (
      {stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83], stage0_24[84], stage0_24[85]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[17],stage1_26[26],stage1_25[48],stage1_24[87]}
   );
   gpc606_5 gpc488 (
      {stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89], stage0_24[90], stage0_24[91]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[18],stage1_26[27],stage1_25[49],stage1_24[88]}
   );
   gpc606_5 gpc489 (
      {stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95], stage0_24[96], stage0_24[97]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[19],stage1_26[28],stage1_25[50],stage1_24[89]}
   );
   gpc606_5 gpc490 (
      {stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101], stage0_24[102], stage0_24[103]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[20],stage1_26[29],stage1_25[51],stage1_24[90]}
   );
   gpc606_5 gpc491 (
      {stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107], stage0_24[108], stage0_24[109]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[21],stage1_26[30],stage1_25[52],stage1_24[91]}
   );
   gpc606_5 gpc492 (
      {stage0_24[110], stage0_24[111], stage0_24[112], stage0_24[113], stage0_24[114], stage0_24[115]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[22],stage1_26[31],stage1_25[53],stage1_24[92]}
   );
   gpc606_5 gpc493 (
      {stage0_24[116], stage0_24[117], stage0_24[118], stage0_24[119], stage0_24[120], stage0_24[121]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[23],stage1_26[32],stage1_25[54],stage1_24[93]}
   );
   gpc606_5 gpc494 (
      {stage0_24[122], stage0_24[123], stage0_24[124], stage0_24[125], stage0_24[126], stage0_24[127]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[24],stage1_26[33],stage1_25[55],stage1_24[94]}
   );
   gpc606_5 gpc495 (
      {stage0_24[128], stage0_24[129], stage0_24[130], stage0_24[131], stage0_24[132], stage0_24[133]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[25],stage1_26[34],stage1_25[56],stage1_24[95]}
   );
   gpc606_5 gpc496 (
      {stage0_24[134], stage0_24[135], stage0_24[136], stage0_24[137], stage0_24[138], stage0_24[139]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[26],stage1_26[35],stage1_25[57],stage1_24[96]}
   );
   gpc606_5 gpc497 (
      {stage0_24[140], stage0_24[141], stage0_24[142], stage0_24[143], stage0_24[144], stage0_24[145]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[27],stage1_26[36],stage1_25[58],stage1_24[97]}
   );
   gpc615_5 gpc498 (
      {stage0_24[146], stage0_24[147], stage0_24[148], stage0_24[149], stage0_24[150]},
      {stage0_25[90]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[28],stage1_26[37],stage1_25[59],stage1_24[98]}
   );
   gpc615_5 gpc499 (
      {stage0_24[151], stage0_24[152], stage0_24[153], stage0_24[154], stage0_24[155]},
      {stage0_25[91]},
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88], stage0_26[89]},
      {stage1_28[14],stage1_27[29],stage1_26[38],stage1_25[60],stage1_24[99]}
   );
   gpc615_5 gpc500 (
      {stage0_24[156], stage0_24[157], stage0_24[158], stage0_24[159], stage0_24[160]},
      {stage0_25[92]},
      {stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93], stage0_26[94], stage0_26[95]},
      {stage1_28[15],stage1_27[30],stage1_26[39],stage1_25[61],stage1_24[100]}
   );
   gpc615_5 gpc501 (
      {stage0_24[161], stage0_24[162], stage0_24[163], stage0_24[164], stage0_24[165]},
      {stage0_25[93]},
      {stage0_26[96], stage0_26[97], stage0_26[98], stage0_26[99], stage0_26[100], stage0_26[101]},
      {stage1_28[16],stage1_27[31],stage1_26[40],stage1_25[62],stage1_24[101]}
   );
   gpc615_5 gpc502 (
      {stage0_24[166], stage0_24[167], stage0_24[168], stage0_24[169], stage0_24[170]},
      {stage0_25[94]},
      {stage0_26[102], stage0_26[103], stage0_26[104], stage0_26[105], stage0_26[106], stage0_26[107]},
      {stage1_28[17],stage1_27[32],stage1_26[41],stage1_25[63],stage1_24[102]}
   );
   gpc615_5 gpc503 (
      {stage0_24[171], stage0_24[172], stage0_24[173], stage0_24[174], stage0_24[175]},
      {stage0_25[95]},
      {stage0_26[108], stage0_26[109], stage0_26[110], stage0_26[111], stage0_26[112], stage0_26[113]},
      {stage1_28[18],stage1_27[33],stage1_26[42],stage1_25[64],stage1_24[103]}
   );
   gpc615_5 gpc504 (
      {stage0_24[176], stage0_24[177], stage0_24[178], stage0_24[179], stage0_24[180]},
      {stage0_25[96]},
      {stage0_26[114], stage0_26[115], stage0_26[116], stage0_26[117], stage0_26[118], stage0_26[119]},
      {stage1_28[19],stage1_27[34],stage1_26[43],stage1_25[65],stage1_24[104]}
   );
   gpc615_5 gpc505 (
      {stage0_24[181], stage0_24[182], stage0_24[183], stage0_24[184], stage0_24[185]},
      {stage0_25[97]},
      {stage0_26[120], stage0_26[121], stage0_26[122], stage0_26[123], stage0_26[124], stage0_26[125]},
      {stage1_28[20],stage1_27[35],stage1_26[44],stage1_25[66],stage1_24[105]}
   );
   gpc615_5 gpc506 (
      {stage0_24[186], stage0_24[187], stage0_24[188], stage0_24[189], stage0_24[190]},
      {stage0_25[98]},
      {stage0_26[126], stage0_26[127], stage0_26[128], stage0_26[129], stage0_26[130], stage0_26[131]},
      {stage1_28[21],stage1_27[36],stage1_26[45],stage1_25[67],stage1_24[106]}
   );
   gpc615_5 gpc507 (
      {stage0_24[191], stage0_24[192], stage0_24[193], stage0_24[194], stage0_24[195]},
      {stage0_25[99]},
      {stage0_26[132], stage0_26[133], stage0_26[134], stage0_26[135], stage0_26[136], stage0_26[137]},
      {stage1_28[22],stage1_27[37],stage1_26[46],stage1_25[68],stage1_24[107]}
   );
   gpc615_5 gpc508 (
      {stage0_24[196], stage0_24[197], stage0_24[198], stage0_24[199], stage0_24[200]},
      {stage0_25[100]},
      {stage0_26[138], stage0_26[139], stage0_26[140], stage0_26[141], stage0_26[142], stage0_26[143]},
      {stage1_28[23],stage1_27[38],stage1_26[47],stage1_25[69],stage1_24[108]}
   );
   gpc615_5 gpc509 (
      {stage0_24[201], stage0_24[202], stage0_24[203], stage0_24[204], stage0_24[205]},
      {stage0_25[101]},
      {stage0_26[144], stage0_26[145], stage0_26[146], stage0_26[147], stage0_26[148], stage0_26[149]},
      {stage1_28[24],stage1_27[39],stage1_26[48],stage1_25[70],stage1_24[109]}
   );
   gpc615_5 gpc510 (
      {stage0_24[206], stage0_24[207], stage0_24[208], stage0_24[209], stage0_24[210]},
      {stage0_25[102]},
      {stage0_26[150], stage0_26[151], stage0_26[152], stage0_26[153], stage0_26[154], stage0_26[155]},
      {stage1_28[25],stage1_27[40],stage1_26[49],stage1_25[71],stage1_24[110]}
   );
   gpc615_5 gpc511 (
      {stage0_24[211], stage0_24[212], stage0_24[213], stage0_24[214], stage0_24[215]},
      {stage0_25[103]},
      {stage0_26[156], stage0_26[157], stage0_26[158], stage0_26[159], stage0_26[160], stage0_26[161]},
      {stage1_28[26],stage1_27[41],stage1_26[50],stage1_25[72],stage1_24[111]}
   );
   gpc615_5 gpc512 (
      {stage0_24[216], stage0_24[217], stage0_24[218], stage0_24[219], stage0_24[220]},
      {stage0_25[104]},
      {stage0_26[162], stage0_26[163], stage0_26[164], stage0_26[165], stage0_26[166], stage0_26[167]},
      {stage1_28[27],stage1_27[42],stage1_26[51],stage1_25[73],stage1_24[112]}
   );
   gpc615_5 gpc513 (
      {stage0_24[221], stage0_24[222], stage0_24[223], stage0_24[224], stage0_24[225]},
      {stage0_25[105]},
      {stage0_26[168], stage0_26[169], stage0_26[170], stage0_26[171], stage0_26[172], stage0_26[173]},
      {stage1_28[28],stage1_27[43],stage1_26[52],stage1_25[74],stage1_24[113]}
   );
   gpc615_5 gpc514 (
      {stage0_24[226], stage0_24[227], stage0_24[228], stage0_24[229], stage0_24[230]},
      {stage0_25[106]},
      {stage0_26[174], stage0_26[175], stage0_26[176], stage0_26[177], stage0_26[178], stage0_26[179]},
      {stage1_28[29],stage1_27[44],stage1_26[53],stage1_25[75],stage1_24[114]}
   );
   gpc606_5 gpc515 (
      {stage0_25[107], stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[30],stage1_27[45],stage1_26[54],stage1_25[76]}
   );
   gpc606_5 gpc516 (
      {stage0_25[113], stage0_25[114], stage0_25[115], stage0_25[116], stage0_25[117], stage0_25[118]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[31],stage1_27[46],stage1_26[55],stage1_25[77]}
   );
   gpc606_5 gpc517 (
      {stage0_25[119], stage0_25[120], stage0_25[121], stage0_25[122], stage0_25[123], stage0_25[124]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[32],stage1_27[47],stage1_26[56],stage1_25[78]}
   );
   gpc606_5 gpc518 (
      {stage0_25[125], stage0_25[126], stage0_25[127], stage0_25[128], stage0_25[129], stage0_25[130]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[33],stage1_27[48],stage1_26[57],stage1_25[79]}
   );
   gpc606_5 gpc519 (
      {stage0_25[131], stage0_25[132], stage0_25[133], stage0_25[134], stage0_25[135], stage0_25[136]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[34],stage1_27[49],stage1_26[58],stage1_25[80]}
   );
   gpc606_5 gpc520 (
      {stage0_25[137], stage0_25[138], stage0_25[139], stage0_25[140], stage0_25[141], stage0_25[142]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[35],stage1_27[50],stage1_26[59],stage1_25[81]}
   );
   gpc606_5 gpc521 (
      {stage0_25[143], stage0_25[144], stage0_25[145], stage0_25[146], stage0_25[147], stage0_25[148]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[36],stage1_27[51],stage1_26[60],stage1_25[82]}
   );
   gpc606_5 gpc522 (
      {stage0_25[149], stage0_25[150], stage0_25[151], stage0_25[152], stage0_25[153], stage0_25[154]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[37],stage1_27[52],stage1_26[61],stage1_25[83]}
   );
   gpc606_5 gpc523 (
      {stage0_25[155], stage0_25[156], stage0_25[157], stage0_25[158], stage0_25[159], stage0_25[160]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[38],stage1_27[53],stage1_26[62],stage1_25[84]}
   );
   gpc606_5 gpc524 (
      {stage0_25[161], stage0_25[162], stage0_25[163], stage0_25[164], stage0_25[165], stage0_25[166]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[39],stage1_27[54],stage1_26[63],stage1_25[85]}
   );
   gpc606_5 gpc525 (
      {stage0_25[167], stage0_25[168], stage0_25[169], stage0_25[170], stage0_25[171], stage0_25[172]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[40],stage1_27[55],stage1_26[64],stage1_25[86]}
   );
   gpc606_5 gpc526 (
      {stage0_25[173], stage0_25[174], stage0_25[175], stage0_25[176], stage0_25[177], stage0_25[178]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[41],stage1_27[56],stage1_26[65],stage1_25[87]}
   );
   gpc606_5 gpc527 (
      {stage0_25[179], stage0_25[180], stage0_25[181], stage0_25[182], stage0_25[183], stage0_25[184]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[42],stage1_27[57],stage1_26[66],stage1_25[88]}
   );
   gpc606_5 gpc528 (
      {stage0_25[185], stage0_25[186], stage0_25[187], stage0_25[188], stage0_25[189], stage0_25[190]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[43],stage1_27[58],stage1_26[67],stage1_25[89]}
   );
   gpc606_5 gpc529 (
      {stage0_25[191], stage0_25[192], stage0_25[193], stage0_25[194], stage0_25[195], stage0_25[196]},
      {stage0_27[84], stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage1_29[14],stage1_28[44],stage1_27[59],stage1_26[68],stage1_25[90]}
   );
   gpc606_5 gpc530 (
      {stage0_25[197], stage0_25[198], stage0_25[199], stage0_25[200], stage0_25[201], stage0_25[202]},
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage1_29[15],stage1_28[45],stage1_27[60],stage1_26[69],stage1_25[91]}
   );
   gpc606_5 gpc531 (
      {stage0_25[203], stage0_25[204], stage0_25[205], stage0_25[206], stage0_25[207], stage0_25[208]},
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage1_29[16],stage1_28[46],stage1_27[61],stage1_26[70],stage1_25[92]}
   );
   gpc606_5 gpc532 (
      {stage0_25[209], stage0_25[210], stage0_25[211], stage0_25[212], stage0_25[213], stage0_25[214]},
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage1_29[17],stage1_28[47],stage1_27[62],stage1_26[71],stage1_25[93]}
   );
   gpc606_5 gpc533 (
      {stage0_25[215], stage0_25[216], stage0_25[217], stage0_25[218], stage0_25[219], stage0_25[220]},
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage1_29[18],stage1_28[48],stage1_27[63],stage1_26[72],stage1_25[94]}
   );
   gpc606_5 gpc534 (
      {stage0_25[221], stage0_25[222], stage0_25[223], stage0_25[224], stage0_25[225], stage0_25[226]},
      {stage0_27[114], stage0_27[115], stage0_27[116], stage0_27[117], stage0_27[118], stage0_27[119]},
      {stage1_29[19],stage1_28[49],stage1_27[64],stage1_26[73],stage1_25[95]}
   );
   gpc606_5 gpc535 (
      {stage0_25[227], stage0_25[228], stage0_25[229], stage0_25[230], stage0_25[231], stage0_25[232]},
      {stage0_27[120], stage0_27[121], stage0_27[122], stage0_27[123], stage0_27[124], stage0_27[125]},
      {stage1_29[20],stage1_28[50],stage1_27[65],stage1_26[74],stage1_25[96]}
   );
   gpc606_5 gpc536 (
      {stage0_25[233], stage0_25[234], stage0_25[235], stage0_25[236], stage0_25[237], stage0_25[238]},
      {stage0_27[126], stage0_27[127], stage0_27[128], stage0_27[129], stage0_27[130], stage0_27[131]},
      {stage1_29[21],stage1_28[51],stage1_27[66],stage1_26[75],stage1_25[97]}
   );
   gpc606_5 gpc537 (
      {stage0_25[239], stage0_25[240], stage0_25[241], stage0_25[242], stage0_25[243], stage0_25[244]},
      {stage0_27[132], stage0_27[133], stage0_27[134], stage0_27[135], stage0_27[136], stage0_27[137]},
      {stage1_29[22],stage1_28[52],stage1_27[67],stage1_26[76],stage1_25[98]}
   );
   gpc615_5 gpc538 (
      {stage0_26[180], stage0_26[181], stage0_26[182], stage0_26[183], stage0_26[184]},
      {stage0_27[138]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[23],stage1_28[53],stage1_27[68],stage1_26[77]}
   );
   gpc615_5 gpc539 (
      {stage0_26[185], stage0_26[186], stage0_26[187], stage0_26[188], stage0_26[189]},
      {stage0_27[139]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[24],stage1_28[54],stage1_27[69],stage1_26[78]}
   );
   gpc615_5 gpc540 (
      {stage0_26[190], stage0_26[191], stage0_26[192], stage0_26[193], stage0_26[194]},
      {stage0_27[140]},
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage1_30[2],stage1_29[25],stage1_28[55],stage1_27[70],stage1_26[79]}
   );
   gpc606_5 gpc541 (
      {stage0_27[141], stage0_27[142], stage0_27[143], stage0_27[144], stage0_27[145], stage0_27[146]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[3],stage1_29[26],stage1_28[56],stage1_27[71]}
   );
   gpc606_5 gpc542 (
      {stage0_27[147], stage0_27[148], stage0_27[149], stage0_27[150], stage0_27[151], stage0_27[152]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[4],stage1_29[27],stage1_28[57],stage1_27[72]}
   );
   gpc606_5 gpc543 (
      {stage0_27[153], stage0_27[154], stage0_27[155], stage0_27[156], stage0_27[157], stage0_27[158]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[5],stage1_29[28],stage1_28[58],stage1_27[73]}
   );
   gpc615_5 gpc544 (
      {stage0_27[159], stage0_27[160], stage0_27[161], stage0_27[162], stage0_27[163]},
      {stage0_28[18]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[6],stage1_29[29],stage1_28[59],stage1_27[74]}
   );
   gpc615_5 gpc545 (
      {stage0_27[164], stage0_27[165], stage0_27[166], stage0_27[167], stage0_27[168]},
      {stage0_28[19]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[7],stage1_29[30],stage1_28[60],stage1_27[75]}
   );
   gpc615_5 gpc546 (
      {stage0_27[169], stage0_27[170], stage0_27[171], stage0_27[172], stage0_27[173]},
      {stage0_28[20]},
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage1_31[5],stage1_30[8],stage1_29[31],stage1_28[61],stage1_27[76]}
   );
   gpc615_5 gpc547 (
      {stage0_27[174], stage0_27[175], stage0_27[176], stage0_27[177], stage0_27[178]},
      {stage0_28[21]},
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage1_31[6],stage1_30[9],stage1_29[32],stage1_28[62],stage1_27[77]}
   );
   gpc615_5 gpc548 (
      {stage0_27[179], stage0_27[180], stage0_27[181], stage0_27[182], stage0_27[183]},
      {stage0_28[22]},
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage1_31[7],stage1_30[10],stage1_29[33],stage1_28[63],stage1_27[78]}
   );
   gpc615_5 gpc549 (
      {stage0_27[184], stage0_27[185], stage0_27[186], stage0_27[187], stage0_27[188]},
      {stage0_28[23]},
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage1_31[8],stage1_30[11],stage1_29[34],stage1_28[64],stage1_27[79]}
   );
   gpc615_5 gpc550 (
      {stage0_27[189], stage0_27[190], stage0_27[191], stage0_27[192], stage0_27[193]},
      {stage0_28[24]},
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage1_31[9],stage1_30[12],stage1_29[35],stage1_28[65],stage1_27[80]}
   );
   gpc615_5 gpc551 (
      {stage0_27[194], stage0_27[195], stage0_27[196], stage0_27[197], stage0_27[198]},
      {stage0_28[25]},
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage1_31[10],stage1_30[13],stage1_29[36],stage1_28[66],stage1_27[81]}
   );
   gpc615_5 gpc552 (
      {stage0_27[199], stage0_27[200], stage0_27[201], stage0_27[202], stage0_27[203]},
      {stage0_28[26]},
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage1_31[11],stage1_30[14],stage1_29[37],stage1_28[67],stage1_27[82]}
   );
   gpc615_5 gpc553 (
      {stage0_27[204], stage0_27[205], stage0_27[206], stage0_27[207], stage0_27[208]},
      {stage0_28[27]},
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage1_31[12],stage1_30[15],stage1_29[38],stage1_28[68],stage1_27[83]}
   );
   gpc615_5 gpc554 (
      {stage0_27[209], stage0_27[210], stage0_27[211], stage0_27[212], stage0_27[213]},
      {stage0_28[28]},
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage1_31[13],stage1_30[16],stage1_29[39],stage1_28[69],stage1_27[84]}
   );
   gpc615_5 gpc555 (
      {stage0_27[214], stage0_27[215], stage0_27[216], stage0_27[217], stage0_27[218]},
      {stage0_28[29]},
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage1_31[14],stage1_30[17],stage1_29[40],stage1_28[70],stage1_27[85]}
   );
   gpc615_5 gpc556 (
      {stage0_27[219], stage0_27[220], stage0_27[221], stage0_27[222], stage0_27[223]},
      {stage0_28[30]},
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage1_31[15],stage1_30[18],stage1_29[41],stage1_28[71],stage1_27[86]}
   );
   gpc2116_5 gpc557 (
      {stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35], stage0_28[36]},
      {stage0_29[96]},
      {stage0_30[0]},
      {stage0_31[0], stage0_31[1]},
      {stage1_32[0],stage1_31[16],stage1_30[19],stage1_29[42],stage1_28[72]}
   );
   gpc606_5 gpc558 (
      {stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42]},
      {stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5], stage0_30[6]},
      {stage1_32[1],stage1_31[17],stage1_30[20],stage1_29[43],stage1_28[73]}
   );
   gpc606_5 gpc559 (
      {stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47], stage0_28[48]},
      {stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11], stage0_30[12]},
      {stage1_32[2],stage1_31[18],stage1_30[21],stage1_29[44],stage1_28[74]}
   );
   gpc606_5 gpc560 (
      {stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53], stage0_28[54]},
      {stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17], stage0_30[18]},
      {stage1_32[3],stage1_31[19],stage1_30[22],stage1_29[45],stage1_28[75]}
   );
   gpc606_5 gpc561 (
      {stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58], stage0_28[59], stage0_28[60]},
      {stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23], stage0_30[24]},
      {stage1_32[4],stage1_31[20],stage1_30[23],stage1_29[46],stage1_28[76]}
   );
   gpc606_5 gpc562 (
      {stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64], stage0_28[65], stage0_28[66]},
      {stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29], stage0_30[30]},
      {stage1_32[5],stage1_31[21],stage1_30[24],stage1_29[47],stage1_28[77]}
   );
   gpc606_5 gpc563 (
      {stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70], stage0_28[71], stage0_28[72]},
      {stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35], stage0_30[36]},
      {stage1_32[6],stage1_31[22],stage1_30[25],stage1_29[48],stage1_28[78]}
   );
   gpc606_5 gpc564 (
      {stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76], stage0_28[77], stage0_28[78]},
      {stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41], stage0_30[42]},
      {stage1_32[7],stage1_31[23],stage1_30[26],stage1_29[49],stage1_28[79]}
   );
   gpc606_5 gpc565 (
      {stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82], stage0_28[83], stage0_28[84]},
      {stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47], stage0_30[48]},
      {stage1_32[8],stage1_31[24],stage1_30[27],stage1_29[50],stage1_28[80]}
   );
   gpc606_5 gpc566 (
      {stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88], stage0_28[89], stage0_28[90]},
      {stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53], stage0_30[54]},
      {stage1_32[9],stage1_31[25],stage1_30[28],stage1_29[51],stage1_28[81]}
   );
   gpc606_5 gpc567 (
      {stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94], stage0_28[95], stage0_28[96]},
      {stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60]},
      {stage1_32[10],stage1_31[26],stage1_30[29],stage1_29[52],stage1_28[82]}
   );
   gpc606_5 gpc568 (
      {stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100], stage0_28[101], stage0_28[102]},
      {stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66]},
      {stage1_32[11],stage1_31[27],stage1_30[30],stage1_29[53],stage1_28[83]}
   );
   gpc606_5 gpc569 (
      {stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106], stage0_28[107], stage0_28[108]},
      {stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72]},
      {stage1_32[12],stage1_31[28],stage1_30[31],stage1_29[54],stage1_28[84]}
   );
   gpc606_5 gpc570 (
      {stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114]},
      {stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78]},
      {stage1_32[13],stage1_31[29],stage1_30[32],stage1_29[55],stage1_28[85]}
   );
   gpc606_5 gpc571 (
      {stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83], stage0_30[84]},
      {stage1_32[14],stage1_31[30],stage1_30[33],stage1_29[56],stage1_28[86]}
   );
   gpc606_5 gpc572 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125], stage0_28[126]},
      {stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89], stage0_30[90]},
      {stage1_32[15],stage1_31[31],stage1_30[34],stage1_29[57],stage1_28[87]}
   );
   gpc606_5 gpc573 (
      {stage0_28[127], stage0_28[128], stage0_28[129], stage0_28[130], stage0_28[131], stage0_28[132]},
      {stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95], stage0_30[96]},
      {stage1_32[16],stage1_31[32],stage1_30[35],stage1_29[58],stage1_28[88]}
   );
   gpc606_5 gpc574 (
      {stage0_28[133], stage0_28[134], stage0_28[135], stage0_28[136], stage0_28[137], stage0_28[138]},
      {stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101], stage0_30[102]},
      {stage1_32[17],stage1_31[33],stage1_30[36],stage1_29[59],stage1_28[89]}
   );
   gpc606_5 gpc575 (
      {stage0_28[139], stage0_28[140], stage0_28[141], stage0_28[142], stage0_28[143], stage0_28[144]},
      {stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107], stage0_30[108]},
      {stage1_32[18],stage1_31[34],stage1_30[37],stage1_29[60],stage1_28[90]}
   );
   gpc606_5 gpc576 (
      {stage0_28[145], stage0_28[146], stage0_28[147], stage0_28[148], stage0_28[149], stage0_28[150]},
      {stage0_30[109], stage0_30[110], stage0_30[111], stage0_30[112], stage0_30[113], stage0_30[114]},
      {stage1_32[19],stage1_31[35],stage1_30[38],stage1_29[61],stage1_28[91]}
   );
   gpc606_5 gpc577 (
      {stage0_28[151], stage0_28[152], stage0_28[153], stage0_28[154], stage0_28[155], stage0_28[156]},
      {stage0_30[115], stage0_30[116], stage0_30[117], stage0_30[118], stage0_30[119], stage0_30[120]},
      {stage1_32[20],stage1_31[36],stage1_30[39],stage1_29[62],stage1_28[92]}
   );
   gpc606_5 gpc578 (
      {stage0_28[157], stage0_28[158], stage0_28[159], stage0_28[160], stage0_28[161], stage0_28[162]},
      {stage0_30[121], stage0_30[122], stage0_30[123], stage0_30[124], stage0_30[125], stage0_30[126]},
      {stage1_32[21],stage1_31[37],stage1_30[40],stage1_29[63],stage1_28[93]}
   );
   gpc606_5 gpc579 (
      {stage0_28[163], stage0_28[164], stage0_28[165], stage0_28[166], stage0_28[167], stage0_28[168]},
      {stage0_30[127], stage0_30[128], stage0_30[129], stage0_30[130], stage0_30[131], stage0_30[132]},
      {stage1_32[22],stage1_31[38],stage1_30[41],stage1_29[64],stage1_28[94]}
   );
   gpc606_5 gpc580 (
      {stage0_28[169], stage0_28[170], stage0_28[171], stage0_28[172], stage0_28[173], stage0_28[174]},
      {stage0_30[133], stage0_30[134], stage0_30[135], stage0_30[136], stage0_30[137], stage0_30[138]},
      {stage1_32[23],stage1_31[39],stage1_30[42],stage1_29[65],stage1_28[95]}
   );
   gpc606_5 gpc581 (
      {stage0_28[175], stage0_28[176], stage0_28[177], stage0_28[178], stage0_28[179], stage0_28[180]},
      {stage0_30[139], stage0_30[140], stage0_30[141], stage0_30[142], stage0_30[143], stage0_30[144]},
      {stage1_32[24],stage1_31[40],stage1_30[43],stage1_29[66],stage1_28[96]}
   );
   gpc606_5 gpc582 (
      {stage0_28[181], stage0_28[182], stage0_28[183], stage0_28[184], stage0_28[185], stage0_28[186]},
      {stage0_30[145], stage0_30[146], stage0_30[147], stage0_30[148], stage0_30[149], stage0_30[150]},
      {stage1_32[25],stage1_31[41],stage1_30[44],stage1_29[67],stage1_28[97]}
   );
   gpc606_5 gpc583 (
      {stage0_28[187], stage0_28[188], stage0_28[189], stage0_28[190], stage0_28[191], stage0_28[192]},
      {stage0_30[151], stage0_30[152], stage0_30[153], stage0_30[154], stage0_30[155], stage0_30[156]},
      {stage1_32[26],stage1_31[42],stage1_30[45],stage1_29[68],stage1_28[98]}
   );
   gpc606_5 gpc584 (
      {stage0_28[193], stage0_28[194], stage0_28[195], stage0_28[196], stage0_28[197], stage0_28[198]},
      {stage0_30[157], stage0_30[158], stage0_30[159], stage0_30[160], stage0_30[161], stage0_30[162]},
      {stage1_32[27],stage1_31[43],stage1_30[46],stage1_29[69],stage1_28[99]}
   );
   gpc606_5 gpc585 (
      {stage0_28[199], stage0_28[200], stage0_28[201], stage0_28[202], stage0_28[203], stage0_28[204]},
      {stage0_30[163], stage0_30[164], stage0_30[165], stage0_30[166], stage0_30[167], stage0_30[168]},
      {stage1_32[28],stage1_31[44],stage1_30[47],stage1_29[70],stage1_28[100]}
   );
   gpc606_5 gpc586 (
      {stage0_28[205], stage0_28[206], stage0_28[207], stage0_28[208], stage0_28[209], stage0_28[210]},
      {stage0_30[169], stage0_30[170], stage0_30[171], stage0_30[172], stage0_30[173], stage0_30[174]},
      {stage1_32[29],stage1_31[45],stage1_30[48],stage1_29[71],stage1_28[101]}
   );
   gpc606_5 gpc587 (
      {stage0_28[211], stage0_28[212], stage0_28[213], stage0_28[214], stage0_28[215], stage0_28[216]},
      {stage0_30[175], stage0_30[176], stage0_30[177], stage0_30[178], stage0_30[179], stage0_30[180]},
      {stage1_32[30],stage1_31[46],stage1_30[49],stage1_29[72],stage1_28[102]}
   );
   gpc606_5 gpc588 (
      {stage0_28[217], stage0_28[218], stage0_28[219], stage0_28[220], stage0_28[221], stage0_28[222]},
      {stage0_30[181], stage0_30[182], stage0_30[183], stage0_30[184], stage0_30[185], stage0_30[186]},
      {stage1_32[31],stage1_31[47],stage1_30[50],stage1_29[73],stage1_28[103]}
   );
   gpc606_5 gpc589 (
      {stage0_28[223], stage0_28[224], stage0_28[225], stage0_28[226], stage0_28[227], stage0_28[228]},
      {stage0_30[187], stage0_30[188], stage0_30[189], stage0_30[190], stage0_30[191], stage0_30[192]},
      {stage1_32[32],stage1_31[48],stage1_30[51],stage1_29[74],stage1_28[104]}
   );
   gpc606_5 gpc590 (
      {stage0_28[229], stage0_28[230], stage0_28[231], stage0_28[232], stage0_28[233], stage0_28[234]},
      {stage0_30[193], stage0_30[194], stage0_30[195], stage0_30[196], stage0_30[197], stage0_30[198]},
      {stage1_32[33],stage1_31[49],stage1_30[52],stage1_29[75],stage1_28[105]}
   );
   gpc606_5 gpc591 (
      {stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101], stage0_29[102]},
      {stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6], stage0_31[7]},
      {stage1_33[0],stage1_32[34],stage1_31[50],stage1_30[53],stage1_29[76]}
   );
   gpc606_5 gpc592 (
      {stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107], stage0_29[108]},
      {stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12], stage0_31[13]},
      {stage1_33[1],stage1_32[35],stage1_31[51],stage1_30[54],stage1_29[77]}
   );
   gpc606_5 gpc593 (
      {stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113], stage0_29[114]},
      {stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17], stage0_31[18], stage0_31[19]},
      {stage1_33[2],stage1_32[36],stage1_31[52],stage1_30[55],stage1_29[78]}
   );
   gpc606_5 gpc594 (
      {stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119], stage0_29[120]},
      {stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23], stage0_31[24], stage0_31[25]},
      {stage1_33[3],stage1_32[37],stage1_31[53],stage1_30[56],stage1_29[79]}
   );
   gpc606_5 gpc595 (
      {stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125], stage0_29[126]},
      {stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29], stage0_31[30], stage0_31[31]},
      {stage1_33[4],stage1_32[38],stage1_31[54],stage1_30[57],stage1_29[80]}
   );
   gpc606_5 gpc596 (
      {stage0_29[127], stage0_29[128], stage0_29[129], stage0_29[130], stage0_29[131], stage0_29[132]},
      {stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35], stage0_31[36], stage0_31[37]},
      {stage1_33[5],stage1_32[39],stage1_31[55],stage1_30[58],stage1_29[81]}
   );
   gpc606_5 gpc597 (
      {stage0_29[133], stage0_29[134], stage0_29[135], stage0_29[136], stage0_29[137], stage0_29[138]},
      {stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41], stage0_31[42], stage0_31[43]},
      {stage1_33[6],stage1_32[40],stage1_31[56],stage1_30[59],stage1_29[82]}
   );
   gpc606_5 gpc598 (
      {stage0_29[139], stage0_29[140], stage0_29[141], stage0_29[142], stage0_29[143], stage0_29[144]},
      {stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47], stage0_31[48], stage0_31[49]},
      {stage1_33[7],stage1_32[41],stage1_31[57],stage1_30[60],stage1_29[83]}
   );
   gpc606_5 gpc599 (
      {stage0_29[145], stage0_29[146], stage0_29[147], stage0_29[148], stage0_29[149], stage0_29[150]},
      {stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53], stage0_31[54], stage0_31[55]},
      {stage1_33[8],stage1_32[42],stage1_31[58],stage1_30[61],stage1_29[84]}
   );
   gpc606_5 gpc600 (
      {stage0_29[151], stage0_29[152], stage0_29[153], stage0_29[154], stage0_29[155], stage0_29[156]},
      {stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59], stage0_31[60], stage0_31[61]},
      {stage1_33[9],stage1_32[43],stage1_31[59],stage1_30[62],stage1_29[85]}
   );
   gpc606_5 gpc601 (
      {stage0_29[157], stage0_29[158], stage0_29[159], stage0_29[160], stage0_29[161], stage0_29[162]},
      {stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65], stage0_31[66], stage0_31[67]},
      {stage1_33[10],stage1_32[44],stage1_31[60],stage1_30[63],stage1_29[86]}
   );
   gpc606_5 gpc602 (
      {stage0_29[163], stage0_29[164], stage0_29[165], stage0_29[166], stage0_29[167], stage0_29[168]},
      {stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71], stage0_31[72], stage0_31[73]},
      {stage1_33[11],stage1_32[45],stage1_31[61],stage1_30[64],stage1_29[87]}
   );
   gpc606_5 gpc603 (
      {stage0_29[169], stage0_29[170], stage0_29[171], stage0_29[172], stage0_29[173], stage0_29[174]},
      {stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77], stage0_31[78], stage0_31[79]},
      {stage1_33[12],stage1_32[46],stage1_31[62],stage1_30[65],stage1_29[88]}
   );
   gpc606_5 gpc604 (
      {stage0_29[175], stage0_29[176], stage0_29[177], stage0_29[178], stage0_29[179], stage0_29[180]},
      {stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83], stage0_31[84], stage0_31[85]},
      {stage1_33[13],stage1_32[47],stage1_31[63],stage1_30[66],stage1_29[89]}
   );
   gpc606_5 gpc605 (
      {stage0_29[181], stage0_29[182], stage0_29[183], stage0_29[184], stage0_29[185], stage0_29[186]},
      {stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89], stage0_31[90], stage0_31[91]},
      {stage1_33[14],stage1_32[48],stage1_31[64],stage1_30[67],stage1_29[90]}
   );
   gpc606_5 gpc606 (
      {stage0_29[187], stage0_29[188], stage0_29[189], stage0_29[190], stage0_29[191], stage0_29[192]},
      {stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95], stage0_31[96], stage0_31[97]},
      {stage1_33[15],stage1_32[49],stage1_31[65],stage1_30[68],stage1_29[91]}
   );
   gpc606_5 gpc607 (
      {stage0_29[193], stage0_29[194], stage0_29[195], stage0_29[196], stage0_29[197], stage0_29[198]},
      {stage0_31[98], stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage1_33[16],stage1_32[50],stage1_31[66],stage1_30[69],stage1_29[92]}
   );
   gpc606_5 gpc608 (
      {stage0_29[199], stage0_29[200], stage0_29[201], stage0_29[202], stage0_29[203], stage0_29[204]},
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108], stage0_31[109]},
      {stage1_33[17],stage1_32[51],stage1_31[67],stage1_30[70],stage1_29[93]}
   );
   gpc606_5 gpc609 (
      {stage0_29[205], stage0_29[206], stage0_29[207], stage0_29[208], stage0_29[209], stage0_29[210]},
      {stage0_31[110], stage0_31[111], stage0_31[112], stage0_31[113], stage0_31[114], stage0_31[115]},
      {stage1_33[18],stage1_32[52],stage1_31[68],stage1_30[71],stage1_29[94]}
   );
   gpc606_5 gpc610 (
      {stage0_29[211], stage0_29[212], stage0_29[213], stage0_29[214], stage0_29[215], stage0_29[216]},
      {stage0_31[116], stage0_31[117], stage0_31[118], stage0_31[119], stage0_31[120], stage0_31[121]},
      {stage1_33[19],stage1_32[53],stage1_31[69],stage1_30[72],stage1_29[95]}
   );
   gpc606_5 gpc611 (
      {stage0_29[217], stage0_29[218], stage0_29[219], stage0_29[220], stage0_29[221], stage0_29[222]},
      {stage0_31[122], stage0_31[123], stage0_31[124], stage0_31[125], stage0_31[126], stage0_31[127]},
      {stage1_33[20],stage1_32[54],stage1_31[70],stage1_30[73],stage1_29[96]}
   );
   gpc606_5 gpc612 (
      {stage0_29[223], stage0_29[224], stage0_29[225], stage0_29[226], stage0_29[227], stage0_29[228]},
      {stage0_31[128], stage0_31[129], stage0_31[130], stage0_31[131], stage0_31[132], stage0_31[133]},
      {stage1_33[21],stage1_32[55],stage1_31[71],stage1_30[74],stage1_29[97]}
   );
   gpc606_5 gpc613 (
      {stage0_29[229], stage0_29[230], stage0_29[231], stage0_29[232], stage0_29[233], stage0_29[234]},
      {stage0_31[134], stage0_31[135], stage0_31[136], stage0_31[137], stage0_31[138], stage0_31[139]},
      {stage1_33[22],stage1_32[56],stage1_31[72],stage1_30[75],stage1_29[98]}
   );
   gpc606_5 gpc614 (
      {stage0_29[235], stage0_29[236], stage0_29[237], stage0_29[238], stage0_29[239], stage0_29[240]},
      {stage0_31[140], stage0_31[141], stage0_31[142], stage0_31[143], stage0_31[144], stage0_31[145]},
      {stage1_33[23],stage1_32[57],stage1_31[73],stage1_30[76],stage1_29[99]}
   );
   gpc606_5 gpc615 (
      {stage0_29[241], stage0_29[242], stage0_29[243], stage0_29[244], stage0_29[245], stage0_29[246]},
      {stage0_31[146], stage0_31[147], stage0_31[148], stage0_31[149], stage0_31[150], stage0_31[151]},
      {stage1_33[24],stage1_32[58],stage1_31[74],stage1_30[77],stage1_29[100]}
   );
   gpc615_5 gpc616 (
      {stage0_30[199], stage0_30[200], stage0_30[201], stage0_30[202], stage0_30[203]},
      {stage0_31[152]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[25],stage1_32[59],stage1_31[75],stage1_30[78]}
   );
   gpc615_5 gpc617 (
      {stage0_30[204], stage0_30[205], stage0_30[206], stage0_30[207], stage0_30[208]},
      {stage0_31[153]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[26],stage1_32[60],stage1_31[76],stage1_30[79]}
   );
   gpc615_5 gpc618 (
      {stage0_30[209], stage0_30[210], stage0_30[211], stage0_30[212], stage0_30[213]},
      {stage0_31[154]},
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage1_34[2],stage1_33[27],stage1_32[61],stage1_31[77],stage1_30[80]}
   );
   gpc615_5 gpc619 (
      {stage0_30[214], stage0_30[215], stage0_30[216], stage0_30[217], stage0_30[218]},
      {stage0_31[155]},
      {stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21], stage0_32[22], stage0_32[23]},
      {stage1_34[3],stage1_33[28],stage1_32[62],stage1_31[78],stage1_30[81]}
   );
   gpc615_5 gpc620 (
      {stage0_30[219], stage0_30[220], stage0_30[221], stage0_30[222], stage0_30[223]},
      {stage0_31[156]},
      {stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27], stage0_32[28], stage0_32[29]},
      {stage1_34[4],stage1_33[29],stage1_32[63],stage1_31[79],stage1_30[82]}
   );
   gpc615_5 gpc621 (
      {stage0_30[224], stage0_30[225], stage0_30[226], stage0_30[227], stage0_30[228]},
      {stage0_31[157]},
      {stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33], stage0_32[34], stage0_32[35]},
      {stage1_34[5],stage1_33[30],stage1_32[64],stage1_31[80],stage1_30[83]}
   );
   gpc615_5 gpc622 (
      {stage0_30[229], stage0_30[230], stage0_30[231], stage0_30[232], stage0_30[233]},
      {stage0_31[158]},
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage1_34[6],stage1_33[31],stage1_32[65],stage1_31[81],stage1_30[84]}
   );
   gpc615_5 gpc623 (
      {stage0_30[234], stage0_30[235], stage0_30[236], stage0_30[237], stage0_30[238]},
      {stage0_31[159]},
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage1_34[7],stage1_33[32],stage1_32[66],stage1_31[82],stage1_30[85]}
   );
   gpc615_5 gpc624 (
      {stage0_30[239], stage0_30[240], stage0_30[241], stage0_30[242], stage0_30[243]},
      {stage0_31[160]},
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52], stage0_32[53]},
      {stage1_34[8],stage1_33[33],stage1_32[67],stage1_31[83],stage1_30[86]}
   );
   gpc615_5 gpc625 (
      {stage0_30[244], stage0_30[245], stage0_30[246], stage0_30[247], stage0_30[248]},
      {stage0_31[161]},
      {stage0_32[54], stage0_32[55], stage0_32[56], stage0_32[57], stage0_32[58], stage0_32[59]},
      {stage1_34[9],stage1_33[34],stage1_32[68],stage1_31[84],stage1_30[87]}
   );
   gpc615_5 gpc626 (
      {stage0_30[249], stage0_30[250], stage0_30[251], stage0_30[252], stage0_30[253]},
      {stage0_31[162]},
      {stage0_32[60], stage0_32[61], stage0_32[62], stage0_32[63], stage0_32[64], stage0_32[65]},
      {stage1_34[10],stage1_33[35],stage1_32[69],stage1_31[85],stage1_30[88]}
   );
   gpc615_5 gpc627 (
      {stage0_31[163], stage0_31[164], stage0_31[165], stage0_31[166], stage0_31[167]},
      {stage0_32[66]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[11],stage1_33[36],stage1_32[70],stage1_31[86]}
   );
   gpc615_5 gpc628 (
      {stage0_31[168], stage0_31[169], stage0_31[170], stage0_31[171], stage0_31[172]},
      {stage0_32[67]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[12],stage1_33[37],stage1_32[71],stage1_31[87]}
   );
   gpc615_5 gpc629 (
      {stage0_31[173], stage0_31[174], stage0_31[175], stage0_31[176], stage0_31[177]},
      {stage0_32[68]},
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage1_35[2],stage1_34[13],stage1_33[38],stage1_32[72],stage1_31[88]}
   );
   gpc615_5 gpc630 (
      {stage0_31[178], stage0_31[179], stage0_31[180], stage0_31[181], stage0_31[182]},
      {stage0_32[69]},
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage1_35[3],stage1_34[14],stage1_33[39],stage1_32[73],stage1_31[89]}
   );
   gpc615_5 gpc631 (
      {stage0_31[183], stage0_31[184], stage0_31[185], stage0_31[186], stage0_31[187]},
      {stage0_32[70]},
      {stage0_33[24], stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29]},
      {stage1_35[4],stage1_34[15],stage1_33[40],stage1_32[74],stage1_31[90]}
   );
   gpc615_5 gpc632 (
      {stage0_31[188], stage0_31[189], stage0_31[190], stage0_31[191], stage0_31[192]},
      {stage0_32[71]},
      {stage0_33[30], stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35]},
      {stage1_35[5],stage1_34[16],stage1_33[41],stage1_32[75],stage1_31[91]}
   );
   gpc615_5 gpc633 (
      {stage0_31[193], stage0_31[194], stage0_31[195], stage0_31[196], stage0_31[197]},
      {stage0_32[72]},
      {stage0_33[36], stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41]},
      {stage1_35[6],stage1_34[17],stage1_33[42],stage1_32[76],stage1_31[92]}
   );
   gpc615_5 gpc634 (
      {stage0_31[198], stage0_31[199], stage0_31[200], stage0_31[201], stage0_31[202]},
      {stage0_32[73]},
      {stage0_33[42], stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47]},
      {stage1_35[7],stage1_34[18],stage1_33[43],stage1_32[77],stage1_31[93]}
   );
   gpc615_5 gpc635 (
      {stage0_31[203], stage0_31[204], stage0_31[205], stage0_31[206], stage0_31[207]},
      {stage0_32[74]},
      {stage0_33[48], stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53]},
      {stage1_35[8],stage1_34[19],stage1_33[44],stage1_32[78],stage1_31[94]}
   );
   gpc615_5 gpc636 (
      {stage0_31[208], stage0_31[209], stage0_31[210], stage0_31[211], stage0_31[212]},
      {stage0_32[75]},
      {stage0_33[54], stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59]},
      {stage1_35[9],stage1_34[20],stage1_33[45],stage1_32[79],stage1_31[95]}
   );
   gpc615_5 gpc637 (
      {stage0_31[213], stage0_31[214], stage0_31[215], stage0_31[216], stage0_31[217]},
      {stage0_32[76]},
      {stage0_33[60], stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65]},
      {stage1_35[10],stage1_34[21],stage1_33[46],stage1_32[80],stage1_31[96]}
   );
   gpc615_5 gpc638 (
      {stage0_31[218], stage0_31[219], stage0_31[220], stage0_31[221], stage0_31[222]},
      {stage0_32[77]},
      {stage0_33[66], stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71]},
      {stage1_35[11],stage1_34[22],stage1_33[47],stage1_32[81],stage1_31[97]}
   );
   gpc615_5 gpc639 (
      {stage0_31[223], stage0_31[224], stage0_31[225], stage0_31[226], stage0_31[227]},
      {stage0_32[78]},
      {stage0_33[72], stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77]},
      {stage1_35[12],stage1_34[23],stage1_33[48],stage1_32[82],stage1_31[98]}
   );
   gpc615_5 gpc640 (
      {stage0_31[228], stage0_31[229], stage0_31[230], stage0_31[231], stage0_31[232]},
      {stage0_32[79]},
      {stage0_33[78], stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83]},
      {stage1_35[13],stage1_34[24],stage1_33[49],stage1_32[83],stage1_31[99]}
   );
   gpc615_5 gpc641 (
      {stage0_31[233], stage0_31[234], stage0_31[235], stage0_31[236], stage0_31[237]},
      {stage0_32[80]},
      {stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88], stage0_33[89]},
      {stage1_35[14],stage1_34[25],stage1_33[50],stage1_32[84],stage1_31[100]}
   );
   gpc615_5 gpc642 (
      {stage0_31[238], stage0_31[239], stage0_31[240], stage0_31[241], stage0_31[242]},
      {stage0_32[81]},
      {stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93], stage0_33[94], stage0_33[95]},
      {stage1_35[15],stage1_34[26],stage1_33[51],stage1_32[85],stage1_31[101]}
   );
   gpc606_5 gpc643 (
      {stage0_32[82], stage0_32[83], stage0_32[84], stage0_32[85], stage0_32[86], stage0_32[87]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[16],stage1_34[27],stage1_33[52],stage1_32[86]}
   );
   gpc606_5 gpc644 (
      {stage0_32[88], stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92], stage0_32[93]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[17],stage1_34[28],stage1_33[53],stage1_32[87]}
   );
   gpc606_5 gpc645 (
      {stage0_32[94], stage0_32[95], stage0_32[96], stage0_32[97], stage0_32[98], stage0_32[99]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[18],stage1_34[29],stage1_33[54],stage1_32[88]}
   );
   gpc606_5 gpc646 (
      {stage0_32[100], stage0_32[101], stage0_32[102], stage0_32[103], stage0_32[104], stage0_32[105]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[19],stage1_34[30],stage1_33[55],stage1_32[89]}
   );
   gpc606_5 gpc647 (
      {stage0_32[106], stage0_32[107], stage0_32[108], stage0_32[109], stage0_32[110], stage0_32[111]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[20],stage1_34[31],stage1_33[56],stage1_32[90]}
   );
   gpc606_5 gpc648 (
      {stage0_32[112], stage0_32[113], stage0_32[114], stage0_32[115], stage0_32[116], stage0_32[117]},
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35]},
      {stage1_36[5],stage1_35[21],stage1_34[32],stage1_33[57],stage1_32[91]}
   );
   gpc606_5 gpc649 (
      {stage0_32[118], stage0_32[119], stage0_32[120], stage0_32[121], stage0_32[122], stage0_32[123]},
      {stage0_34[36], stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41]},
      {stage1_36[6],stage1_35[22],stage1_34[33],stage1_33[58],stage1_32[92]}
   );
   gpc606_5 gpc650 (
      {stage0_32[124], stage0_32[125], stage0_32[126], stage0_32[127], stage0_32[128], stage0_32[129]},
      {stage0_34[42], stage0_34[43], stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47]},
      {stage1_36[7],stage1_35[23],stage1_34[34],stage1_33[59],stage1_32[93]}
   );
   gpc606_5 gpc651 (
      {stage0_32[130], stage0_32[131], stage0_32[132], stage0_32[133], stage0_32[134], stage0_32[135]},
      {stage0_34[48], stage0_34[49], stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53]},
      {stage1_36[8],stage1_35[24],stage1_34[35],stage1_33[60],stage1_32[94]}
   );
   gpc606_5 gpc652 (
      {stage0_32[136], stage0_32[137], stage0_32[138], stage0_32[139], stage0_32[140], stage0_32[141]},
      {stage0_34[54], stage0_34[55], stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59]},
      {stage1_36[9],stage1_35[25],stage1_34[36],stage1_33[61],stage1_32[95]}
   );
   gpc606_5 gpc653 (
      {stage0_32[142], stage0_32[143], stage0_32[144], stage0_32[145], stage0_32[146], stage0_32[147]},
      {stage0_34[60], stage0_34[61], stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65]},
      {stage1_36[10],stage1_35[26],stage1_34[37],stage1_33[62],stage1_32[96]}
   );
   gpc606_5 gpc654 (
      {stage0_32[148], stage0_32[149], stage0_32[150], stage0_32[151], stage0_32[152], stage0_32[153]},
      {stage0_34[66], stage0_34[67], stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71]},
      {stage1_36[11],stage1_35[27],stage1_34[38],stage1_33[63],stage1_32[97]}
   );
   gpc606_5 gpc655 (
      {stage0_32[154], stage0_32[155], stage0_32[156], stage0_32[157], stage0_32[158], stage0_32[159]},
      {stage0_34[72], stage0_34[73], stage0_34[74], stage0_34[75], stage0_34[76], stage0_34[77]},
      {stage1_36[12],stage1_35[28],stage1_34[39],stage1_33[64],stage1_32[98]}
   );
   gpc606_5 gpc656 (
      {stage0_32[160], stage0_32[161], stage0_32[162], stage0_32[163], stage0_32[164], stage0_32[165]},
      {stage0_34[78], stage0_34[79], stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83]},
      {stage1_36[13],stage1_35[29],stage1_34[40],stage1_33[65],stage1_32[99]}
   );
   gpc606_5 gpc657 (
      {stage0_32[166], stage0_32[167], stage0_32[168], stage0_32[169], stage0_32[170], stage0_32[171]},
      {stage0_34[84], stage0_34[85], stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89]},
      {stage1_36[14],stage1_35[30],stage1_34[41],stage1_33[66],stage1_32[100]}
   );
   gpc606_5 gpc658 (
      {stage0_32[172], stage0_32[173], stage0_32[174], stage0_32[175], stage0_32[176], stage0_32[177]},
      {stage0_34[90], stage0_34[91], stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95]},
      {stage1_36[15],stage1_35[31],stage1_34[42],stage1_33[67],stage1_32[101]}
   );
   gpc606_5 gpc659 (
      {stage0_32[178], stage0_32[179], stage0_32[180], stage0_32[181], stage0_32[182], stage0_32[183]},
      {stage0_34[96], stage0_34[97], stage0_34[98], stage0_34[99], stage0_34[100], stage0_34[101]},
      {stage1_36[16],stage1_35[32],stage1_34[43],stage1_33[68],stage1_32[102]}
   );
   gpc606_5 gpc660 (
      {stage0_32[184], stage0_32[185], stage0_32[186], stage0_32[187], stage0_32[188], stage0_32[189]},
      {stage0_34[102], stage0_34[103], stage0_34[104], stage0_34[105], stage0_34[106], stage0_34[107]},
      {stage1_36[17],stage1_35[33],stage1_34[44],stage1_33[69],stage1_32[103]}
   );
   gpc606_5 gpc661 (
      {stage0_32[190], stage0_32[191], stage0_32[192], stage0_32[193], stage0_32[194], stage0_32[195]},
      {stage0_34[108], stage0_34[109], stage0_34[110], stage0_34[111], stage0_34[112], stage0_34[113]},
      {stage1_36[18],stage1_35[34],stage1_34[45],stage1_33[70],stage1_32[104]}
   );
   gpc606_5 gpc662 (
      {stage0_32[196], stage0_32[197], stage0_32[198], stage0_32[199], stage0_32[200], stage0_32[201]},
      {stage0_34[114], stage0_34[115], stage0_34[116], stage0_34[117], stage0_34[118], stage0_34[119]},
      {stage1_36[19],stage1_35[35],stage1_34[46],stage1_33[71],stage1_32[105]}
   );
   gpc606_5 gpc663 (
      {stage0_32[202], stage0_32[203], stage0_32[204], stage0_32[205], stage0_32[206], stage0_32[207]},
      {stage0_34[120], stage0_34[121], stage0_34[122], stage0_34[123], stage0_34[124], stage0_34[125]},
      {stage1_36[20],stage1_35[36],stage1_34[47],stage1_33[72],stage1_32[106]}
   );
   gpc606_5 gpc664 (
      {stage0_32[208], stage0_32[209], stage0_32[210], stage0_32[211], stage0_32[212], stage0_32[213]},
      {stage0_34[126], stage0_34[127], stage0_34[128], stage0_34[129], stage0_34[130], stage0_34[131]},
      {stage1_36[21],stage1_35[37],stage1_34[48],stage1_33[73],stage1_32[107]}
   );
   gpc606_5 gpc665 (
      {stage0_32[214], stage0_32[215], stage0_32[216], stage0_32[217], stage0_32[218], stage0_32[219]},
      {stage0_34[132], stage0_34[133], stage0_34[134], stage0_34[135], stage0_34[136], stage0_34[137]},
      {stage1_36[22],stage1_35[38],stage1_34[49],stage1_33[74],stage1_32[108]}
   );
   gpc606_5 gpc666 (
      {stage0_32[220], stage0_32[221], stage0_32[222], stage0_32[223], stage0_32[224], stage0_32[225]},
      {stage0_34[138], stage0_34[139], stage0_34[140], stage0_34[141], stage0_34[142], stage0_34[143]},
      {stage1_36[23],stage1_35[39],stage1_34[50],stage1_33[75],stage1_32[109]}
   );
   gpc606_5 gpc667 (
      {stage0_32[226], stage0_32[227], stage0_32[228], stage0_32[229], stage0_32[230], stage0_32[231]},
      {stage0_34[144], stage0_34[145], stage0_34[146], stage0_34[147], stage0_34[148], stage0_34[149]},
      {stage1_36[24],stage1_35[40],stage1_34[51],stage1_33[76],stage1_32[110]}
   );
   gpc606_5 gpc668 (
      {stage0_32[232], stage0_32[233], stage0_32[234], stage0_32[235], stage0_32[236], stage0_32[237]},
      {stage0_34[150], stage0_34[151], stage0_34[152], stage0_34[153], stage0_34[154], stage0_34[155]},
      {stage1_36[25],stage1_35[41],stage1_34[52],stage1_33[77],stage1_32[111]}
   );
   gpc606_5 gpc669 (
      {stage0_32[238], stage0_32[239], stage0_32[240], stage0_32[241], stage0_32[242], stage0_32[243]},
      {stage0_34[156], stage0_34[157], stage0_34[158], stage0_34[159], stage0_34[160], stage0_34[161]},
      {stage1_36[26],stage1_35[42],stage1_34[53],stage1_33[78],stage1_32[112]}
   );
   gpc606_5 gpc670 (
      {stage0_32[244], stage0_32[245], stage0_32[246], stage0_32[247], stage0_32[248], stage0_32[249]},
      {stage0_34[162], stage0_34[163], stage0_34[164], stage0_34[165], stage0_34[166], stage0_34[167]},
      {stage1_36[27],stage1_35[43],stage1_34[54],stage1_33[79],stage1_32[113]}
   );
   gpc606_5 gpc671 (
      {stage0_32[250], stage0_32[251], stage0_32[252], stage0_32[253], stage0_32[254], stage0_32[255]},
      {stage0_34[168], stage0_34[169], stage0_34[170], stage0_34[171], stage0_34[172], stage0_34[173]},
      {stage1_36[28],stage1_35[44],stage1_34[55],stage1_33[80],stage1_32[114]}
   );
   gpc606_5 gpc672 (
      {stage0_33[96], stage0_33[97], stage0_33[98], stage0_33[99], stage0_33[100], stage0_33[101]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[29],stage1_35[45],stage1_34[56],stage1_33[81]}
   );
   gpc606_5 gpc673 (
      {stage0_33[102], stage0_33[103], stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[30],stage1_35[46],stage1_34[57],stage1_33[82]}
   );
   gpc606_5 gpc674 (
      {stage0_33[108], stage0_33[109], stage0_33[110], stage0_33[111], stage0_33[112], stage0_33[113]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[31],stage1_35[47],stage1_34[58],stage1_33[83]}
   );
   gpc606_5 gpc675 (
      {stage0_33[114], stage0_33[115], stage0_33[116], stage0_33[117], stage0_33[118], stage0_33[119]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[32],stage1_35[48],stage1_34[59],stage1_33[84]}
   );
   gpc606_5 gpc676 (
      {stage0_33[120], stage0_33[121], stage0_33[122], stage0_33[123], stage0_33[124], stage0_33[125]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[33],stage1_35[49],stage1_34[60],stage1_33[85]}
   );
   gpc606_5 gpc677 (
      {stage0_33[126], stage0_33[127], stage0_33[128], stage0_33[129], stage0_33[130], stage0_33[131]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[34],stage1_35[50],stage1_34[61],stage1_33[86]}
   );
   gpc606_5 gpc678 (
      {stage0_33[132], stage0_33[133], stage0_33[134], stage0_33[135], stage0_33[136], stage0_33[137]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[35],stage1_35[51],stage1_34[62],stage1_33[87]}
   );
   gpc606_5 gpc679 (
      {stage0_33[138], stage0_33[139], stage0_33[140], stage0_33[141], stage0_33[142], stage0_33[143]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[36],stage1_35[52],stage1_34[63],stage1_33[88]}
   );
   gpc606_5 gpc680 (
      {stage0_33[144], stage0_33[145], stage0_33[146], stage0_33[147], stage0_33[148], stage0_33[149]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[37],stage1_35[53],stage1_34[64],stage1_33[89]}
   );
   gpc606_5 gpc681 (
      {stage0_33[150], stage0_33[151], stage0_33[152], stage0_33[153], stage0_33[154], stage0_33[155]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[38],stage1_35[54],stage1_34[65],stage1_33[90]}
   );
   gpc606_5 gpc682 (
      {stage0_33[156], stage0_33[157], stage0_33[158], stage0_33[159], stage0_33[160], stage0_33[161]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[39],stage1_35[55],stage1_34[66],stage1_33[91]}
   );
   gpc606_5 gpc683 (
      {stage0_33[162], stage0_33[163], stage0_33[164], stage0_33[165], stage0_33[166], stage0_33[167]},
      {stage0_35[66], stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage1_37[11],stage1_36[40],stage1_35[56],stage1_34[67],stage1_33[92]}
   );
   gpc606_5 gpc684 (
      {stage0_33[168], stage0_33[169], stage0_33[170], stage0_33[171], stage0_33[172], stage0_33[173]},
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76], stage0_35[77]},
      {stage1_37[12],stage1_36[41],stage1_35[57],stage1_34[68],stage1_33[93]}
   );
   gpc606_5 gpc685 (
      {stage0_33[174], stage0_33[175], stage0_33[176], stage0_33[177], stage0_33[178], stage0_33[179]},
      {stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81], stage0_35[82], stage0_35[83]},
      {stage1_37[13],stage1_36[42],stage1_35[58],stage1_34[69],stage1_33[94]}
   );
   gpc606_5 gpc686 (
      {stage0_33[180], stage0_33[181], stage0_33[182], stage0_33[183], stage0_33[184], stage0_33[185]},
      {stage0_35[84], stage0_35[85], stage0_35[86], stage0_35[87], stage0_35[88], stage0_35[89]},
      {stage1_37[14],stage1_36[43],stage1_35[59],stage1_34[70],stage1_33[95]}
   );
   gpc606_5 gpc687 (
      {stage0_33[186], stage0_33[187], stage0_33[188], stage0_33[189], stage0_33[190], stage0_33[191]},
      {stage0_35[90], stage0_35[91], stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95]},
      {stage1_37[15],stage1_36[44],stage1_35[60],stage1_34[71],stage1_33[96]}
   );
   gpc606_5 gpc688 (
      {stage0_33[192], stage0_33[193], stage0_33[194], stage0_33[195], stage0_33[196], stage0_33[197]},
      {stage0_35[96], stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage1_37[16],stage1_36[45],stage1_35[61],stage1_34[72],stage1_33[97]}
   );
   gpc606_5 gpc689 (
      {stage0_33[198], stage0_33[199], stage0_33[200], stage0_33[201], stage0_33[202], stage0_33[203]},
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106], stage0_35[107]},
      {stage1_37[17],stage1_36[46],stage1_35[62],stage1_34[73],stage1_33[98]}
   );
   gpc606_5 gpc690 (
      {stage0_33[204], stage0_33[205], stage0_33[206], stage0_33[207], stage0_33[208], stage0_33[209]},
      {stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111], stage0_35[112], stage0_35[113]},
      {stage1_37[18],stage1_36[47],stage1_35[63],stage1_34[74],stage1_33[99]}
   );
   gpc606_5 gpc691 (
      {stage0_33[210], stage0_33[211], stage0_33[212], stage0_33[213], stage0_33[214], stage0_33[215]},
      {stage0_35[114], stage0_35[115], stage0_35[116], stage0_35[117], stage0_35[118], stage0_35[119]},
      {stage1_37[19],stage1_36[48],stage1_35[64],stage1_34[75],stage1_33[100]}
   );
   gpc606_5 gpc692 (
      {stage0_33[216], stage0_33[217], stage0_33[218], stage0_33[219], stage0_33[220], stage0_33[221]},
      {stage0_35[120], stage0_35[121], stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125]},
      {stage1_37[20],stage1_36[49],stage1_35[65],stage1_34[76],stage1_33[101]}
   );
   gpc606_5 gpc693 (
      {stage0_33[222], stage0_33[223], stage0_33[224], stage0_33[225], stage0_33[226], stage0_33[227]},
      {stage0_35[126], stage0_35[127], stage0_35[128], stage0_35[129], stage0_35[130], stage0_35[131]},
      {stage1_37[21],stage1_36[50],stage1_35[66],stage1_34[77],stage1_33[102]}
   );
   gpc606_5 gpc694 (
      {stage0_33[228], stage0_33[229], stage0_33[230], stage0_33[231], stage0_33[232], stage0_33[233]},
      {stage0_35[132], stage0_35[133], stage0_35[134], stage0_35[135], stage0_35[136], stage0_35[137]},
      {stage1_37[22],stage1_36[51],stage1_35[67],stage1_34[78],stage1_33[103]}
   );
   gpc606_5 gpc695 (
      {stage0_33[234], stage0_33[235], stage0_33[236], stage0_33[237], stage0_33[238], stage0_33[239]},
      {stage0_35[138], stage0_35[139], stage0_35[140], stage0_35[141], stage0_35[142], stage0_35[143]},
      {stage1_37[23],stage1_36[52],stage1_35[68],stage1_34[79],stage1_33[104]}
   );
   gpc606_5 gpc696 (
      {stage0_33[240], stage0_33[241], stage0_33[242], stage0_33[243], stage0_33[244], stage0_33[245]},
      {stage0_35[144], stage0_35[145], stage0_35[146], stage0_35[147], stage0_35[148], stage0_35[149]},
      {stage1_37[24],stage1_36[53],stage1_35[69],stage1_34[80],stage1_33[105]}
   );
   gpc606_5 gpc697 (
      {stage0_33[246], stage0_33[247], stage0_33[248], stage0_33[249], stage0_33[250], stage0_33[251]},
      {stage0_35[150], stage0_35[151], stage0_35[152], stage0_35[153], stage0_35[154], stage0_35[155]},
      {stage1_37[25],stage1_36[54],stage1_35[70],stage1_34[81],stage1_33[106]}
   );
   gpc615_5 gpc698 (
      {stage0_34[174], stage0_34[175], stage0_34[176], stage0_34[177], stage0_34[178]},
      {stage0_35[156]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[26],stage1_36[55],stage1_35[71],stage1_34[82]}
   );
   gpc615_5 gpc699 (
      {stage0_34[179], stage0_34[180], stage0_34[181], stage0_34[182], stage0_34[183]},
      {stage0_35[157]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[27],stage1_36[56],stage1_35[72],stage1_34[83]}
   );
   gpc615_5 gpc700 (
      {stage0_34[184], stage0_34[185], stage0_34[186], stage0_34[187], stage0_34[188]},
      {stage0_35[158]},
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17]},
      {stage1_38[2],stage1_37[28],stage1_36[57],stage1_35[73],stage1_34[84]}
   );
   gpc615_5 gpc701 (
      {stage0_34[189], stage0_34[190], stage0_34[191], stage0_34[192], stage0_34[193]},
      {stage0_35[159]},
      {stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23]},
      {stage1_38[3],stage1_37[29],stage1_36[58],stage1_35[74],stage1_34[85]}
   );
   gpc615_5 gpc702 (
      {stage0_34[194], stage0_34[195], stage0_34[196], stage0_34[197], stage0_34[198]},
      {stage0_35[160]},
      {stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29]},
      {stage1_38[4],stage1_37[30],stage1_36[59],stage1_35[75],stage1_34[86]}
   );
   gpc615_5 gpc703 (
      {stage0_34[199], stage0_34[200], stage0_34[201], stage0_34[202], stage0_34[203]},
      {stage0_35[161]},
      {stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35]},
      {stage1_38[5],stage1_37[31],stage1_36[60],stage1_35[76],stage1_34[87]}
   );
   gpc615_5 gpc704 (
      {stage0_34[204], stage0_34[205], stage0_34[206], stage0_34[207], stage0_34[208]},
      {stage0_35[162]},
      {stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41]},
      {stage1_38[6],stage1_37[32],stage1_36[61],stage1_35[77],stage1_34[88]}
   );
   gpc615_5 gpc705 (
      {stage0_34[209], stage0_34[210], stage0_34[211], stage0_34[212], stage0_34[213]},
      {stage0_35[163]},
      {stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47]},
      {stage1_38[7],stage1_37[33],stage1_36[62],stage1_35[78],stage1_34[89]}
   );
   gpc615_5 gpc706 (
      {stage0_34[214], stage0_34[215], stage0_34[216], stage0_34[217], stage0_34[218]},
      {stage0_35[164]},
      {stage0_36[48], stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53]},
      {stage1_38[8],stage1_37[34],stage1_36[63],stage1_35[79],stage1_34[90]}
   );
   gpc615_5 gpc707 (
      {stage0_34[219], stage0_34[220], stage0_34[221], stage0_34[222], stage0_34[223]},
      {stage0_35[165]},
      {stage0_36[54], stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59]},
      {stage1_38[9],stage1_37[35],stage1_36[64],stage1_35[80],stage1_34[91]}
   );
   gpc615_5 gpc708 (
      {stage0_34[224], stage0_34[225], stage0_34[226], stage0_34[227], stage0_34[228]},
      {stage0_35[166]},
      {stage0_36[60], stage0_36[61], stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65]},
      {stage1_38[10],stage1_37[36],stage1_36[65],stage1_35[81],stage1_34[92]}
   );
   gpc615_5 gpc709 (
      {stage0_34[229], stage0_34[230], stage0_34[231], stage0_34[232], stage0_34[233]},
      {stage0_35[167]},
      {stage0_36[66], stage0_36[67], stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71]},
      {stage1_38[11],stage1_37[37],stage1_36[66],stage1_35[82],stage1_34[93]}
   );
   gpc615_5 gpc710 (
      {stage0_34[234], stage0_34[235], stage0_34[236], stage0_34[237], stage0_34[238]},
      {stage0_35[168]},
      {stage0_36[72], stage0_36[73], stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77]},
      {stage1_38[12],stage1_37[38],stage1_36[67],stage1_35[83],stage1_34[94]}
   );
   gpc615_5 gpc711 (
      {stage0_34[239], stage0_34[240], stage0_34[241], stage0_34[242], stage0_34[243]},
      {stage0_35[169]},
      {stage0_36[78], stage0_36[79], stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83]},
      {stage1_38[13],stage1_37[39],stage1_36[68],stage1_35[84],stage1_34[95]}
   );
   gpc615_5 gpc712 (
      {stage0_34[244], stage0_34[245], stage0_34[246], stage0_34[247], stage0_34[248]},
      {stage0_35[170]},
      {stage0_36[84], stage0_36[85], stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89]},
      {stage1_38[14],stage1_37[40],stage1_36[69],stage1_35[85],stage1_34[96]}
   );
   gpc615_5 gpc713 (
      {stage0_35[171], stage0_35[172], stage0_35[173], stage0_35[174], stage0_35[175]},
      {stage0_36[90]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[15],stage1_37[41],stage1_36[70],stage1_35[86]}
   );
   gpc615_5 gpc714 (
      {stage0_35[176], stage0_35[177], stage0_35[178], stage0_35[179], stage0_35[180]},
      {stage0_36[91]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[16],stage1_37[42],stage1_36[71],stage1_35[87]}
   );
   gpc615_5 gpc715 (
      {stage0_35[181], stage0_35[182], stage0_35[183], stage0_35[184], stage0_35[185]},
      {stage0_36[92]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[17],stage1_37[43],stage1_36[72],stage1_35[88]}
   );
   gpc615_5 gpc716 (
      {stage0_35[186], stage0_35[187], stage0_35[188], stage0_35[189], stage0_35[190]},
      {stage0_36[93]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[18],stage1_37[44],stage1_36[73],stage1_35[89]}
   );
   gpc615_5 gpc717 (
      {stage0_35[191], stage0_35[192], stage0_35[193], stage0_35[194], stage0_35[195]},
      {stage0_36[94]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[19],stage1_37[45],stage1_36[74],stage1_35[90]}
   );
   gpc615_5 gpc718 (
      {stage0_35[196], stage0_35[197], stage0_35[198], stage0_35[199], stage0_35[200]},
      {stage0_36[95]},
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage1_39[5],stage1_38[20],stage1_37[46],stage1_36[75],stage1_35[91]}
   );
   gpc615_5 gpc719 (
      {stage0_35[201], stage0_35[202], stage0_35[203], stage0_35[204], stage0_35[205]},
      {stage0_36[96]},
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage1_39[6],stage1_38[21],stage1_37[47],stage1_36[76],stage1_35[92]}
   );
   gpc615_5 gpc720 (
      {stage0_35[206], stage0_35[207], stage0_35[208], stage0_35[209], stage0_35[210]},
      {stage0_36[97]},
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage1_39[7],stage1_38[22],stage1_37[48],stage1_36[77],stage1_35[93]}
   );
   gpc615_5 gpc721 (
      {stage0_35[211], stage0_35[212], stage0_35[213], stage0_35[214], stage0_35[215]},
      {stage0_36[98]},
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage1_39[8],stage1_38[23],stage1_37[49],stage1_36[78],stage1_35[94]}
   );
   gpc615_5 gpc722 (
      {stage0_35[216], stage0_35[217], stage0_35[218], stage0_35[219], stage0_35[220]},
      {stage0_36[99]},
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage1_39[9],stage1_38[24],stage1_37[50],stage1_36[79],stage1_35[95]}
   );
   gpc615_5 gpc723 (
      {stage0_35[221], stage0_35[222], stage0_35[223], stage0_35[224], stage0_35[225]},
      {stage0_36[100]},
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65]},
      {stage1_39[10],stage1_38[25],stage1_37[51],stage1_36[80],stage1_35[96]}
   );
   gpc615_5 gpc724 (
      {stage0_35[226], stage0_35[227], stage0_35[228], stage0_35[229], stage0_35[230]},
      {stage0_36[101]},
      {stage0_37[66], stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71]},
      {stage1_39[11],stage1_38[26],stage1_37[52],stage1_36[81],stage1_35[97]}
   );
   gpc615_5 gpc725 (
      {stage0_35[231], stage0_35[232], stage0_35[233], stage0_35[234], stage0_35[235]},
      {stage0_36[102]},
      {stage0_37[72], stage0_37[73], stage0_37[74], stage0_37[75], stage0_37[76], stage0_37[77]},
      {stage1_39[12],stage1_38[27],stage1_37[53],stage1_36[82],stage1_35[98]}
   );
   gpc207_4 gpc726 (
      {stage0_36[103], stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107], stage0_36[108], stage0_36[109]},
      {stage0_38[0], stage0_38[1]},
      {stage1_39[13],stage1_38[28],stage1_37[54],stage1_36[83]}
   );
   gpc606_5 gpc727 (
      {stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113], stage0_36[114], stage0_36[115]},
      {stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5], stage0_38[6], stage0_38[7]},
      {stage1_40[0],stage1_39[14],stage1_38[29],stage1_37[55],stage1_36[84]}
   );
   gpc606_5 gpc728 (
      {stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119], stage0_36[120], stage0_36[121]},
      {stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11], stage0_38[12], stage0_38[13]},
      {stage1_40[1],stage1_39[15],stage1_38[30],stage1_37[56],stage1_36[85]}
   );
   gpc606_5 gpc729 (
      {stage0_36[122], stage0_36[123], stage0_36[124], stage0_36[125], stage0_36[126], stage0_36[127]},
      {stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17], stage0_38[18], stage0_38[19]},
      {stage1_40[2],stage1_39[16],stage1_38[31],stage1_37[57],stage1_36[86]}
   );
   gpc606_5 gpc730 (
      {stage0_36[128], stage0_36[129], stage0_36[130], stage0_36[131], stage0_36[132], stage0_36[133]},
      {stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23], stage0_38[24], stage0_38[25]},
      {stage1_40[3],stage1_39[17],stage1_38[32],stage1_37[58],stage1_36[87]}
   );
   gpc606_5 gpc731 (
      {stage0_36[134], stage0_36[135], stage0_36[136], stage0_36[137], stage0_36[138], stage0_36[139]},
      {stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29], stage0_38[30], stage0_38[31]},
      {stage1_40[4],stage1_39[18],stage1_38[33],stage1_37[59],stage1_36[88]}
   );
   gpc606_5 gpc732 (
      {stage0_36[140], stage0_36[141], stage0_36[142], stage0_36[143], stage0_36[144], stage0_36[145]},
      {stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35], stage0_38[36], stage0_38[37]},
      {stage1_40[5],stage1_39[19],stage1_38[34],stage1_37[60],stage1_36[89]}
   );
   gpc606_5 gpc733 (
      {stage0_36[146], stage0_36[147], stage0_36[148], stage0_36[149], stage0_36[150], stage0_36[151]},
      {stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41], stage0_38[42], stage0_38[43]},
      {stage1_40[6],stage1_39[20],stage1_38[35],stage1_37[61],stage1_36[90]}
   );
   gpc606_5 gpc734 (
      {stage0_36[152], stage0_36[153], stage0_36[154], stage0_36[155], stage0_36[156], stage0_36[157]},
      {stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47], stage0_38[48], stage0_38[49]},
      {stage1_40[7],stage1_39[21],stage1_38[36],stage1_37[62],stage1_36[91]}
   );
   gpc606_5 gpc735 (
      {stage0_36[158], stage0_36[159], stage0_36[160], stage0_36[161], stage0_36[162], stage0_36[163]},
      {stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53], stage0_38[54], stage0_38[55]},
      {stage1_40[8],stage1_39[22],stage1_38[37],stage1_37[63],stage1_36[92]}
   );
   gpc606_5 gpc736 (
      {stage0_36[164], stage0_36[165], stage0_36[166], stage0_36[167], stage0_36[168], stage0_36[169]},
      {stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59], stage0_38[60], stage0_38[61]},
      {stage1_40[9],stage1_39[23],stage1_38[38],stage1_37[64],stage1_36[93]}
   );
   gpc606_5 gpc737 (
      {stage0_36[170], stage0_36[171], stage0_36[172], stage0_36[173], stage0_36[174], stage0_36[175]},
      {stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65], stage0_38[66], stage0_38[67]},
      {stage1_40[10],stage1_39[24],stage1_38[39],stage1_37[65],stage1_36[94]}
   );
   gpc606_5 gpc738 (
      {stage0_36[176], stage0_36[177], stage0_36[178], stage0_36[179], stage0_36[180], stage0_36[181]},
      {stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71], stage0_38[72], stage0_38[73]},
      {stage1_40[11],stage1_39[25],stage1_38[40],stage1_37[66],stage1_36[95]}
   );
   gpc606_5 gpc739 (
      {stage0_36[182], stage0_36[183], stage0_36[184], stage0_36[185], stage0_36[186], stage0_36[187]},
      {stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77], stage0_38[78], stage0_38[79]},
      {stage1_40[12],stage1_39[26],stage1_38[41],stage1_37[67],stage1_36[96]}
   );
   gpc606_5 gpc740 (
      {stage0_36[188], stage0_36[189], stage0_36[190], stage0_36[191], stage0_36[192], stage0_36[193]},
      {stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83], stage0_38[84], stage0_38[85]},
      {stage1_40[13],stage1_39[27],stage1_38[42],stage1_37[68],stage1_36[97]}
   );
   gpc606_5 gpc741 (
      {stage0_36[194], stage0_36[195], stage0_36[196], stage0_36[197], stage0_36[198], stage0_36[199]},
      {stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89], stage0_38[90], stage0_38[91]},
      {stage1_40[14],stage1_39[28],stage1_38[43],stage1_37[69],stage1_36[98]}
   );
   gpc606_5 gpc742 (
      {stage0_36[200], stage0_36[201], stage0_36[202], stage0_36[203], stage0_36[204], stage0_36[205]},
      {stage0_38[92], stage0_38[93], stage0_38[94], stage0_38[95], stage0_38[96], stage0_38[97]},
      {stage1_40[15],stage1_39[29],stage1_38[44],stage1_37[70],stage1_36[99]}
   );
   gpc606_5 gpc743 (
      {stage0_36[206], stage0_36[207], stage0_36[208], stage0_36[209], stage0_36[210], stage0_36[211]},
      {stage0_38[98], stage0_38[99], stage0_38[100], stage0_38[101], stage0_38[102], stage0_38[103]},
      {stage1_40[16],stage1_39[30],stage1_38[45],stage1_37[71],stage1_36[100]}
   );
   gpc606_5 gpc744 (
      {stage0_37[78], stage0_37[79], stage0_37[80], stage0_37[81], stage0_37[82], stage0_37[83]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[17],stage1_39[31],stage1_38[46],stage1_37[72]}
   );
   gpc606_5 gpc745 (
      {stage0_37[84], stage0_37[85], stage0_37[86], stage0_37[87], stage0_37[88], stage0_37[89]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[18],stage1_39[32],stage1_38[47],stage1_37[73]}
   );
   gpc606_5 gpc746 (
      {stage0_37[90], stage0_37[91], stage0_37[92], stage0_37[93], stage0_37[94], stage0_37[95]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[19],stage1_39[33],stage1_38[48],stage1_37[74]}
   );
   gpc606_5 gpc747 (
      {stage0_37[96], stage0_37[97], stage0_37[98], stage0_37[99], stage0_37[100], stage0_37[101]},
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23]},
      {stage1_41[3],stage1_40[20],stage1_39[34],stage1_38[49],stage1_37[75]}
   );
   gpc606_5 gpc748 (
      {stage0_37[102], stage0_37[103], stage0_37[104], stage0_37[105], stage0_37[106], stage0_37[107]},
      {stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29]},
      {stage1_41[4],stage1_40[21],stage1_39[35],stage1_38[50],stage1_37[76]}
   );
   gpc606_5 gpc749 (
      {stage0_37[108], stage0_37[109], stage0_37[110], stage0_37[111], stage0_37[112], stage0_37[113]},
      {stage0_39[30], stage0_39[31], stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35]},
      {stage1_41[5],stage1_40[22],stage1_39[36],stage1_38[51],stage1_37[77]}
   );
   gpc606_5 gpc750 (
      {stage0_37[114], stage0_37[115], stage0_37[116], stage0_37[117], stage0_37[118], stage0_37[119]},
      {stage0_39[36], stage0_39[37], stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41]},
      {stage1_41[6],stage1_40[23],stage1_39[37],stage1_38[52],stage1_37[78]}
   );
   gpc606_5 gpc751 (
      {stage0_37[120], stage0_37[121], stage0_37[122], stage0_37[123], stage0_37[124], stage0_37[125]},
      {stage0_39[42], stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage1_41[7],stage1_40[24],stage1_39[38],stage1_38[53],stage1_37[79]}
   );
   gpc606_5 gpc752 (
      {stage0_37[126], stage0_37[127], stage0_37[128], stage0_37[129], stage0_37[130], stage0_37[131]},
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52], stage0_39[53]},
      {stage1_41[8],stage1_40[25],stage1_39[39],stage1_38[54],stage1_37[80]}
   );
   gpc606_5 gpc753 (
      {stage0_37[132], stage0_37[133], stage0_37[134], stage0_37[135], stage0_37[136], stage0_37[137]},
      {stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57], stage0_39[58], stage0_39[59]},
      {stage1_41[9],stage1_40[26],stage1_39[40],stage1_38[55],stage1_37[81]}
   );
   gpc606_5 gpc754 (
      {stage0_37[138], stage0_37[139], stage0_37[140], stage0_37[141], stage0_37[142], stage0_37[143]},
      {stage0_39[60], stage0_39[61], stage0_39[62], stage0_39[63], stage0_39[64], stage0_39[65]},
      {stage1_41[10],stage1_40[27],stage1_39[41],stage1_38[56],stage1_37[82]}
   );
   gpc606_5 gpc755 (
      {stage0_37[144], stage0_37[145], stage0_37[146], stage0_37[147], stage0_37[148], stage0_37[149]},
      {stage0_39[66], stage0_39[67], stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71]},
      {stage1_41[11],stage1_40[28],stage1_39[42],stage1_38[57],stage1_37[83]}
   );
   gpc606_5 gpc756 (
      {stage0_37[150], stage0_37[151], stage0_37[152], stage0_37[153], stage0_37[154], stage0_37[155]},
      {stage0_39[72], stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage1_41[12],stage1_40[29],stage1_39[43],stage1_38[58],stage1_37[84]}
   );
   gpc606_5 gpc757 (
      {stage0_37[156], stage0_37[157], stage0_37[158], stage0_37[159], stage0_37[160], stage0_37[161]},
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82], stage0_39[83]},
      {stage1_41[13],stage1_40[30],stage1_39[44],stage1_38[59],stage1_37[85]}
   );
   gpc606_5 gpc758 (
      {stage0_37[162], stage0_37[163], stage0_37[164], stage0_37[165], stage0_37[166], stage0_37[167]},
      {stage0_39[84], stage0_39[85], stage0_39[86], stage0_39[87], stage0_39[88], stage0_39[89]},
      {stage1_41[14],stage1_40[31],stage1_39[45],stage1_38[60],stage1_37[86]}
   );
   gpc606_5 gpc759 (
      {stage0_37[168], stage0_37[169], stage0_37[170], stage0_37[171], stage0_37[172], stage0_37[173]},
      {stage0_39[90], stage0_39[91], stage0_39[92], stage0_39[93], stage0_39[94], stage0_39[95]},
      {stage1_41[15],stage1_40[32],stage1_39[46],stage1_38[61],stage1_37[87]}
   );
   gpc606_5 gpc760 (
      {stage0_37[174], stage0_37[175], stage0_37[176], stage0_37[177], stage0_37[178], stage0_37[179]},
      {stage0_39[96], stage0_39[97], stage0_39[98], stage0_39[99], stage0_39[100], stage0_39[101]},
      {stage1_41[16],stage1_40[33],stage1_39[47],stage1_38[62],stage1_37[88]}
   );
   gpc606_5 gpc761 (
      {stage0_37[180], stage0_37[181], stage0_37[182], stage0_37[183], stage0_37[184], stage0_37[185]},
      {stage0_39[102], stage0_39[103], stage0_39[104], stage0_39[105], stage0_39[106], stage0_39[107]},
      {stage1_41[17],stage1_40[34],stage1_39[48],stage1_38[63],stage1_37[89]}
   );
   gpc606_5 gpc762 (
      {stage0_37[186], stage0_37[187], stage0_37[188], stage0_37[189], stage0_37[190], stage0_37[191]},
      {stage0_39[108], stage0_39[109], stage0_39[110], stage0_39[111], stage0_39[112], stage0_39[113]},
      {stage1_41[18],stage1_40[35],stage1_39[49],stage1_38[64],stage1_37[90]}
   );
   gpc606_5 gpc763 (
      {stage0_37[192], stage0_37[193], stage0_37[194], stage0_37[195], stage0_37[196], stage0_37[197]},
      {stage0_39[114], stage0_39[115], stage0_39[116], stage0_39[117], stage0_39[118], stage0_39[119]},
      {stage1_41[19],stage1_40[36],stage1_39[50],stage1_38[65],stage1_37[91]}
   );
   gpc606_5 gpc764 (
      {stage0_37[198], stage0_37[199], stage0_37[200], stage0_37[201], stage0_37[202], stage0_37[203]},
      {stage0_39[120], stage0_39[121], stage0_39[122], stage0_39[123], stage0_39[124], stage0_39[125]},
      {stage1_41[20],stage1_40[37],stage1_39[51],stage1_38[66],stage1_37[92]}
   );
   gpc606_5 gpc765 (
      {stage0_37[204], stage0_37[205], stage0_37[206], stage0_37[207], stage0_37[208], stage0_37[209]},
      {stage0_39[126], stage0_39[127], stage0_39[128], stage0_39[129], stage0_39[130], stage0_39[131]},
      {stage1_41[21],stage1_40[38],stage1_39[52],stage1_38[67],stage1_37[93]}
   );
   gpc606_5 gpc766 (
      {stage0_37[210], stage0_37[211], stage0_37[212], stage0_37[213], stage0_37[214], stage0_37[215]},
      {stage0_39[132], stage0_39[133], stage0_39[134], stage0_39[135], stage0_39[136], stage0_39[137]},
      {stage1_41[22],stage1_40[39],stage1_39[53],stage1_38[68],stage1_37[94]}
   );
   gpc606_5 gpc767 (
      {stage0_37[216], stage0_37[217], stage0_37[218], stage0_37[219], stage0_37[220], stage0_37[221]},
      {stage0_39[138], stage0_39[139], stage0_39[140], stage0_39[141], stage0_39[142], stage0_39[143]},
      {stage1_41[23],stage1_40[40],stage1_39[54],stage1_38[69],stage1_37[95]}
   );
   gpc606_5 gpc768 (
      {stage0_37[222], stage0_37[223], stage0_37[224], stage0_37[225], stage0_37[226], stage0_37[227]},
      {stage0_39[144], stage0_39[145], stage0_39[146], stage0_39[147], stage0_39[148], stage0_39[149]},
      {stage1_41[24],stage1_40[41],stage1_39[55],stage1_38[70],stage1_37[96]}
   );
   gpc606_5 gpc769 (
      {stage0_37[228], stage0_37[229], stage0_37[230], stage0_37[231], stage0_37[232], stage0_37[233]},
      {stage0_39[150], stage0_39[151], stage0_39[152], stage0_39[153], stage0_39[154], stage0_39[155]},
      {stage1_41[25],stage1_40[42],stage1_39[56],stage1_38[71],stage1_37[97]}
   );
   gpc606_5 gpc770 (
      {stage0_37[234], stage0_37[235], stage0_37[236], stage0_37[237], stage0_37[238], stage0_37[239]},
      {stage0_39[156], stage0_39[157], stage0_39[158], stage0_39[159], stage0_39[160], stage0_39[161]},
      {stage1_41[26],stage1_40[43],stage1_39[57],stage1_38[72],stage1_37[98]}
   );
   gpc606_5 gpc771 (
      {stage0_37[240], stage0_37[241], stage0_37[242], stage0_37[243], stage0_37[244], stage0_37[245]},
      {stage0_39[162], stage0_39[163], stage0_39[164], stage0_39[165], stage0_39[166], stage0_39[167]},
      {stage1_41[27],stage1_40[44],stage1_39[58],stage1_38[73],stage1_37[99]}
   );
   gpc606_5 gpc772 (
      {stage0_37[246], stage0_37[247], stage0_37[248], stage0_37[249], stage0_37[250], stage0_37[251]},
      {stage0_39[168], stage0_39[169], stage0_39[170], stage0_39[171], stage0_39[172], stage0_39[173]},
      {stage1_41[28],stage1_40[45],stage1_39[59],stage1_38[74],stage1_37[100]}
   );
   gpc615_5 gpc773 (
      {stage0_38[104], stage0_38[105], stage0_38[106], stage0_38[107], stage0_38[108]},
      {stage0_39[174]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[29],stage1_40[46],stage1_39[60],stage1_38[75]}
   );
   gpc615_5 gpc774 (
      {stage0_38[109], stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113]},
      {stage0_39[175]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[30],stage1_40[47],stage1_39[61],stage1_38[76]}
   );
   gpc615_5 gpc775 (
      {stage0_38[114], stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118]},
      {stage0_39[176]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[31],stage1_40[48],stage1_39[62],stage1_38[77]}
   );
   gpc615_5 gpc776 (
      {stage0_38[119], stage0_38[120], stage0_38[121], stage0_38[122], stage0_38[123]},
      {stage0_39[177]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[32],stage1_40[49],stage1_39[63],stage1_38[78]}
   );
   gpc615_5 gpc777 (
      {stage0_38[124], stage0_38[125], stage0_38[126], stage0_38[127], stage0_38[128]},
      {stage0_39[178]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[33],stage1_40[50],stage1_39[64],stage1_38[79]}
   );
   gpc615_5 gpc778 (
      {stage0_38[129], stage0_38[130], stage0_38[131], stage0_38[132], stage0_38[133]},
      {stage0_39[179]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[34],stage1_40[51],stage1_39[65],stage1_38[80]}
   );
   gpc615_5 gpc779 (
      {stage0_38[134], stage0_38[135], stage0_38[136], stage0_38[137], stage0_38[138]},
      {stage0_39[180]},
      {stage0_40[36], stage0_40[37], stage0_40[38], stage0_40[39], stage0_40[40], stage0_40[41]},
      {stage1_42[6],stage1_41[35],stage1_40[52],stage1_39[66],stage1_38[81]}
   );
   gpc615_5 gpc780 (
      {stage0_38[139], stage0_38[140], stage0_38[141], stage0_38[142], stage0_38[143]},
      {stage0_39[181]},
      {stage0_40[42], stage0_40[43], stage0_40[44], stage0_40[45], stage0_40[46], stage0_40[47]},
      {stage1_42[7],stage1_41[36],stage1_40[53],stage1_39[67],stage1_38[82]}
   );
   gpc615_5 gpc781 (
      {stage0_38[144], stage0_38[145], stage0_38[146], stage0_38[147], stage0_38[148]},
      {stage0_39[182]},
      {stage0_40[48], stage0_40[49], stage0_40[50], stage0_40[51], stage0_40[52], stage0_40[53]},
      {stage1_42[8],stage1_41[37],stage1_40[54],stage1_39[68],stage1_38[83]}
   );
   gpc615_5 gpc782 (
      {stage0_38[149], stage0_38[150], stage0_38[151], stage0_38[152], stage0_38[153]},
      {stage0_39[183]},
      {stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57], stage0_40[58], stage0_40[59]},
      {stage1_42[9],stage1_41[38],stage1_40[55],stage1_39[69],stage1_38[84]}
   );
   gpc615_5 gpc783 (
      {stage0_38[154], stage0_38[155], stage0_38[156], stage0_38[157], stage0_38[158]},
      {stage0_39[184]},
      {stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63], stage0_40[64], stage0_40[65]},
      {stage1_42[10],stage1_41[39],stage1_40[56],stage1_39[70],stage1_38[85]}
   );
   gpc615_5 gpc784 (
      {stage0_38[159], stage0_38[160], stage0_38[161], stage0_38[162], stage0_38[163]},
      {stage0_39[185]},
      {stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69], stage0_40[70], stage0_40[71]},
      {stage1_42[11],stage1_41[40],stage1_40[57],stage1_39[71],stage1_38[86]}
   );
   gpc615_5 gpc785 (
      {stage0_38[164], stage0_38[165], stage0_38[166], stage0_38[167], stage0_38[168]},
      {stage0_39[186]},
      {stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75], stage0_40[76], stage0_40[77]},
      {stage1_42[12],stage1_41[41],stage1_40[58],stage1_39[72],stage1_38[87]}
   );
   gpc615_5 gpc786 (
      {stage0_38[169], stage0_38[170], stage0_38[171], stage0_38[172], stage0_38[173]},
      {stage0_39[187]},
      {stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81], stage0_40[82], stage0_40[83]},
      {stage1_42[13],stage1_41[42],stage1_40[59],stage1_39[73],stage1_38[88]}
   );
   gpc615_5 gpc787 (
      {stage0_38[174], stage0_38[175], stage0_38[176], stage0_38[177], stage0_38[178]},
      {stage0_39[188]},
      {stage0_40[84], stage0_40[85], stage0_40[86], stage0_40[87], stage0_40[88], stage0_40[89]},
      {stage1_42[14],stage1_41[43],stage1_40[60],stage1_39[74],stage1_38[89]}
   );
   gpc615_5 gpc788 (
      {stage0_38[179], stage0_38[180], stage0_38[181], stage0_38[182], stage0_38[183]},
      {stage0_39[189]},
      {stage0_40[90], stage0_40[91], stage0_40[92], stage0_40[93], stage0_40[94], stage0_40[95]},
      {stage1_42[15],stage1_41[44],stage1_40[61],stage1_39[75],stage1_38[90]}
   );
   gpc615_5 gpc789 (
      {stage0_38[184], stage0_38[185], stage0_38[186], stage0_38[187], stage0_38[188]},
      {stage0_39[190]},
      {stage0_40[96], stage0_40[97], stage0_40[98], stage0_40[99], stage0_40[100], stage0_40[101]},
      {stage1_42[16],stage1_41[45],stage1_40[62],stage1_39[76],stage1_38[91]}
   );
   gpc615_5 gpc790 (
      {stage0_38[189], stage0_38[190], stage0_38[191], stage0_38[192], stage0_38[193]},
      {stage0_39[191]},
      {stage0_40[102], stage0_40[103], stage0_40[104], stage0_40[105], stage0_40[106], stage0_40[107]},
      {stage1_42[17],stage1_41[46],stage1_40[63],stage1_39[77],stage1_38[92]}
   );
   gpc615_5 gpc791 (
      {stage0_38[194], stage0_38[195], stage0_38[196], stage0_38[197], stage0_38[198]},
      {stage0_39[192]},
      {stage0_40[108], stage0_40[109], stage0_40[110], stage0_40[111], stage0_40[112], stage0_40[113]},
      {stage1_42[18],stage1_41[47],stage1_40[64],stage1_39[78],stage1_38[93]}
   );
   gpc615_5 gpc792 (
      {stage0_38[199], stage0_38[200], stage0_38[201], stage0_38[202], stage0_38[203]},
      {stage0_39[193]},
      {stage0_40[114], stage0_40[115], stage0_40[116], stage0_40[117], stage0_40[118], stage0_40[119]},
      {stage1_42[19],stage1_41[48],stage1_40[65],stage1_39[79],stage1_38[94]}
   );
   gpc615_5 gpc793 (
      {stage0_38[204], stage0_38[205], stage0_38[206], stage0_38[207], stage0_38[208]},
      {stage0_39[194]},
      {stage0_40[120], stage0_40[121], stage0_40[122], stage0_40[123], stage0_40[124], stage0_40[125]},
      {stage1_42[20],stage1_41[49],stage1_40[66],stage1_39[80],stage1_38[95]}
   );
   gpc615_5 gpc794 (
      {stage0_38[209], stage0_38[210], stage0_38[211], stage0_38[212], stage0_38[213]},
      {stage0_39[195]},
      {stage0_40[126], stage0_40[127], stage0_40[128], stage0_40[129], stage0_40[130], stage0_40[131]},
      {stage1_42[21],stage1_41[50],stage1_40[67],stage1_39[81],stage1_38[96]}
   );
   gpc623_5 gpc795 (
      {stage0_38[214], stage0_38[215], stage0_38[216]},
      {stage0_39[196], stage0_39[197]},
      {stage0_40[132], stage0_40[133], stage0_40[134], stage0_40[135], stage0_40[136], stage0_40[137]},
      {stage1_42[22],stage1_41[51],stage1_40[68],stage1_39[82],stage1_38[97]}
   );
   gpc615_5 gpc796 (
      {stage0_39[198], stage0_39[199], stage0_39[200], stage0_39[201], stage0_39[202]},
      {stage0_40[138]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[23],stage1_41[52],stage1_40[69],stage1_39[83]}
   );
   gpc615_5 gpc797 (
      {stage0_39[203], stage0_39[204], stage0_39[205], stage0_39[206], stage0_39[207]},
      {stage0_40[139]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[24],stage1_41[53],stage1_40[70],stage1_39[84]}
   );
   gpc615_5 gpc798 (
      {stage0_39[208], stage0_39[209], stage0_39[210], stage0_39[211], stage0_39[212]},
      {stage0_40[140]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[25],stage1_41[54],stage1_40[71],stage1_39[85]}
   );
   gpc615_5 gpc799 (
      {stage0_39[213], stage0_39[214], stage0_39[215], stage0_39[216], stage0_39[217]},
      {stage0_40[141]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[26],stage1_41[55],stage1_40[72],stage1_39[86]}
   );
   gpc606_5 gpc800 (
      {stage0_40[142], stage0_40[143], stage0_40[144], stage0_40[145], stage0_40[146], stage0_40[147]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[4],stage1_42[27],stage1_41[56],stage1_40[73]}
   );
   gpc606_5 gpc801 (
      {stage0_40[148], stage0_40[149], stage0_40[150], stage0_40[151], stage0_40[152], stage0_40[153]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[5],stage1_42[28],stage1_41[57],stage1_40[74]}
   );
   gpc606_5 gpc802 (
      {stage0_40[154], stage0_40[155], stage0_40[156], stage0_40[157], stage0_40[158], stage0_40[159]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[6],stage1_42[29],stage1_41[58],stage1_40[75]}
   );
   gpc606_5 gpc803 (
      {stage0_40[160], stage0_40[161], stage0_40[162], stage0_40[163], stage0_40[164], stage0_40[165]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[7],stage1_42[30],stage1_41[59],stage1_40[76]}
   );
   gpc606_5 gpc804 (
      {stage0_40[166], stage0_40[167], stage0_40[168], stage0_40[169], stage0_40[170], stage0_40[171]},
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29]},
      {stage1_44[4],stage1_43[8],stage1_42[31],stage1_41[60],stage1_40[77]}
   );
   gpc606_5 gpc805 (
      {stage0_40[172], stage0_40[173], stage0_40[174], stage0_40[175], stage0_40[176], stage0_40[177]},
      {stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35]},
      {stage1_44[5],stage1_43[9],stage1_42[32],stage1_41[61],stage1_40[78]}
   );
   gpc606_5 gpc806 (
      {stage0_40[178], stage0_40[179], stage0_40[180], stage0_40[181], stage0_40[182], stage0_40[183]},
      {stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41]},
      {stage1_44[6],stage1_43[10],stage1_42[33],stage1_41[62],stage1_40[79]}
   );
   gpc606_5 gpc807 (
      {stage0_40[184], stage0_40[185], stage0_40[186], stage0_40[187], stage0_40[188], stage0_40[189]},
      {stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47]},
      {stage1_44[7],stage1_43[11],stage1_42[34],stage1_41[63],stage1_40[80]}
   );
   gpc606_5 gpc808 (
      {stage0_40[190], stage0_40[191], stage0_40[192], stage0_40[193], stage0_40[194], stage0_40[195]},
      {stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53]},
      {stage1_44[8],stage1_43[12],stage1_42[35],stage1_41[64],stage1_40[81]}
   );
   gpc606_5 gpc809 (
      {stage0_40[196], stage0_40[197], stage0_40[198], stage0_40[199], stage0_40[200], stage0_40[201]},
      {stage0_42[54], stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59]},
      {stage1_44[9],stage1_43[13],stage1_42[36],stage1_41[65],stage1_40[82]}
   );
   gpc606_5 gpc810 (
      {stage0_40[202], stage0_40[203], stage0_40[204], stage0_40[205], stage0_40[206], stage0_40[207]},
      {stage0_42[60], stage0_42[61], stage0_42[62], stage0_42[63], stage0_42[64], stage0_42[65]},
      {stage1_44[10],stage1_43[14],stage1_42[37],stage1_41[66],stage1_40[83]}
   );
   gpc606_5 gpc811 (
      {stage0_40[208], stage0_40[209], stage0_40[210], stage0_40[211], stage0_40[212], stage0_40[213]},
      {stage0_42[66], stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage1_44[11],stage1_43[15],stage1_42[38],stage1_41[67],stage1_40[84]}
   );
   gpc606_5 gpc812 (
      {stage0_40[214], stage0_40[215], stage0_40[216], stage0_40[217], stage0_40[218], stage0_40[219]},
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76], stage0_42[77]},
      {stage1_44[12],stage1_43[16],stage1_42[39],stage1_41[68],stage1_40[85]}
   );
   gpc606_5 gpc813 (
      {stage0_40[220], stage0_40[221], stage0_40[222], stage0_40[223], stage0_40[224], stage0_40[225]},
      {stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81], stage0_42[82], stage0_42[83]},
      {stage1_44[13],stage1_43[17],stage1_42[40],stage1_41[69],stage1_40[86]}
   );
   gpc606_5 gpc814 (
      {stage0_40[226], stage0_40[227], stage0_40[228], stage0_40[229], stage0_40[230], stage0_40[231]},
      {stage0_42[84], stage0_42[85], stage0_42[86], stage0_42[87], stage0_42[88], stage0_42[89]},
      {stage1_44[14],stage1_43[18],stage1_42[41],stage1_41[70],stage1_40[87]}
   );
   gpc606_5 gpc815 (
      {stage0_40[232], stage0_40[233], stage0_40[234], stage0_40[235], stage0_40[236], stage0_40[237]},
      {stage0_42[90], stage0_42[91], stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95]},
      {stage1_44[15],stage1_43[19],stage1_42[42],stage1_41[71],stage1_40[88]}
   );
   gpc606_5 gpc816 (
      {stage0_40[238], stage0_40[239], stage0_40[240], stage0_40[241], stage0_40[242], stage0_40[243]},
      {stage0_42[96], stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage1_44[16],stage1_43[20],stage1_42[43],stage1_41[72],stage1_40[89]}
   );
   gpc606_5 gpc817 (
      {stage0_40[244], stage0_40[245], stage0_40[246], stage0_40[247], stage0_40[248], stage0_40[249]},
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106], stage0_42[107]},
      {stage1_44[17],stage1_43[21],stage1_42[44],stage1_41[73],stage1_40[90]}
   );
   gpc606_5 gpc818 (
      {stage0_40[250], stage0_40[251], stage0_40[252], stage0_40[253], stage0_40[254], stage0_40[255]},
      {stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111], stage0_42[112], stage0_42[113]},
      {stage1_44[18],stage1_43[22],stage1_42[45],stage1_41[74],stage1_40[91]}
   );
   gpc606_5 gpc819 (
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[19],stage1_43[23],stage1_42[46],stage1_41[75]}
   );
   gpc606_5 gpc820 (
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[20],stage1_43[24],stage1_42[47],stage1_41[76]}
   );
   gpc606_5 gpc821 (
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[21],stage1_43[25],stage1_42[48],stage1_41[77]}
   );
   gpc606_5 gpc822 (
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage0_43[18], stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage1_45[3],stage1_44[22],stage1_43[26],stage1_42[49],stage1_41[78]}
   );
   gpc606_5 gpc823 (
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage1_45[4],stage1_44[23],stage1_43[27],stage1_42[50],stage1_41[79]}
   );
   gpc606_5 gpc824 (
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35]},
      {stage1_45[5],stage1_44[24],stage1_43[28],stage1_42[51],stage1_41[80]}
   );
   gpc606_5 gpc825 (
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39], stage0_43[40], stage0_43[41]},
      {stage1_45[6],stage1_44[25],stage1_43[29],stage1_42[52],stage1_41[81]}
   );
   gpc606_5 gpc826 (
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage0_43[42], stage0_43[43], stage0_43[44], stage0_43[45], stage0_43[46], stage0_43[47]},
      {stage1_45[7],stage1_44[26],stage1_43[30],stage1_42[53],stage1_41[82]}
   );
   gpc606_5 gpc827 (
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage0_43[48], stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage1_45[8],stage1_44[27],stage1_43[31],stage1_42[54],stage1_41[83]}
   );
   gpc606_5 gpc828 (
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58], stage0_43[59]},
      {stage1_45[9],stage1_44[28],stage1_43[32],stage1_42[55],stage1_41[84]}
   );
   gpc606_5 gpc829 (
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63], stage0_43[64], stage0_43[65]},
      {stage1_45[10],stage1_44[29],stage1_43[33],stage1_42[56],stage1_41[85]}
   );
   gpc606_5 gpc830 (
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage0_43[66], stage0_43[67], stage0_43[68], stage0_43[69], stage0_43[70], stage0_43[71]},
      {stage1_45[11],stage1_44[30],stage1_43[34],stage1_42[57],stage1_41[86]}
   );
   gpc606_5 gpc831 (
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100], stage0_41[101]},
      {stage0_43[72], stage0_43[73], stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77]},
      {stage1_45[12],stage1_44[31],stage1_43[35],stage1_42[58],stage1_41[87]}
   );
   gpc606_5 gpc832 (
      {stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105], stage0_41[106], stage0_41[107]},
      {stage0_43[78], stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage1_45[13],stage1_44[32],stage1_43[36],stage1_42[59],stage1_41[88]}
   );
   gpc606_5 gpc833 (
      {stage0_41[108], stage0_41[109], stage0_41[110], stage0_41[111], stage0_41[112], stage0_41[113]},
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88], stage0_43[89]},
      {stage1_45[14],stage1_44[33],stage1_43[37],stage1_42[60],stage1_41[89]}
   );
   gpc606_5 gpc834 (
      {stage0_41[114], stage0_41[115], stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119]},
      {stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93], stage0_43[94], stage0_43[95]},
      {stage1_45[15],stage1_44[34],stage1_43[38],stage1_42[61],stage1_41[90]}
   );
   gpc606_5 gpc835 (
      {stage0_41[120], stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage0_43[96], stage0_43[97], stage0_43[98], stage0_43[99], stage0_43[100], stage0_43[101]},
      {stage1_45[16],stage1_44[35],stage1_43[39],stage1_42[62],stage1_41[91]}
   );
   gpc606_5 gpc836 (
      {stage0_41[126], stage0_41[127], stage0_41[128], stage0_41[129], stage0_41[130], stage0_41[131]},
      {stage0_43[102], stage0_43[103], stage0_43[104], stage0_43[105], stage0_43[106], stage0_43[107]},
      {stage1_45[17],stage1_44[36],stage1_43[40],stage1_42[63],stage1_41[92]}
   );
   gpc606_5 gpc837 (
      {stage0_41[132], stage0_41[133], stage0_41[134], stage0_41[135], stage0_41[136], stage0_41[137]},
      {stage0_43[108], stage0_43[109], stage0_43[110], stage0_43[111], stage0_43[112], stage0_43[113]},
      {stage1_45[18],stage1_44[37],stage1_43[41],stage1_42[64],stage1_41[93]}
   );
   gpc606_5 gpc838 (
      {stage0_41[138], stage0_41[139], stage0_41[140], stage0_41[141], stage0_41[142], stage0_41[143]},
      {stage0_43[114], stage0_43[115], stage0_43[116], stage0_43[117], stage0_43[118], stage0_43[119]},
      {stage1_45[19],stage1_44[38],stage1_43[42],stage1_42[65],stage1_41[94]}
   );
   gpc615_5 gpc839 (
      {stage0_41[144], stage0_41[145], stage0_41[146], stage0_41[147], stage0_41[148]},
      {stage0_42[114]},
      {stage0_43[120], stage0_43[121], stage0_43[122], stage0_43[123], stage0_43[124], stage0_43[125]},
      {stage1_45[20],stage1_44[39],stage1_43[43],stage1_42[66],stage1_41[95]}
   );
   gpc615_5 gpc840 (
      {stage0_41[149], stage0_41[150], stage0_41[151], stage0_41[152], stage0_41[153]},
      {stage0_42[115]},
      {stage0_43[126], stage0_43[127], stage0_43[128], stage0_43[129], stage0_43[130], stage0_43[131]},
      {stage1_45[21],stage1_44[40],stage1_43[44],stage1_42[67],stage1_41[96]}
   );
   gpc615_5 gpc841 (
      {stage0_41[154], stage0_41[155], stage0_41[156], stage0_41[157], stage0_41[158]},
      {stage0_42[116]},
      {stage0_43[132], stage0_43[133], stage0_43[134], stage0_43[135], stage0_43[136], stage0_43[137]},
      {stage1_45[22],stage1_44[41],stage1_43[45],stage1_42[68],stage1_41[97]}
   );
   gpc615_5 gpc842 (
      {stage0_41[159], stage0_41[160], stage0_41[161], stage0_41[162], stage0_41[163]},
      {stage0_42[117]},
      {stage0_43[138], stage0_43[139], stage0_43[140], stage0_43[141], stage0_43[142], stage0_43[143]},
      {stage1_45[23],stage1_44[42],stage1_43[46],stage1_42[69],stage1_41[98]}
   );
   gpc615_5 gpc843 (
      {stage0_41[164], stage0_41[165], stage0_41[166], stage0_41[167], stage0_41[168]},
      {stage0_42[118]},
      {stage0_43[144], stage0_43[145], stage0_43[146], stage0_43[147], stage0_43[148], stage0_43[149]},
      {stage1_45[24],stage1_44[43],stage1_43[47],stage1_42[70],stage1_41[99]}
   );
   gpc615_5 gpc844 (
      {stage0_41[169], stage0_41[170], stage0_41[171], stage0_41[172], stage0_41[173]},
      {stage0_42[119]},
      {stage0_43[150], stage0_43[151], stage0_43[152], stage0_43[153], stage0_43[154], stage0_43[155]},
      {stage1_45[25],stage1_44[44],stage1_43[48],stage1_42[71],stage1_41[100]}
   );
   gpc615_5 gpc845 (
      {stage0_41[174], stage0_41[175], stage0_41[176], stage0_41[177], stage0_41[178]},
      {stage0_42[120]},
      {stage0_43[156], stage0_43[157], stage0_43[158], stage0_43[159], stage0_43[160], stage0_43[161]},
      {stage1_45[26],stage1_44[45],stage1_43[49],stage1_42[72],stage1_41[101]}
   );
   gpc615_5 gpc846 (
      {stage0_41[179], stage0_41[180], stage0_41[181], stage0_41[182], stage0_41[183]},
      {stage0_42[121]},
      {stage0_43[162], stage0_43[163], stage0_43[164], stage0_43[165], stage0_43[166], stage0_43[167]},
      {stage1_45[27],stage1_44[46],stage1_43[50],stage1_42[73],stage1_41[102]}
   );
   gpc615_5 gpc847 (
      {stage0_41[184], stage0_41[185], stage0_41[186], stage0_41[187], stage0_41[188]},
      {stage0_42[122]},
      {stage0_43[168], stage0_43[169], stage0_43[170], stage0_43[171], stage0_43[172], stage0_43[173]},
      {stage1_45[28],stage1_44[47],stage1_43[51],stage1_42[74],stage1_41[103]}
   );
   gpc615_5 gpc848 (
      {stage0_41[189], stage0_41[190], stage0_41[191], stage0_41[192], stage0_41[193]},
      {stage0_42[123]},
      {stage0_43[174], stage0_43[175], stage0_43[176], stage0_43[177], stage0_43[178], stage0_43[179]},
      {stage1_45[29],stage1_44[48],stage1_43[52],stage1_42[75],stage1_41[104]}
   );
   gpc615_5 gpc849 (
      {stage0_41[194], stage0_41[195], stage0_41[196], stage0_41[197], stage0_41[198]},
      {stage0_42[124]},
      {stage0_43[180], stage0_43[181], stage0_43[182], stage0_43[183], stage0_43[184], stage0_43[185]},
      {stage1_45[30],stage1_44[49],stage1_43[53],stage1_42[76],stage1_41[105]}
   );
   gpc615_5 gpc850 (
      {stage0_41[199], stage0_41[200], stage0_41[201], stage0_41[202], stage0_41[203]},
      {stage0_42[125]},
      {stage0_43[186], stage0_43[187], stage0_43[188], stage0_43[189], stage0_43[190], stage0_43[191]},
      {stage1_45[31],stage1_44[50],stage1_43[54],stage1_42[77],stage1_41[106]}
   );
   gpc615_5 gpc851 (
      {stage0_41[204], stage0_41[205], stage0_41[206], stage0_41[207], stage0_41[208]},
      {stage0_42[126]},
      {stage0_43[192], stage0_43[193], stage0_43[194], stage0_43[195], stage0_43[196], stage0_43[197]},
      {stage1_45[32],stage1_44[51],stage1_43[55],stage1_42[78],stage1_41[107]}
   );
   gpc615_5 gpc852 (
      {stage0_41[209], stage0_41[210], stage0_41[211], stage0_41[212], stage0_41[213]},
      {stage0_42[127]},
      {stage0_43[198], stage0_43[199], stage0_43[200], stage0_43[201], stage0_43[202], stage0_43[203]},
      {stage1_45[33],stage1_44[52],stage1_43[56],stage1_42[79],stage1_41[108]}
   );
   gpc615_5 gpc853 (
      {stage0_41[214], stage0_41[215], stage0_41[216], stage0_41[217], stage0_41[218]},
      {stage0_42[128]},
      {stage0_43[204], stage0_43[205], stage0_43[206], stage0_43[207], stage0_43[208], stage0_43[209]},
      {stage1_45[34],stage1_44[53],stage1_43[57],stage1_42[80],stage1_41[109]}
   );
   gpc615_5 gpc854 (
      {stage0_41[219], stage0_41[220], stage0_41[221], stage0_41[222], stage0_41[223]},
      {stage0_42[129]},
      {stage0_43[210], stage0_43[211], stage0_43[212], stage0_43[213], stage0_43[214], stage0_43[215]},
      {stage1_45[35],stage1_44[54],stage1_43[58],stage1_42[81],stage1_41[110]}
   );
   gpc615_5 gpc855 (
      {stage0_42[130], stage0_42[131], stage0_42[132], stage0_42[133], stage0_42[134]},
      {stage0_43[216]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[36],stage1_44[55],stage1_43[59],stage1_42[82]}
   );
   gpc615_5 gpc856 (
      {stage0_42[135], stage0_42[136], stage0_42[137], stage0_42[138], stage0_42[139]},
      {stage0_43[217]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[37],stage1_44[56],stage1_43[60],stage1_42[83]}
   );
   gpc615_5 gpc857 (
      {stage0_42[140], stage0_42[141], stage0_42[142], stage0_42[143], stage0_42[144]},
      {stage0_43[218]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[38],stage1_44[57],stage1_43[61],stage1_42[84]}
   );
   gpc615_5 gpc858 (
      {stage0_42[145], stage0_42[146], stage0_42[147], stage0_42[148], stage0_42[149]},
      {stage0_43[219]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[39],stage1_44[58],stage1_43[62],stage1_42[85]}
   );
   gpc615_5 gpc859 (
      {stage0_42[150], stage0_42[151], stage0_42[152], stage0_42[153], stage0_42[154]},
      {stage0_43[220]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[40],stage1_44[59],stage1_43[63],stage1_42[86]}
   );
   gpc615_5 gpc860 (
      {stage0_42[155], stage0_42[156], stage0_42[157], stage0_42[158], stage0_42[159]},
      {stage0_43[221]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[41],stage1_44[60],stage1_43[64],stage1_42[87]}
   );
   gpc615_5 gpc861 (
      {stage0_42[160], stage0_42[161], stage0_42[162], stage0_42[163], stage0_42[164]},
      {stage0_43[222]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[42],stage1_44[61],stage1_43[65],stage1_42[88]}
   );
   gpc615_5 gpc862 (
      {stage0_42[165], stage0_42[166], stage0_42[167], stage0_42[168], stage0_42[169]},
      {stage0_43[223]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[43],stage1_44[62],stage1_43[66],stage1_42[89]}
   );
   gpc615_5 gpc863 (
      {stage0_42[170], stage0_42[171], stage0_42[172], stage0_42[173], stage0_42[174]},
      {stage0_43[224]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[44],stage1_44[63],stage1_43[67],stage1_42[90]}
   );
   gpc615_5 gpc864 (
      {stage0_43[225], stage0_43[226], stage0_43[227], stage0_43[228], stage0_43[229]},
      {stage0_44[54]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[9],stage1_45[45],stage1_44[64],stage1_43[68]}
   );
   gpc615_5 gpc865 (
      {stage0_43[230], stage0_43[231], stage0_43[232], stage0_43[233], stage0_43[234]},
      {stage0_44[55]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[10],stage1_45[46],stage1_44[65],stage1_43[69]}
   );
   gpc615_5 gpc866 (
      {stage0_43[235], stage0_43[236], stage0_43[237], stage0_43[238], stage0_43[239]},
      {stage0_44[56]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[11],stage1_45[47],stage1_44[66],stage1_43[70]}
   );
   gpc615_5 gpc867 (
      {stage0_43[240], stage0_43[241], stage0_43[242], stage0_43[243], stage0_43[244]},
      {stage0_44[57]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[12],stage1_45[48],stage1_44[67],stage1_43[71]}
   );
   gpc615_5 gpc868 (
      {stage0_43[245], stage0_43[246], stage0_43[247], stage0_43[248], stage0_43[249]},
      {stage0_44[58]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[13],stage1_45[49],stage1_44[68],stage1_43[72]}
   );
   gpc606_5 gpc869 (
      {stage0_44[59], stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[5],stage1_46[14],stage1_45[50],stage1_44[69]}
   );
   gpc606_5 gpc870 (
      {stage0_44[65], stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[6],stage1_46[15],stage1_45[51],stage1_44[70]}
   );
   gpc606_5 gpc871 (
      {stage0_44[71], stage0_44[72], stage0_44[73], stage0_44[74], stage0_44[75], stage0_44[76]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[7],stage1_46[16],stage1_45[52],stage1_44[71]}
   );
   gpc606_5 gpc872 (
      {stage0_44[77], stage0_44[78], stage0_44[79], stage0_44[80], stage0_44[81], stage0_44[82]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[8],stage1_46[17],stage1_45[53],stage1_44[72]}
   );
   gpc606_5 gpc873 (
      {stage0_44[83], stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[9],stage1_46[18],stage1_45[54],stage1_44[73]}
   );
   gpc606_5 gpc874 (
      {stage0_44[89], stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[10],stage1_46[19],stage1_45[55],stage1_44[74]}
   );
   gpc606_5 gpc875 (
      {stage0_44[95], stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[11],stage1_46[20],stage1_45[56],stage1_44[75]}
   );
   gpc606_5 gpc876 (
      {stage0_44[101], stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106]},
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage1_48[7],stage1_47[12],stage1_46[21],stage1_45[57],stage1_44[76]}
   );
   gpc606_5 gpc877 (
      {stage0_44[107], stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112]},
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage1_48[8],stage1_47[13],stage1_46[22],stage1_45[58],stage1_44[77]}
   );
   gpc606_5 gpc878 (
      {stage0_44[113], stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118]},
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage1_48[9],stage1_47[14],stage1_46[23],stage1_45[59],stage1_44[78]}
   );
   gpc606_5 gpc879 (
      {stage0_44[119], stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124]},
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage1_48[10],stage1_47[15],stage1_46[24],stage1_45[60],stage1_44[79]}
   );
   gpc606_5 gpc880 (
      {stage0_44[125], stage0_44[126], stage0_44[127], stage0_44[128], stage0_44[129], stage0_44[130]},
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70], stage0_46[71]},
      {stage1_48[11],stage1_47[16],stage1_46[25],stage1_45[61],stage1_44[80]}
   );
   gpc606_5 gpc881 (
      {stage0_44[131], stage0_44[132], stage0_44[133], stage0_44[134], stage0_44[135], stage0_44[136]},
      {stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75], stage0_46[76], stage0_46[77]},
      {stage1_48[12],stage1_47[17],stage1_46[26],stage1_45[62],stage1_44[81]}
   );
   gpc606_5 gpc882 (
      {stage0_44[137], stage0_44[138], stage0_44[139], stage0_44[140], stage0_44[141], stage0_44[142]},
      {stage0_46[78], stage0_46[79], stage0_46[80], stage0_46[81], stage0_46[82], stage0_46[83]},
      {stage1_48[13],stage1_47[18],stage1_46[27],stage1_45[63],stage1_44[82]}
   );
   gpc606_5 gpc883 (
      {stage0_44[143], stage0_44[144], stage0_44[145], stage0_44[146], stage0_44[147], stage0_44[148]},
      {stage0_46[84], stage0_46[85], stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89]},
      {stage1_48[14],stage1_47[19],stage1_46[28],stage1_45[64],stage1_44[83]}
   );
   gpc606_5 gpc884 (
      {stage0_44[149], stage0_44[150], stage0_44[151], stage0_44[152], stage0_44[153], stage0_44[154]},
      {stage0_46[90], stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage1_48[15],stage1_47[20],stage1_46[29],stage1_45[65],stage1_44[84]}
   );
   gpc606_5 gpc885 (
      {stage0_44[155], stage0_44[156], stage0_44[157], stage0_44[158], stage0_44[159], stage0_44[160]},
      {stage0_46[96], stage0_46[97], stage0_46[98], stage0_46[99], stage0_46[100], stage0_46[101]},
      {stage1_48[16],stage1_47[21],stage1_46[30],stage1_45[66],stage1_44[85]}
   );
   gpc606_5 gpc886 (
      {stage0_44[161], stage0_44[162], stage0_44[163], stage0_44[164], stage0_44[165], stage0_44[166]},
      {stage0_46[102], stage0_46[103], stage0_46[104], stage0_46[105], stage0_46[106], stage0_46[107]},
      {stage1_48[17],stage1_47[22],stage1_46[31],stage1_45[67],stage1_44[86]}
   );
   gpc606_5 gpc887 (
      {stage0_44[167], stage0_44[168], stage0_44[169], stage0_44[170], stage0_44[171], stage0_44[172]},
      {stage0_46[108], stage0_46[109], stage0_46[110], stage0_46[111], stage0_46[112], stage0_46[113]},
      {stage1_48[18],stage1_47[23],stage1_46[32],stage1_45[68],stage1_44[87]}
   );
   gpc606_5 gpc888 (
      {stage0_44[173], stage0_44[174], stage0_44[175], stage0_44[176], stage0_44[177], stage0_44[178]},
      {stage0_46[114], stage0_46[115], stage0_46[116], stage0_46[117], stage0_46[118], stage0_46[119]},
      {stage1_48[19],stage1_47[24],stage1_46[33],stage1_45[69],stage1_44[88]}
   );
   gpc606_5 gpc889 (
      {stage0_44[179], stage0_44[180], stage0_44[181], stage0_44[182], stage0_44[183], stage0_44[184]},
      {stage0_46[120], stage0_46[121], stage0_46[122], stage0_46[123], stage0_46[124], stage0_46[125]},
      {stage1_48[20],stage1_47[25],stage1_46[34],stage1_45[70],stage1_44[89]}
   );
   gpc606_5 gpc890 (
      {stage0_44[185], stage0_44[186], stage0_44[187], stage0_44[188], stage0_44[189], stage0_44[190]},
      {stage0_46[126], stage0_46[127], stage0_46[128], stage0_46[129], stage0_46[130], stage0_46[131]},
      {stage1_48[21],stage1_47[26],stage1_46[35],stage1_45[71],stage1_44[90]}
   );
   gpc606_5 gpc891 (
      {stage0_44[191], stage0_44[192], stage0_44[193], stage0_44[194], stage0_44[195], stage0_44[196]},
      {stage0_46[132], stage0_46[133], stage0_46[134], stage0_46[135], stage0_46[136], stage0_46[137]},
      {stage1_48[22],stage1_47[27],stage1_46[36],stage1_45[72],stage1_44[91]}
   );
   gpc606_5 gpc892 (
      {stage0_44[197], stage0_44[198], stage0_44[199], stage0_44[200], stage0_44[201], stage0_44[202]},
      {stage0_46[138], stage0_46[139], stage0_46[140], stage0_46[141], stage0_46[142], stage0_46[143]},
      {stage1_48[23],stage1_47[28],stage1_46[37],stage1_45[73],stage1_44[92]}
   );
   gpc606_5 gpc893 (
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[24],stage1_47[29],stage1_46[38],stage1_45[74]}
   );
   gpc606_5 gpc894 (
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[25],stage1_47[30],stage1_46[39],stage1_45[75]}
   );
   gpc606_5 gpc895 (
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[26],stage1_47[31],stage1_46[40],stage1_45[76]}
   );
   gpc606_5 gpc896 (
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[27],stage1_47[32],stage1_46[41],stage1_45[77]}
   );
   gpc606_5 gpc897 (
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[28],stage1_47[33],stage1_46[42],stage1_45[78]}
   );
   gpc606_5 gpc898 (
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[29],stage1_47[34],stage1_46[43],stage1_45[79]}
   );
   gpc606_5 gpc899 (
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[30],stage1_47[35],stage1_46[44],stage1_45[80]}
   );
   gpc606_5 gpc900 (
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[31],stage1_47[36],stage1_46[45],stage1_45[81]}
   );
   gpc606_5 gpc901 (
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage0_47[48], stage0_47[49], stage0_47[50], stage0_47[51], stage0_47[52], stage0_47[53]},
      {stage1_49[8],stage1_48[32],stage1_47[37],stage1_46[46],stage1_45[82]}
   );
   gpc606_5 gpc902 (
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage0_47[54], stage0_47[55], stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59]},
      {stage1_49[9],stage1_48[33],stage1_47[38],stage1_46[47],stage1_45[83]}
   );
   gpc606_5 gpc903 (
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage0_47[60], stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65]},
      {stage1_49[10],stage1_48[34],stage1_47[39],stage1_46[48],stage1_45[84]}
   );
   gpc606_5 gpc904 (
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage0_47[66], stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71]},
      {stage1_49[11],stage1_48[35],stage1_47[40],stage1_46[49],stage1_45[85]}
   );
   gpc606_5 gpc905 (
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage0_47[72], stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage1_49[12],stage1_48[36],stage1_47[41],stage1_46[50],stage1_45[86]}
   );
   gpc606_5 gpc906 (
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82], stage0_47[83]},
      {stage1_49[13],stage1_48[37],stage1_47[42],stage1_46[51],stage1_45[87]}
   );
   gpc606_5 gpc907 (
      {stage0_45[114], stage0_45[115], stage0_45[116], stage0_45[117], stage0_45[118], stage0_45[119]},
      {stage0_47[84], stage0_47[85], stage0_47[86], stage0_47[87], stage0_47[88], stage0_47[89]},
      {stage1_49[14],stage1_48[38],stage1_47[43],stage1_46[52],stage1_45[88]}
   );
   gpc606_5 gpc908 (
      {stage0_45[120], stage0_45[121], stage0_45[122], stage0_45[123], stage0_45[124], stage0_45[125]},
      {stage0_47[90], stage0_47[91], stage0_47[92], stage0_47[93], stage0_47[94], stage0_47[95]},
      {stage1_49[15],stage1_48[39],stage1_47[44],stage1_46[53],stage1_45[89]}
   );
   gpc606_5 gpc909 (
      {stage0_45[126], stage0_45[127], stage0_45[128], stage0_45[129], stage0_45[130], stage0_45[131]},
      {stage0_47[96], stage0_47[97], stage0_47[98], stage0_47[99], stage0_47[100], stage0_47[101]},
      {stage1_49[16],stage1_48[40],stage1_47[45],stage1_46[54],stage1_45[90]}
   );
   gpc606_5 gpc910 (
      {stage0_45[132], stage0_45[133], stage0_45[134], stage0_45[135], stage0_45[136], stage0_45[137]},
      {stage0_47[102], stage0_47[103], stage0_47[104], stage0_47[105], stage0_47[106], stage0_47[107]},
      {stage1_49[17],stage1_48[41],stage1_47[46],stage1_46[55],stage1_45[91]}
   );
   gpc606_5 gpc911 (
      {stage0_45[138], stage0_45[139], stage0_45[140], stage0_45[141], stage0_45[142], stage0_45[143]},
      {stage0_47[108], stage0_47[109], stage0_47[110], stage0_47[111], stage0_47[112], stage0_47[113]},
      {stage1_49[18],stage1_48[42],stage1_47[47],stage1_46[56],stage1_45[92]}
   );
   gpc606_5 gpc912 (
      {stage0_45[144], stage0_45[145], stage0_45[146], stage0_45[147], stage0_45[148], stage0_45[149]},
      {stage0_47[114], stage0_47[115], stage0_47[116], stage0_47[117], stage0_47[118], stage0_47[119]},
      {stage1_49[19],stage1_48[43],stage1_47[48],stage1_46[57],stage1_45[93]}
   );
   gpc606_5 gpc913 (
      {stage0_45[150], stage0_45[151], stage0_45[152], stage0_45[153], stage0_45[154], stage0_45[155]},
      {stage0_47[120], stage0_47[121], stage0_47[122], stage0_47[123], stage0_47[124], stage0_47[125]},
      {stage1_49[20],stage1_48[44],stage1_47[49],stage1_46[58],stage1_45[94]}
   );
   gpc606_5 gpc914 (
      {stage0_45[156], stage0_45[157], stage0_45[158], stage0_45[159], stage0_45[160], stage0_45[161]},
      {stage0_47[126], stage0_47[127], stage0_47[128], stage0_47[129], stage0_47[130], stage0_47[131]},
      {stage1_49[21],stage1_48[45],stage1_47[50],stage1_46[59],stage1_45[95]}
   );
   gpc606_5 gpc915 (
      {stage0_45[162], stage0_45[163], stage0_45[164], stage0_45[165], stage0_45[166], stage0_45[167]},
      {stage0_47[132], stage0_47[133], stage0_47[134], stage0_47[135], stage0_47[136], stage0_47[137]},
      {stage1_49[22],stage1_48[46],stage1_47[51],stage1_46[60],stage1_45[96]}
   );
   gpc606_5 gpc916 (
      {stage0_45[168], stage0_45[169], stage0_45[170], stage0_45[171], stage0_45[172], stage0_45[173]},
      {stage0_47[138], stage0_47[139], stage0_47[140], stage0_47[141], stage0_47[142], stage0_47[143]},
      {stage1_49[23],stage1_48[47],stage1_47[52],stage1_46[61],stage1_45[97]}
   );
   gpc606_5 gpc917 (
      {stage0_45[174], stage0_45[175], stage0_45[176], stage0_45[177], stage0_45[178], stage0_45[179]},
      {stage0_47[144], stage0_47[145], stage0_47[146], stage0_47[147], stage0_47[148], stage0_47[149]},
      {stage1_49[24],stage1_48[48],stage1_47[53],stage1_46[62],stage1_45[98]}
   );
   gpc615_5 gpc918 (
      {stage0_45[180], stage0_45[181], stage0_45[182], stage0_45[183], stage0_45[184]},
      {stage0_46[144]},
      {stage0_47[150], stage0_47[151], stage0_47[152], stage0_47[153], stage0_47[154], stage0_47[155]},
      {stage1_49[25],stage1_48[49],stage1_47[54],stage1_46[63],stage1_45[99]}
   );
   gpc615_5 gpc919 (
      {stage0_45[185], stage0_45[186], stage0_45[187], stage0_45[188], stage0_45[189]},
      {stage0_46[145]},
      {stage0_47[156], stage0_47[157], stage0_47[158], stage0_47[159], stage0_47[160], stage0_47[161]},
      {stage1_49[26],stage1_48[50],stage1_47[55],stage1_46[64],stage1_45[100]}
   );
   gpc615_5 gpc920 (
      {stage0_45[190], stage0_45[191], stage0_45[192], stage0_45[193], stage0_45[194]},
      {stage0_46[146]},
      {stage0_47[162], stage0_47[163], stage0_47[164], stage0_47[165], stage0_47[166], stage0_47[167]},
      {stage1_49[27],stage1_48[51],stage1_47[56],stage1_46[65],stage1_45[101]}
   );
   gpc615_5 gpc921 (
      {stage0_45[195], stage0_45[196], stage0_45[197], stage0_45[198], stage0_45[199]},
      {stage0_46[147]},
      {stage0_47[168], stage0_47[169], stage0_47[170], stage0_47[171], stage0_47[172], stage0_47[173]},
      {stage1_49[28],stage1_48[52],stage1_47[57],stage1_46[66],stage1_45[102]}
   );
   gpc606_5 gpc922 (
      {stage0_46[148], stage0_46[149], stage0_46[150], stage0_46[151], stage0_46[152], stage0_46[153]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[29],stage1_48[53],stage1_47[58],stage1_46[67]}
   );
   gpc606_5 gpc923 (
      {stage0_46[154], stage0_46[155], stage0_46[156], stage0_46[157], stage0_46[158], stage0_46[159]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[30],stage1_48[54],stage1_47[59],stage1_46[68]}
   );
   gpc606_5 gpc924 (
      {stage0_46[160], stage0_46[161], stage0_46[162], stage0_46[163], stage0_46[164], stage0_46[165]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[31],stage1_48[55],stage1_47[60],stage1_46[69]}
   );
   gpc606_5 gpc925 (
      {stage0_46[166], stage0_46[167], stage0_46[168], stage0_46[169], stage0_46[170], stage0_46[171]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[32],stage1_48[56],stage1_47[61],stage1_46[70]}
   );
   gpc606_5 gpc926 (
      {stage0_46[172], stage0_46[173], stage0_46[174], stage0_46[175], stage0_46[176], stage0_46[177]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[33],stage1_48[57],stage1_47[62],stage1_46[71]}
   );
   gpc606_5 gpc927 (
      {stage0_46[178], stage0_46[179], stage0_46[180], stage0_46[181], stage0_46[182], stage0_46[183]},
      {stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35]},
      {stage1_50[5],stage1_49[34],stage1_48[58],stage1_47[63],stage1_46[72]}
   );
   gpc606_5 gpc928 (
      {stage0_46[184], stage0_46[185], stage0_46[186], stage0_46[187], stage0_46[188], stage0_46[189]},
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage1_50[6],stage1_49[35],stage1_48[59],stage1_47[64],stage1_46[73]}
   );
   gpc606_5 gpc929 (
      {stage0_46[190], stage0_46[191], stage0_46[192], stage0_46[193], stage0_46[194], stage0_46[195]},
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage1_50[7],stage1_49[36],stage1_48[60],stage1_47[65],stage1_46[74]}
   );
   gpc606_5 gpc930 (
      {stage0_46[196], stage0_46[197], stage0_46[198], stage0_46[199], stage0_46[200], stage0_46[201]},
      {stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage1_50[8],stage1_49[37],stage1_48[61],stage1_47[66],stage1_46[75]}
   );
   gpc606_5 gpc931 (
      {stage0_46[202], stage0_46[203], stage0_46[204], stage0_46[205], stage0_46[206], stage0_46[207]},
      {stage0_48[54], stage0_48[55], stage0_48[56], stage0_48[57], stage0_48[58], stage0_48[59]},
      {stage1_50[9],stage1_49[38],stage1_48[62],stage1_47[67],stage1_46[76]}
   );
   gpc606_5 gpc932 (
      {stage0_46[208], stage0_46[209], stage0_46[210], stage0_46[211], stage0_46[212], stage0_46[213]},
      {stage0_48[60], stage0_48[61], stage0_48[62], stage0_48[63], stage0_48[64], stage0_48[65]},
      {stage1_50[10],stage1_49[39],stage1_48[63],stage1_47[68],stage1_46[77]}
   );
   gpc606_5 gpc933 (
      {stage0_46[214], stage0_46[215], stage0_46[216], stage0_46[217], stage0_46[218], stage0_46[219]},
      {stage0_48[66], stage0_48[67], stage0_48[68], stage0_48[69], stage0_48[70], stage0_48[71]},
      {stage1_50[11],stage1_49[40],stage1_48[64],stage1_47[69],stage1_46[78]}
   );
   gpc606_5 gpc934 (
      {stage0_46[220], stage0_46[221], stage0_46[222], stage0_46[223], stage0_46[224], stage0_46[225]},
      {stage0_48[72], stage0_48[73], stage0_48[74], stage0_48[75], stage0_48[76], stage0_48[77]},
      {stage1_50[12],stage1_49[41],stage1_48[65],stage1_47[70],stage1_46[79]}
   );
   gpc606_5 gpc935 (
      {stage0_46[226], stage0_46[227], stage0_46[228], stage0_46[229], stage0_46[230], stage0_46[231]},
      {stage0_48[78], stage0_48[79], stage0_48[80], stage0_48[81], stage0_48[82], stage0_48[83]},
      {stage1_50[13],stage1_49[42],stage1_48[66],stage1_47[71],stage1_46[80]}
   );
   gpc615_5 gpc936 (
      {stage0_46[232], stage0_46[233], stage0_46[234], stage0_46[235], stage0_46[236]},
      {stage0_47[174]},
      {stage0_48[84], stage0_48[85], stage0_48[86], stage0_48[87], stage0_48[88], stage0_48[89]},
      {stage1_50[14],stage1_49[43],stage1_48[67],stage1_47[72],stage1_46[81]}
   );
   gpc615_5 gpc937 (
      {stage0_47[175], stage0_47[176], stage0_47[177], stage0_47[178], stage0_47[179]},
      {stage0_48[90]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[15],stage1_49[44],stage1_48[68],stage1_47[73]}
   );
   gpc615_5 gpc938 (
      {stage0_47[180], stage0_47[181], stage0_47[182], stage0_47[183], stage0_47[184]},
      {stage0_48[91]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[16],stage1_49[45],stage1_48[69],stage1_47[74]}
   );
   gpc615_5 gpc939 (
      {stage0_47[185], stage0_47[186], stage0_47[187], stage0_47[188], stage0_47[189]},
      {stage0_48[92]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[17],stage1_49[46],stage1_48[70],stage1_47[75]}
   );
   gpc615_5 gpc940 (
      {stage0_47[190], stage0_47[191], stage0_47[192], stage0_47[193], stage0_47[194]},
      {stage0_48[93]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[18],stage1_49[47],stage1_48[71],stage1_47[76]}
   );
   gpc615_5 gpc941 (
      {stage0_47[195], stage0_47[196], stage0_47[197], stage0_47[198], stage0_47[199]},
      {stage0_48[94]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[19],stage1_49[48],stage1_48[72],stage1_47[77]}
   );
   gpc615_5 gpc942 (
      {stage0_47[200], stage0_47[201], stage0_47[202], stage0_47[203], stage0_47[204]},
      {stage0_48[95]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[20],stage1_49[49],stage1_48[73],stage1_47[78]}
   );
   gpc606_5 gpc943 (
      {stage0_48[96], stage0_48[97], stage0_48[98], stage0_48[99], stage0_48[100], stage0_48[101]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[6],stage1_50[21],stage1_49[50],stage1_48[74]}
   );
   gpc606_5 gpc944 (
      {stage0_48[102], stage0_48[103], stage0_48[104], stage0_48[105], stage0_48[106], stage0_48[107]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[7],stage1_50[22],stage1_49[51],stage1_48[75]}
   );
   gpc615_5 gpc945 (
      {stage0_48[108], stage0_48[109], stage0_48[110], stage0_48[111], stage0_48[112]},
      {stage0_49[36]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[8],stage1_50[23],stage1_49[52],stage1_48[76]}
   );
   gpc615_5 gpc946 (
      {stage0_48[113], stage0_48[114], stage0_48[115], stage0_48[116], stage0_48[117]},
      {stage0_49[37]},
      {stage0_50[18], stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage1_52[3],stage1_51[9],stage1_50[24],stage1_49[53],stage1_48[77]}
   );
   gpc615_5 gpc947 (
      {stage0_48[118], stage0_48[119], stage0_48[120], stage0_48[121], stage0_48[122]},
      {stage0_49[38]},
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage1_52[4],stage1_51[10],stage1_50[25],stage1_49[54],stage1_48[78]}
   );
   gpc615_5 gpc948 (
      {stage0_48[123], stage0_48[124], stage0_48[125], stage0_48[126], stage0_48[127]},
      {stage0_49[39]},
      {stage0_50[30], stage0_50[31], stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35]},
      {stage1_52[5],stage1_51[11],stage1_50[26],stage1_49[55],stage1_48[79]}
   );
   gpc615_5 gpc949 (
      {stage0_48[128], stage0_48[129], stage0_48[130], stage0_48[131], stage0_48[132]},
      {stage0_49[40]},
      {stage0_50[36], stage0_50[37], stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41]},
      {stage1_52[6],stage1_51[12],stage1_50[27],stage1_49[56],stage1_48[80]}
   );
   gpc615_5 gpc950 (
      {stage0_48[133], stage0_48[134], stage0_48[135], stage0_48[136], stage0_48[137]},
      {stage0_49[41]},
      {stage0_50[42], stage0_50[43], stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47]},
      {stage1_52[7],stage1_51[13],stage1_50[28],stage1_49[57],stage1_48[81]}
   );
   gpc615_5 gpc951 (
      {stage0_48[138], stage0_48[139], stage0_48[140], stage0_48[141], stage0_48[142]},
      {stage0_49[42]},
      {stage0_50[48], stage0_50[49], stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53]},
      {stage1_52[8],stage1_51[14],stage1_50[29],stage1_49[58],stage1_48[82]}
   );
   gpc615_5 gpc952 (
      {stage0_48[143], stage0_48[144], stage0_48[145], stage0_48[146], stage0_48[147]},
      {stage0_49[43]},
      {stage0_50[54], stage0_50[55], stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59]},
      {stage1_52[9],stage1_51[15],stage1_50[30],stage1_49[59],stage1_48[83]}
   );
   gpc615_5 gpc953 (
      {stage0_48[148], stage0_48[149], stage0_48[150], stage0_48[151], stage0_48[152]},
      {stage0_49[44]},
      {stage0_50[60], stage0_50[61], stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65]},
      {stage1_52[10],stage1_51[16],stage1_50[31],stage1_49[60],stage1_48[84]}
   );
   gpc615_5 gpc954 (
      {stage0_48[153], stage0_48[154], stage0_48[155], stage0_48[156], stage0_48[157]},
      {stage0_49[45]},
      {stage0_50[66], stage0_50[67], stage0_50[68], stage0_50[69], stage0_50[70], stage0_50[71]},
      {stage1_52[11],stage1_51[17],stage1_50[32],stage1_49[61],stage1_48[85]}
   );
   gpc615_5 gpc955 (
      {stage0_48[158], stage0_48[159], stage0_48[160], stage0_48[161], stage0_48[162]},
      {stage0_49[46]},
      {stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75], stage0_50[76], stage0_50[77]},
      {stage1_52[12],stage1_51[18],stage1_50[33],stage1_49[62],stage1_48[86]}
   );
   gpc615_5 gpc956 (
      {stage0_48[163], stage0_48[164], stage0_48[165], stage0_48[166], stage0_48[167]},
      {stage0_49[47]},
      {stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81], stage0_50[82], stage0_50[83]},
      {stage1_52[13],stage1_51[19],stage1_50[34],stage1_49[63],stage1_48[87]}
   );
   gpc615_5 gpc957 (
      {stage0_48[168], stage0_48[169], stage0_48[170], stage0_48[171], stage0_48[172]},
      {stage0_49[48]},
      {stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87], stage0_50[88], stage0_50[89]},
      {stage1_52[14],stage1_51[20],stage1_50[35],stage1_49[64],stage1_48[88]}
   );
   gpc615_5 gpc958 (
      {stage0_48[173], stage0_48[174], stage0_48[175], stage0_48[176], stage0_48[177]},
      {stage0_49[49]},
      {stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93], stage0_50[94], stage0_50[95]},
      {stage1_52[15],stage1_51[21],stage1_50[36],stage1_49[65],stage1_48[89]}
   );
   gpc615_5 gpc959 (
      {stage0_48[178], stage0_48[179], stage0_48[180], stage0_48[181], stage0_48[182]},
      {stage0_49[50]},
      {stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99], stage0_50[100], stage0_50[101]},
      {stage1_52[16],stage1_51[22],stage1_50[37],stage1_49[66],stage1_48[90]}
   );
   gpc615_5 gpc960 (
      {stage0_48[183], stage0_48[184], stage0_48[185], stage0_48[186], stage0_48[187]},
      {stage0_49[51]},
      {stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105], stage0_50[106], stage0_50[107]},
      {stage1_52[17],stage1_51[23],stage1_50[38],stage1_49[67],stage1_48[91]}
   );
   gpc615_5 gpc961 (
      {stage0_48[188], stage0_48[189], stage0_48[190], stage0_48[191], stage0_48[192]},
      {stage0_49[52]},
      {stage0_50[108], stage0_50[109], stage0_50[110], stage0_50[111], stage0_50[112], stage0_50[113]},
      {stage1_52[18],stage1_51[24],stage1_50[39],stage1_49[68],stage1_48[92]}
   );
   gpc615_5 gpc962 (
      {stage0_48[193], stage0_48[194], stage0_48[195], stage0_48[196], stage0_48[197]},
      {stage0_49[53]},
      {stage0_50[114], stage0_50[115], stage0_50[116], stage0_50[117], stage0_50[118], stage0_50[119]},
      {stage1_52[19],stage1_51[25],stage1_50[40],stage1_49[69],stage1_48[93]}
   );
   gpc615_5 gpc963 (
      {stage0_48[198], stage0_48[199], stage0_48[200], stage0_48[201], stage0_48[202]},
      {stage0_49[54]},
      {stage0_50[120], stage0_50[121], stage0_50[122], stage0_50[123], stage0_50[124], stage0_50[125]},
      {stage1_52[20],stage1_51[26],stage1_50[41],stage1_49[70],stage1_48[94]}
   );
   gpc615_5 gpc964 (
      {stage0_48[203], stage0_48[204], stage0_48[205], stage0_48[206], stage0_48[207]},
      {stage0_49[55]},
      {stage0_50[126], stage0_50[127], stage0_50[128], stage0_50[129], stage0_50[130], stage0_50[131]},
      {stage1_52[21],stage1_51[27],stage1_50[42],stage1_49[71],stage1_48[95]}
   );
   gpc615_5 gpc965 (
      {stage0_48[208], stage0_48[209], stage0_48[210], stage0_48[211], stage0_48[212]},
      {stage0_49[56]},
      {stage0_50[132], stage0_50[133], stage0_50[134], stage0_50[135], stage0_50[136], stage0_50[137]},
      {stage1_52[22],stage1_51[28],stage1_50[43],stage1_49[72],stage1_48[96]}
   );
   gpc615_5 gpc966 (
      {stage0_48[213], stage0_48[214], stage0_48[215], stage0_48[216], stage0_48[217]},
      {stage0_49[57]},
      {stage0_50[138], stage0_50[139], stage0_50[140], stage0_50[141], stage0_50[142], stage0_50[143]},
      {stage1_52[23],stage1_51[29],stage1_50[44],stage1_49[73],stage1_48[97]}
   );
   gpc615_5 gpc967 (
      {stage0_48[218], stage0_48[219], stage0_48[220], stage0_48[221], stage0_48[222]},
      {stage0_49[58]},
      {stage0_50[144], stage0_50[145], stage0_50[146], stage0_50[147], stage0_50[148], stage0_50[149]},
      {stage1_52[24],stage1_51[30],stage1_50[45],stage1_49[74],stage1_48[98]}
   );
   gpc615_5 gpc968 (
      {stage0_48[223], stage0_48[224], stage0_48[225], stage0_48[226], stage0_48[227]},
      {stage0_49[59]},
      {stage0_50[150], stage0_50[151], stage0_50[152], stage0_50[153], stage0_50[154], stage0_50[155]},
      {stage1_52[25],stage1_51[31],stage1_50[46],stage1_49[75],stage1_48[99]}
   );
   gpc615_5 gpc969 (
      {stage0_48[228], stage0_48[229], stage0_48[230], stage0_48[231], stage0_48[232]},
      {stage0_49[60]},
      {stage0_50[156], stage0_50[157], stage0_50[158], stage0_50[159], stage0_50[160], stage0_50[161]},
      {stage1_52[26],stage1_51[32],stage1_50[47],stage1_49[76],stage1_48[100]}
   );
   gpc615_5 gpc970 (
      {stage0_48[233], stage0_48[234], stage0_48[235], stage0_48[236], stage0_48[237]},
      {stage0_49[61]},
      {stage0_50[162], stage0_50[163], stage0_50[164], stage0_50[165], stage0_50[166], stage0_50[167]},
      {stage1_52[27],stage1_51[33],stage1_50[48],stage1_49[77],stage1_48[101]}
   );
   gpc615_5 gpc971 (
      {stage0_48[238], stage0_48[239], stage0_48[240], stage0_48[241], stage0_48[242]},
      {stage0_49[62]},
      {stage0_50[168], stage0_50[169], stage0_50[170], stage0_50[171], stage0_50[172], stage0_50[173]},
      {stage1_52[28],stage1_51[34],stage1_50[49],stage1_49[78],stage1_48[102]}
   );
   gpc615_5 gpc972 (
      {stage0_48[243], stage0_48[244], stage0_48[245], stage0_48[246], stage0_48[247]},
      {stage0_49[63]},
      {stage0_50[174], stage0_50[175], stage0_50[176], stage0_50[177], stage0_50[178], stage0_50[179]},
      {stage1_52[29],stage1_51[35],stage1_50[50],stage1_49[79],stage1_48[103]}
   );
   gpc615_5 gpc973 (
      {stage0_48[248], stage0_48[249], stage0_48[250], stage0_48[251], stage0_48[252]},
      {stage0_49[64]},
      {stage0_50[180], stage0_50[181], stage0_50[182], stage0_50[183], stage0_50[184], stage0_50[185]},
      {stage1_52[30],stage1_51[36],stage1_50[51],stage1_49[80],stage1_48[104]}
   );
   gpc606_5 gpc974 (
      {stage0_49[65], stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[31],stage1_51[37],stage1_50[52],stage1_49[81]}
   );
   gpc606_5 gpc975 (
      {stage0_49[71], stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[32],stage1_51[38],stage1_50[53],stage1_49[82]}
   );
   gpc606_5 gpc976 (
      {stage0_49[77], stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[33],stage1_51[39],stage1_50[54],stage1_49[83]}
   );
   gpc606_5 gpc977 (
      {stage0_49[83], stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[34],stage1_51[40],stage1_50[55],stage1_49[84]}
   );
   gpc606_5 gpc978 (
      {stage0_49[89], stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[35],stage1_51[41],stage1_50[56],stage1_49[85]}
   );
   gpc606_5 gpc979 (
      {stage0_49[95], stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[36],stage1_51[42],stage1_50[57],stage1_49[86]}
   );
   gpc606_5 gpc980 (
      {stage0_49[101], stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[37],stage1_51[43],stage1_50[58],stage1_49[87]}
   );
   gpc606_5 gpc981 (
      {stage0_49[107], stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[38],stage1_51[44],stage1_50[59],stage1_49[88]}
   );
   gpc606_5 gpc982 (
      {stage0_49[113], stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[39],stage1_51[45],stage1_50[60],stage1_49[89]}
   );
   gpc606_5 gpc983 (
      {stage0_49[119], stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[40],stage1_51[46],stage1_50[61],stage1_49[90]}
   );
   gpc606_5 gpc984 (
      {stage0_49[125], stage0_49[126], stage0_49[127], stage0_49[128], stage0_49[129], stage0_49[130]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[41],stage1_51[47],stage1_50[62],stage1_49[91]}
   );
   gpc606_5 gpc985 (
      {stage0_49[131], stage0_49[132], stage0_49[133], stage0_49[134], stage0_49[135], stage0_49[136]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[42],stage1_51[48],stage1_50[63],stage1_49[92]}
   );
   gpc606_5 gpc986 (
      {stage0_49[137], stage0_49[138], stage0_49[139], stage0_49[140], stage0_49[141], stage0_49[142]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[43],stage1_51[49],stage1_50[64],stage1_49[93]}
   );
   gpc606_5 gpc987 (
      {stage0_49[143], stage0_49[144], stage0_49[145], stage0_49[146], stage0_49[147], stage0_49[148]},
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage1_53[13],stage1_52[44],stage1_51[50],stage1_50[65],stage1_49[94]}
   );
   gpc606_5 gpc988 (
      {stage0_49[149], stage0_49[150], stage0_49[151], stage0_49[152], stage0_49[153], stage0_49[154]},
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage1_53[14],stage1_52[45],stage1_51[51],stage1_50[66],stage1_49[95]}
   );
   gpc606_5 gpc989 (
      {stage0_49[155], stage0_49[156], stage0_49[157], stage0_49[158], stage0_49[159], stage0_49[160]},
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage1_53[15],stage1_52[46],stage1_51[52],stage1_50[67],stage1_49[96]}
   );
   gpc606_5 gpc990 (
      {stage0_49[161], stage0_49[162], stage0_49[163], stage0_49[164], stage0_49[165], stage0_49[166]},
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage1_53[16],stage1_52[47],stage1_51[53],stage1_50[68],stage1_49[97]}
   );
   gpc606_5 gpc991 (
      {stage0_49[167], stage0_49[168], stage0_49[169], stage0_49[170], stage0_49[171], stage0_49[172]},
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage1_53[17],stage1_52[48],stage1_51[54],stage1_50[69],stage1_49[98]}
   );
   gpc606_5 gpc992 (
      {stage0_49[173], stage0_49[174], stage0_49[175], stage0_49[176], stage0_49[177], stage0_49[178]},
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage1_53[18],stage1_52[49],stage1_51[55],stage1_50[70],stage1_49[99]}
   );
   gpc606_5 gpc993 (
      {stage0_49[179], stage0_49[180], stage0_49[181], stage0_49[182], stage0_49[183], stage0_49[184]},
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage1_53[19],stage1_52[50],stage1_51[56],stage1_50[71],stage1_49[100]}
   );
   gpc606_5 gpc994 (
      {stage0_49[185], stage0_49[186], stage0_49[187], stage0_49[188], stage0_49[189], stage0_49[190]},
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage1_53[20],stage1_52[51],stage1_51[57],stage1_50[72],stage1_49[101]}
   );
   gpc606_5 gpc995 (
      {stage0_49[191], stage0_49[192], stage0_49[193], stage0_49[194], stage0_49[195], stage0_49[196]},
      {stage0_51[126], stage0_51[127], stage0_51[128], stage0_51[129], stage0_51[130], stage0_51[131]},
      {stage1_53[21],stage1_52[52],stage1_51[58],stage1_50[73],stage1_49[102]}
   );
   gpc606_5 gpc996 (
      {stage0_49[197], stage0_49[198], stage0_49[199], stage0_49[200], stage0_49[201], stage0_49[202]},
      {stage0_51[132], stage0_51[133], stage0_51[134], stage0_51[135], stage0_51[136], stage0_51[137]},
      {stage1_53[22],stage1_52[53],stage1_51[59],stage1_50[74],stage1_49[103]}
   );
   gpc606_5 gpc997 (
      {stage0_49[203], stage0_49[204], stage0_49[205], stage0_49[206], stage0_49[207], stage0_49[208]},
      {stage0_51[138], stage0_51[139], stage0_51[140], stage0_51[141], stage0_51[142], stage0_51[143]},
      {stage1_53[23],stage1_52[54],stage1_51[60],stage1_50[75],stage1_49[104]}
   );
   gpc606_5 gpc998 (
      {stage0_50[186], stage0_50[187], stage0_50[188], stage0_50[189], stage0_50[190], stage0_50[191]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[24],stage1_52[55],stage1_51[61],stage1_50[76]}
   );
   gpc606_5 gpc999 (
      {stage0_50[192], stage0_50[193], stage0_50[194], stage0_50[195], stage0_50[196], stage0_50[197]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[25],stage1_52[56],stage1_51[62],stage1_50[77]}
   );
   gpc606_5 gpc1000 (
      {stage0_50[198], stage0_50[199], stage0_50[200], stage0_50[201], stage0_50[202], stage0_50[203]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[26],stage1_52[57],stage1_51[63],stage1_50[78]}
   );
   gpc606_5 gpc1001 (
      {stage0_50[204], stage0_50[205], stage0_50[206], stage0_50[207], stage0_50[208], stage0_50[209]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[27],stage1_52[58],stage1_51[64],stage1_50[79]}
   );
   gpc606_5 gpc1002 (
      {stage0_50[210], stage0_50[211], stage0_50[212], stage0_50[213], stage0_50[214], stage0_50[215]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[28],stage1_52[59],stage1_51[65],stage1_50[80]}
   );
   gpc606_5 gpc1003 (
      {stage0_50[216], stage0_50[217], stage0_50[218], stage0_50[219], stage0_50[220], stage0_50[221]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[29],stage1_52[60],stage1_51[66],stage1_50[81]}
   );
   gpc606_5 gpc1004 (
      {stage0_50[222], stage0_50[223], stage0_50[224], stage0_50[225], stage0_50[226], stage0_50[227]},
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage1_54[6],stage1_53[30],stage1_52[61],stage1_51[67],stage1_50[82]}
   );
   gpc615_5 gpc1005 (
      {stage0_50[228], stage0_50[229], stage0_50[230], stage0_50[231], stage0_50[232]},
      {stage0_51[144]},
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage1_54[7],stage1_53[31],stage1_52[62],stage1_51[68],stage1_50[83]}
   );
   gpc615_5 gpc1006 (
      {stage0_50[233], stage0_50[234], stage0_50[235], stage0_50[236], stage0_50[237]},
      {stage0_51[145]},
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage1_54[8],stage1_53[32],stage1_52[63],stage1_51[69],stage1_50[84]}
   );
   gpc615_5 gpc1007 (
      {stage0_50[238], stage0_50[239], stage0_50[240], stage0_50[241], stage0_50[242]},
      {stage0_51[146]},
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage1_54[9],stage1_53[33],stage1_52[64],stage1_51[70],stage1_50[85]}
   );
   gpc606_5 gpc1008 (
      {stage0_51[147], stage0_51[148], stage0_51[149], stage0_51[150], stage0_51[151], stage0_51[152]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[10],stage1_53[34],stage1_52[65],stage1_51[71]}
   );
   gpc606_5 gpc1009 (
      {stage0_51[153], stage0_51[154], stage0_51[155], stage0_51[156], stage0_51[157], stage0_51[158]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[11],stage1_53[35],stage1_52[66],stage1_51[72]}
   );
   gpc606_5 gpc1010 (
      {stage0_51[159], stage0_51[160], stage0_51[161], stage0_51[162], stage0_51[163], stage0_51[164]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[12],stage1_53[36],stage1_52[67],stage1_51[73]}
   );
   gpc606_5 gpc1011 (
      {stage0_51[165], stage0_51[166], stage0_51[167], stage0_51[168], stage0_51[169], stage0_51[170]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[13],stage1_53[37],stage1_52[68],stage1_51[74]}
   );
   gpc606_5 gpc1012 (
      {stage0_51[171], stage0_51[172], stage0_51[173], stage0_51[174], stage0_51[175], stage0_51[176]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[14],stage1_53[38],stage1_52[69],stage1_51[75]}
   );
   gpc606_5 gpc1013 (
      {stage0_51[177], stage0_51[178], stage0_51[179], stage0_51[180], stage0_51[181], stage0_51[182]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[15],stage1_53[39],stage1_52[70],stage1_51[76]}
   );
   gpc606_5 gpc1014 (
      {stage0_51[183], stage0_51[184], stage0_51[185], stage0_51[186], stage0_51[187], stage0_51[188]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[16],stage1_53[40],stage1_52[71],stage1_51[77]}
   );
   gpc606_5 gpc1015 (
      {stage0_51[189], stage0_51[190], stage0_51[191], stage0_51[192], stage0_51[193], stage0_51[194]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[17],stage1_53[41],stage1_52[72],stage1_51[78]}
   );
   gpc606_5 gpc1016 (
      {stage0_51[195], stage0_51[196], stage0_51[197], stage0_51[198], stage0_51[199], stage0_51[200]},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[18],stage1_53[42],stage1_52[73],stage1_51[79]}
   );
   gpc606_5 gpc1017 (
      {stage0_51[201], stage0_51[202], stage0_51[203], stage0_51[204], stage0_51[205], stage0_51[206]},
      {stage0_53[54], stage0_53[55], stage0_53[56], stage0_53[57], stage0_53[58], stage0_53[59]},
      {stage1_55[9],stage1_54[19],stage1_53[43],stage1_52[74],stage1_51[80]}
   );
   gpc606_5 gpc1018 (
      {stage0_51[207], stage0_51[208], stage0_51[209], stage0_51[210], stage0_51[211], stage0_51[212]},
      {stage0_53[60], stage0_53[61], stage0_53[62], stage0_53[63], stage0_53[64], stage0_53[65]},
      {stage1_55[10],stage1_54[20],stage1_53[44],stage1_52[75],stage1_51[81]}
   );
   gpc606_5 gpc1019 (
      {stage0_51[213], stage0_51[214], stage0_51[215], stage0_51[216], stage0_51[217], stage0_51[218]},
      {stage0_53[66], stage0_53[67], stage0_53[68], stage0_53[69], stage0_53[70], stage0_53[71]},
      {stage1_55[11],stage1_54[21],stage1_53[45],stage1_52[76],stage1_51[82]}
   );
   gpc606_5 gpc1020 (
      {stage0_51[219], stage0_51[220], stage0_51[221], stage0_51[222], stage0_51[223], stage0_51[224]},
      {stage0_53[72], stage0_53[73], stage0_53[74], stage0_53[75], stage0_53[76], stage0_53[77]},
      {stage1_55[12],stage1_54[22],stage1_53[46],stage1_52[77],stage1_51[83]}
   );
   gpc606_5 gpc1021 (
      {stage0_51[225], stage0_51[226], stage0_51[227], stage0_51[228], stage0_51[229], stage0_51[230]},
      {stage0_53[78], stage0_53[79], stage0_53[80], stage0_53[81], stage0_53[82], stage0_53[83]},
      {stage1_55[13],stage1_54[23],stage1_53[47],stage1_52[78],stage1_51[84]}
   );
   gpc615_5 gpc1022 (
      {stage0_51[231], stage0_51[232], stage0_51[233], stage0_51[234], stage0_51[235]},
      {stage0_52[60]},
      {stage0_53[84], stage0_53[85], stage0_53[86], stage0_53[87], stage0_53[88], stage0_53[89]},
      {stage1_55[14],stage1_54[24],stage1_53[48],stage1_52[79],stage1_51[85]}
   );
   gpc606_5 gpc1023 (
      {stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65], stage0_52[66]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[15],stage1_54[25],stage1_53[49],stage1_52[80]}
   );
   gpc606_5 gpc1024 (
      {stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71], stage0_52[72]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[16],stage1_54[26],stage1_53[50],stage1_52[81]}
   );
   gpc606_5 gpc1025 (
      {stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77], stage0_52[78]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[17],stage1_54[27],stage1_53[51],stage1_52[82]}
   );
   gpc606_5 gpc1026 (
      {stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83], stage0_52[84]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[18],stage1_54[28],stage1_53[52],stage1_52[83]}
   );
   gpc606_5 gpc1027 (
      {stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89], stage0_52[90]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[19],stage1_54[29],stage1_53[53],stage1_52[84]}
   );
   gpc606_5 gpc1028 (
      {stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95], stage0_52[96]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[20],stage1_54[30],stage1_53[54],stage1_52[85]}
   );
   gpc606_5 gpc1029 (
      {stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101], stage0_52[102]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[21],stage1_54[31],stage1_53[55],stage1_52[86]}
   );
   gpc606_5 gpc1030 (
      {stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107], stage0_52[108]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[22],stage1_54[32],stage1_53[56],stage1_52[87]}
   );
   gpc606_5 gpc1031 (
      {stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113], stage0_52[114]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[23],stage1_54[33],stage1_53[57],stage1_52[88]}
   );
   gpc606_5 gpc1032 (
      {stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119], stage0_52[120]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[24],stage1_54[34],stage1_53[58],stage1_52[89]}
   );
   gpc606_5 gpc1033 (
      {stage0_52[121], stage0_52[122], stage0_52[123], stage0_52[124], stage0_52[125], stage0_52[126]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[25],stage1_54[35],stage1_53[59],stage1_52[90]}
   );
   gpc606_5 gpc1034 (
      {stage0_52[127], stage0_52[128], stage0_52[129], stage0_52[130], stage0_52[131], stage0_52[132]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[26],stage1_54[36],stage1_53[60],stage1_52[91]}
   );
   gpc606_5 gpc1035 (
      {stage0_52[133], stage0_52[134], stage0_52[135], stage0_52[136], stage0_52[137], stage0_52[138]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[27],stage1_54[37],stage1_53[61],stage1_52[92]}
   );
   gpc606_5 gpc1036 (
      {stage0_52[139], stage0_52[140], stage0_52[141], stage0_52[142], stage0_52[143], stage0_52[144]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[28],stage1_54[38],stage1_53[62],stage1_52[93]}
   );
   gpc606_5 gpc1037 (
      {stage0_52[145], stage0_52[146], stage0_52[147], stage0_52[148], stage0_52[149], stage0_52[150]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87], stage0_54[88], stage0_54[89]},
      {stage1_56[14],stage1_55[29],stage1_54[39],stage1_53[63],stage1_52[94]}
   );
   gpc606_5 gpc1038 (
      {stage0_52[151], stage0_52[152], stage0_52[153], stage0_52[154], stage0_52[155], stage0_52[156]},
      {stage0_54[90], stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95]},
      {stage1_56[15],stage1_55[30],stage1_54[40],stage1_53[64],stage1_52[95]}
   );
   gpc606_5 gpc1039 (
      {stage0_52[157], stage0_52[158], stage0_52[159], stage0_52[160], stage0_52[161], stage0_52[162]},
      {stage0_54[96], stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101]},
      {stage1_56[16],stage1_55[31],stage1_54[41],stage1_53[65],stage1_52[96]}
   );
   gpc606_5 gpc1040 (
      {stage0_52[163], stage0_52[164], stage0_52[165], stage0_52[166], stage0_52[167], stage0_52[168]},
      {stage0_54[102], stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage1_56[17],stage1_55[32],stage1_54[42],stage1_53[66],stage1_52[97]}
   );
   gpc606_5 gpc1041 (
      {stage0_52[169], stage0_52[170], stage0_52[171], stage0_52[172], stage0_52[173], stage0_52[174]},
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112], stage0_54[113]},
      {stage1_56[18],stage1_55[33],stage1_54[43],stage1_53[67],stage1_52[98]}
   );
   gpc606_5 gpc1042 (
      {stage0_52[175], stage0_52[176], stage0_52[177], stage0_52[178], stage0_52[179], stage0_52[180]},
      {stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117], stage0_54[118], stage0_54[119]},
      {stage1_56[19],stage1_55[34],stage1_54[44],stage1_53[68],stage1_52[99]}
   );
   gpc606_5 gpc1043 (
      {stage0_52[181], stage0_52[182], stage0_52[183], stage0_52[184], stage0_52[185], stage0_52[186]},
      {stage0_54[120], stage0_54[121], stage0_54[122], stage0_54[123], stage0_54[124], stage0_54[125]},
      {stage1_56[20],stage1_55[35],stage1_54[45],stage1_53[69],stage1_52[100]}
   );
   gpc606_5 gpc1044 (
      {stage0_52[187], stage0_52[188], stage0_52[189], stage0_52[190], stage0_52[191], stage0_52[192]},
      {stage0_54[126], stage0_54[127], stage0_54[128], stage0_54[129], stage0_54[130], stage0_54[131]},
      {stage1_56[21],stage1_55[36],stage1_54[46],stage1_53[70],stage1_52[101]}
   );
   gpc606_5 gpc1045 (
      {stage0_52[193], stage0_52[194], stage0_52[195], stage0_52[196], stage0_52[197], stage0_52[198]},
      {stage0_54[132], stage0_54[133], stage0_54[134], stage0_54[135], stage0_54[136], stage0_54[137]},
      {stage1_56[22],stage1_55[37],stage1_54[47],stage1_53[71],stage1_52[102]}
   );
   gpc606_5 gpc1046 (
      {stage0_52[199], stage0_52[200], stage0_52[201], stage0_52[202], stage0_52[203], stage0_52[204]},
      {stage0_54[138], stage0_54[139], stage0_54[140], stage0_54[141], stage0_54[142], stage0_54[143]},
      {stage1_56[23],stage1_55[38],stage1_54[48],stage1_53[72],stage1_52[103]}
   );
   gpc606_5 gpc1047 (
      {stage0_52[205], stage0_52[206], stage0_52[207], stage0_52[208], stage0_52[209], stage0_52[210]},
      {stage0_54[144], stage0_54[145], stage0_54[146], stage0_54[147], stage0_54[148], stage0_54[149]},
      {stage1_56[24],stage1_55[39],stage1_54[49],stage1_53[73],stage1_52[104]}
   );
   gpc606_5 gpc1048 (
      {stage0_52[211], stage0_52[212], stage0_52[213], stage0_52[214], stage0_52[215], stage0_52[216]},
      {stage0_54[150], stage0_54[151], stage0_54[152], stage0_54[153], stage0_54[154], stage0_54[155]},
      {stage1_56[25],stage1_55[40],stage1_54[50],stage1_53[74],stage1_52[105]}
   );
   gpc606_5 gpc1049 (
      {stage0_52[217], stage0_52[218], stage0_52[219], stage0_52[220], stage0_52[221], stage0_52[222]},
      {stage0_54[156], stage0_54[157], stage0_54[158], stage0_54[159], stage0_54[160], stage0_54[161]},
      {stage1_56[26],stage1_55[41],stage1_54[51],stage1_53[75],stage1_52[106]}
   );
   gpc606_5 gpc1050 (
      {stage0_53[90], stage0_53[91], stage0_53[92], stage0_53[93], stage0_53[94], stage0_53[95]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[27],stage1_55[42],stage1_54[52],stage1_53[76]}
   );
   gpc606_5 gpc1051 (
      {stage0_53[96], stage0_53[97], stage0_53[98], stage0_53[99], stage0_53[100], stage0_53[101]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[28],stage1_55[43],stage1_54[53],stage1_53[77]}
   );
   gpc606_5 gpc1052 (
      {stage0_53[102], stage0_53[103], stage0_53[104], stage0_53[105], stage0_53[106], stage0_53[107]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[29],stage1_55[44],stage1_54[54],stage1_53[78]}
   );
   gpc606_5 gpc1053 (
      {stage0_53[108], stage0_53[109], stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113]},
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage1_57[3],stage1_56[30],stage1_55[45],stage1_54[55],stage1_53[79]}
   );
   gpc606_5 gpc1054 (
      {stage0_53[114], stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage1_57[4],stage1_56[31],stage1_55[46],stage1_54[56],stage1_53[80]}
   );
   gpc606_5 gpc1055 (
      {stage0_53[120], stage0_53[121], stage0_53[122], stage0_53[123], stage0_53[124], stage0_53[125]},
      {stage0_55[30], stage0_55[31], stage0_55[32], stage0_55[33], stage0_55[34], stage0_55[35]},
      {stage1_57[5],stage1_56[32],stage1_55[47],stage1_54[57],stage1_53[81]}
   );
   gpc606_5 gpc1056 (
      {stage0_53[126], stage0_53[127], stage0_53[128], stage0_53[129], stage0_53[130], stage0_53[131]},
      {stage0_55[36], stage0_55[37], stage0_55[38], stage0_55[39], stage0_55[40], stage0_55[41]},
      {stage1_57[6],stage1_56[33],stage1_55[48],stage1_54[58],stage1_53[82]}
   );
   gpc606_5 gpc1057 (
      {stage0_53[132], stage0_53[133], stage0_53[134], stage0_53[135], stage0_53[136], stage0_53[137]},
      {stage0_55[42], stage0_55[43], stage0_55[44], stage0_55[45], stage0_55[46], stage0_55[47]},
      {stage1_57[7],stage1_56[34],stage1_55[49],stage1_54[59],stage1_53[83]}
   );
   gpc606_5 gpc1058 (
      {stage0_53[138], stage0_53[139], stage0_53[140], stage0_53[141], stage0_53[142], stage0_53[143]},
      {stage0_55[48], stage0_55[49], stage0_55[50], stage0_55[51], stage0_55[52], stage0_55[53]},
      {stage1_57[8],stage1_56[35],stage1_55[50],stage1_54[60],stage1_53[84]}
   );
   gpc606_5 gpc1059 (
      {stage0_53[144], stage0_53[145], stage0_53[146], stage0_53[147], stage0_53[148], stage0_53[149]},
      {stage0_55[54], stage0_55[55], stage0_55[56], stage0_55[57], stage0_55[58], stage0_55[59]},
      {stage1_57[9],stage1_56[36],stage1_55[51],stage1_54[61],stage1_53[85]}
   );
   gpc606_5 gpc1060 (
      {stage0_53[150], stage0_53[151], stage0_53[152], stage0_53[153], stage0_53[154], stage0_53[155]},
      {stage0_55[60], stage0_55[61], stage0_55[62], stage0_55[63], stage0_55[64], stage0_55[65]},
      {stage1_57[10],stage1_56[37],stage1_55[52],stage1_54[62],stage1_53[86]}
   );
   gpc606_5 gpc1061 (
      {stage0_53[156], stage0_53[157], stage0_53[158], stage0_53[159], stage0_53[160], stage0_53[161]},
      {stage0_55[66], stage0_55[67], stage0_55[68], stage0_55[69], stage0_55[70], stage0_55[71]},
      {stage1_57[11],stage1_56[38],stage1_55[53],stage1_54[63],stage1_53[87]}
   );
   gpc606_5 gpc1062 (
      {stage0_53[162], stage0_53[163], stage0_53[164], stage0_53[165], stage0_53[166], stage0_53[167]},
      {stage0_55[72], stage0_55[73], stage0_55[74], stage0_55[75], stage0_55[76], stage0_55[77]},
      {stage1_57[12],stage1_56[39],stage1_55[54],stage1_54[64],stage1_53[88]}
   );
   gpc606_5 gpc1063 (
      {stage0_53[168], stage0_53[169], stage0_53[170], stage0_53[171], stage0_53[172], stage0_53[173]},
      {stage0_55[78], stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83]},
      {stage1_57[13],stage1_56[40],stage1_55[55],stage1_54[65],stage1_53[89]}
   );
   gpc615_5 gpc1064 (
      {stage0_53[174], stage0_53[175], stage0_53[176], stage0_53[177], stage0_53[178]},
      {stage0_54[162]},
      {stage0_55[84], stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89]},
      {stage1_57[14],stage1_56[41],stage1_55[56],stage1_54[66],stage1_53[90]}
   );
   gpc615_5 gpc1065 (
      {stage0_53[179], stage0_53[180], stage0_53[181], stage0_53[182], stage0_53[183]},
      {stage0_54[163]},
      {stage0_55[90], stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95]},
      {stage1_57[15],stage1_56[42],stage1_55[57],stage1_54[67],stage1_53[91]}
   );
   gpc615_5 gpc1066 (
      {stage0_53[184], stage0_53[185], stage0_53[186], stage0_53[187], stage0_53[188]},
      {stage0_54[164]},
      {stage0_55[96], stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101]},
      {stage1_57[16],stage1_56[43],stage1_55[58],stage1_54[68],stage1_53[92]}
   );
   gpc615_5 gpc1067 (
      {stage0_53[189], stage0_53[190], stage0_53[191], stage0_53[192], stage0_53[193]},
      {stage0_54[165]},
      {stage0_55[102], stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage1_57[17],stage1_56[44],stage1_55[59],stage1_54[69],stage1_53[93]}
   );
   gpc615_5 gpc1068 (
      {stage0_53[194], stage0_53[195], stage0_53[196], stage0_53[197], stage0_53[198]},
      {stage0_54[166]},
      {stage0_55[108], stage0_55[109], stage0_55[110], stage0_55[111], stage0_55[112], stage0_55[113]},
      {stage1_57[18],stage1_56[45],stage1_55[60],stage1_54[70],stage1_53[94]}
   );
   gpc615_5 gpc1069 (
      {stage0_53[199], stage0_53[200], stage0_53[201], stage0_53[202], stage0_53[203]},
      {stage0_54[167]},
      {stage0_55[114], stage0_55[115], stage0_55[116], stage0_55[117], stage0_55[118], stage0_55[119]},
      {stage1_57[19],stage1_56[46],stage1_55[61],stage1_54[71],stage1_53[95]}
   );
   gpc615_5 gpc1070 (
      {stage0_53[204], stage0_53[205], stage0_53[206], stage0_53[207], stage0_53[208]},
      {stage0_54[168]},
      {stage0_55[120], stage0_55[121], stage0_55[122], stage0_55[123], stage0_55[124], stage0_55[125]},
      {stage1_57[20],stage1_56[47],stage1_55[62],stage1_54[72],stage1_53[96]}
   );
   gpc615_5 gpc1071 (
      {stage0_53[209], stage0_53[210], stage0_53[211], stage0_53[212], stage0_53[213]},
      {stage0_54[169]},
      {stage0_55[126], stage0_55[127], stage0_55[128], stage0_55[129], stage0_55[130], stage0_55[131]},
      {stage1_57[21],stage1_56[48],stage1_55[63],stage1_54[73],stage1_53[97]}
   );
   gpc615_5 gpc1072 (
      {stage0_53[214], stage0_53[215], stage0_53[216], stage0_53[217], stage0_53[218]},
      {stage0_54[170]},
      {stage0_55[132], stage0_55[133], stage0_55[134], stage0_55[135], stage0_55[136], stage0_55[137]},
      {stage1_57[22],stage1_56[49],stage1_55[64],stage1_54[74],stage1_53[98]}
   );
   gpc615_5 gpc1073 (
      {stage0_53[219], stage0_53[220], stage0_53[221], stage0_53[222], stage0_53[223]},
      {stage0_54[171]},
      {stage0_55[138], stage0_55[139], stage0_55[140], stage0_55[141], stage0_55[142], stage0_55[143]},
      {stage1_57[23],stage1_56[50],stage1_55[65],stage1_54[75],stage1_53[99]}
   );
   gpc615_5 gpc1074 (
      {stage0_53[224], stage0_53[225], stage0_53[226], stage0_53[227], stage0_53[228]},
      {stage0_54[172]},
      {stage0_55[144], stage0_55[145], stage0_55[146], stage0_55[147], stage0_55[148], stage0_55[149]},
      {stage1_57[24],stage1_56[51],stage1_55[66],stage1_54[76],stage1_53[100]}
   );
   gpc615_5 gpc1075 (
      {stage0_53[229], stage0_53[230], stage0_53[231], stage0_53[232], stage0_53[233]},
      {stage0_54[173]},
      {stage0_55[150], stage0_55[151], stage0_55[152], stage0_55[153], stage0_55[154], stage0_55[155]},
      {stage1_57[25],stage1_56[52],stage1_55[67],stage1_54[77],stage1_53[101]}
   );
   gpc615_5 gpc1076 (
      {stage0_53[234], stage0_53[235], stage0_53[236], stage0_53[237], stage0_53[238]},
      {stage0_54[174]},
      {stage0_55[156], stage0_55[157], stage0_55[158], stage0_55[159], stage0_55[160], stage0_55[161]},
      {stage1_57[26],stage1_56[53],stage1_55[68],stage1_54[78],stage1_53[102]}
   );
   gpc615_5 gpc1077 (
      {stage0_53[239], stage0_53[240], stage0_53[241], stage0_53[242], stage0_53[243]},
      {stage0_54[175]},
      {stage0_55[162], stage0_55[163], stage0_55[164], stage0_55[165], stage0_55[166], stage0_55[167]},
      {stage1_57[27],stage1_56[54],stage1_55[69],stage1_54[79],stage1_53[103]}
   );
   gpc615_5 gpc1078 (
      {stage0_53[244], stage0_53[245], stage0_53[246], stage0_53[247], stage0_53[248]},
      {stage0_54[176]},
      {stage0_55[168], stage0_55[169], stage0_55[170], stage0_55[171], stage0_55[172], stage0_55[173]},
      {stage1_57[28],stage1_56[55],stage1_55[70],stage1_54[80],stage1_53[104]}
   );
   gpc615_5 gpc1079 (
      {stage0_53[249], stage0_53[250], stage0_53[251], stage0_53[252], stage0_53[253]},
      {stage0_54[177]},
      {stage0_55[174], stage0_55[175], stage0_55[176], stage0_55[177], stage0_55[178], stage0_55[179]},
      {stage1_57[29],stage1_56[56],stage1_55[71],stage1_54[81],stage1_53[105]}
   );
   gpc606_5 gpc1080 (
      {stage0_55[180], stage0_55[181], stage0_55[182], stage0_55[183], stage0_55[184], stage0_55[185]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[0],stage1_57[30],stage1_56[57],stage1_55[72]}
   );
   gpc606_5 gpc1081 (
      {stage0_55[186], stage0_55[187], stage0_55[188], stage0_55[189], stage0_55[190], stage0_55[191]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[1],stage1_57[31],stage1_56[58],stage1_55[73]}
   );
   gpc606_5 gpc1082 (
      {stage0_55[192], stage0_55[193], stage0_55[194], stage0_55[195], stage0_55[196], stage0_55[197]},
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage1_59[2],stage1_58[2],stage1_57[32],stage1_56[59],stage1_55[74]}
   );
   gpc606_5 gpc1083 (
      {stage0_55[198], stage0_55[199], stage0_55[200], stage0_55[201], stage0_55[202], stage0_55[203]},
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage1_59[3],stage1_58[3],stage1_57[33],stage1_56[60],stage1_55[75]}
   );
   gpc606_5 gpc1084 (
      {stage0_55[204], stage0_55[205], stage0_55[206], stage0_55[207], stage0_55[208], stage0_55[209]},
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage1_59[4],stage1_58[4],stage1_57[34],stage1_56[61],stage1_55[76]}
   );
   gpc606_5 gpc1085 (
      {stage0_55[210], stage0_55[211], stage0_55[212], stage0_55[213], stage0_55[214], stage0_55[215]},
      {stage0_57[30], stage0_57[31], stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35]},
      {stage1_59[5],stage1_58[5],stage1_57[35],stage1_56[62],stage1_55[77]}
   );
   gpc606_5 gpc1086 (
      {stage0_55[216], stage0_55[217], stage0_55[218], stage0_55[219], stage0_55[220], stage0_55[221]},
      {stage0_57[36], stage0_57[37], stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41]},
      {stage1_59[6],stage1_58[6],stage1_57[36],stage1_56[63],stage1_55[78]}
   );
   gpc606_5 gpc1087 (
      {stage0_55[222], stage0_55[223], stage0_55[224], stage0_55[225], stage0_55[226], stage0_55[227]},
      {stage0_57[42], stage0_57[43], stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47]},
      {stage1_59[7],stage1_58[7],stage1_57[37],stage1_56[64],stage1_55[79]}
   );
   gpc606_5 gpc1088 (
      {stage0_55[228], stage0_55[229], stage0_55[230], stage0_55[231], stage0_55[232], stage0_55[233]},
      {stage0_57[48], stage0_57[49], stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53]},
      {stage1_59[8],stage1_58[8],stage1_57[38],stage1_56[65],stage1_55[80]}
   );
   gpc606_5 gpc1089 (
      {stage0_55[234], stage0_55[235], stage0_55[236], stage0_55[237], stage0_55[238], stage0_55[239]},
      {stage0_57[54], stage0_57[55], stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59]},
      {stage1_59[9],stage1_58[9],stage1_57[39],stage1_56[66],stage1_55[81]}
   );
   gpc615_5 gpc1090 (
      {stage0_55[240], stage0_55[241], stage0_55[242], stage0_55[243], stage0_55[244]},
      {stage0_56[0]},
      {stage0_57[60], stage0_57[61], stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65]},
      {stage1_59[10],stage1_58[10],stage1_57[40],stage1_56[67],stage1_55[82]}
   );
   gpc615_5 gpc1091 (
      {stage0_55[245], stage0_55[246], stage0_55[247], stage0_55[248], stage0_55[249]},
      {stage0_56[1]},
      {stage0_57[66], stage0_57[67], stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71]},
      {stage1_59[11],stage1_58[11],stage1_57[41],stage1_56[68],stage1_55[83]}
   );
   gpc606_5 gpc1092 (
      {stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5], stage0_56[6], stage0_56[7]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[12],stage1_58[12],stage1_57[42],stage1_56[69]}
   );
   gpc606_5 gpc1093 (
      {stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11], stage0_56[12], stage0_56[13]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[13],stage1_58[13],stage1_57[43],stage1_56[70]}
   );
   gpc606_5 gpc1094 (
      {stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17], stage0_56[18], stage0_56[19]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[14],stage1_58[14],stage1_57[44],stage1_56[71]}
   );
   gpc606_5 gpc1095 (
      {stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23], stage0_56[24], stage0_56[25]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[15],stage1_58[15],stage1_57[45],stage1_56[72]}
   );
   gpc606_5 gpc1096 (
      {stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29], stage0_56[30], stage0_56[31]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[16],stage1_58[16],stage1_57[46],stage1_56[73]}
   );
   gpc606_5 gpc1097 (
      {stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35], stage0_56[36], stage0_56[37]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[17],stage1_58[17],stage1_57[47],stage1_56[74]}
   );
   gpc606_5 gpc1098 (
      {stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41], stage0_56[42], stage0_56[43]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[18],stage1_58[18],stage1_57[48],stage1_56[75]}
   );
   gpc606_5 gpc1099 (
      {stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47], stage0_56[48], stage0_56[49]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[19],stage1_58[19],stage1_57[49],stage1_56[76]}
   );
   gpc606_5 gpc1100 (
      {stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55]},
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage1_60[8],stage1_59[20],stage1_58[20],stage1_57[50],stage1_56[77]}
   );
   gpc606_5 gpc1101 (
      {stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61]},
      {stage0_58[54], stage0_58[55], stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59]},
      {stage1_60[9],stage1_59[21],stage1_58[21],stage1_57[51],stage1_56[78]}
   );
   gpc606_5 gpc1102 (
      {stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65], stage0_56[66], stage0_56[67]},
      {stage0_58[60], stage0_58[61], stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65]},
      {stage1_60[10],stage1_59[22],stage1_58[22],stage1_57[52],stage1_56[79]}
   );
   gpc606_5 gpc1103 (
      {stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71], stage0_56[72], stage0_56[73]},
      {stage0_58[66], stage0_58[67], stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71]},
      {stage1_60[11],stage1_59[23],stage1_58[23],stage1_57[53],stage1_56[80]}
   );
   gpc606_5 gpc1104 (
      {stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77], stage0_56[78], stage0_56[79]},
      {stage0_58[72], stage0_58[73], stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77]},
      {stage1_60[12],stage1_59[24],stage1_58[24],stage1_57[54],stage1_56[81]}
   );
   gpc606_5 gpc1105 (
      {stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83], stage0_56[84], stage0_56[85]},
      {stage0_58[78], stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage1_60[13],stage1_59[25],stage1_58[25],stage1_57[55],stage1_56[82]}
   );
   gpc606_5 gpc1106 (
      {stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89], stage0_56[90], stage0_56[91]},
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88], stage0_58[89]},
      {stage1_60[14],stage1_59[26],stage1_58[26],stage1_57[56],stage1_56[83]}
   );
   gpc606_5 gpc1107 (
      {stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95], stage0_56[96], stage0_56[97]},
      {stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93], stage0_58[94], stage0_58[95]},
      {stage1_60[15],stage1_59[27],stage1_58[27],stage1_57[57],stage1_56[84]}
   );
   gpc606_5 gpc1108 (
      {stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101], stage0_56[102], stage0_56[103]},
      {stage0_58[96], stage0_58[97], stage0_58[98], stage0_58[99], stage0_58[100], stage0_58[101]},
      {stage1_60[16],stage1_59[28],stage1_58[28],stage1_57[58],stage1_56[85]}
   );
   gpc606_5 gpc1109 (
      {stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107], stage0_56[108], stage0_56[109]},
      {stage0_58[102], stage0_58[103], stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107]},
      {stage1_60[17],stage1_59[29],stage1_58[29],stage1_57[59],stage1_56[86]}
   );
   gpc606_5 gpc1110 (
      {stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113], stage0_56[114], stage0_56[115]},
      {stage0_58[108], stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage1_60[18],stage1_59[30],stage1_58[30],stage1_57[60],stage1_56[87]}
   );
   gpc606_5 gpc1111 (
      {stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119], stage0_56[120], stage0_56[121]},
      {stage0_58[114], stage0_58[115], stage0_58[116], stage0_58[117], stage0_58[118], stage0_58[119]},
      {stage1_60[19],stage1_59[31],stage1_58[31],stage1_57[61],stage1_56[88]}
   );
   gpc606_5 gpc1112 (
      {stage0_56[122], stage0_56[123], stage0_56[124], stage0_56[125], stage0_56[126], stage0_56[127]},
      {stage0_58[120], stage0_58[121], stage0_58[122], stage0_58[123], stage0_58[124], stage0_58[125]},
      {stage1_60[20],stage1_59[32],stage1_58[32],stage1_57[62],stage1_56[89]}
   );
   gpc606_5 gpc1113 (
      {stage0_56[128], stage0_56[129], stage0_56[130], stage0_56[131], stage0_56[132], stage0_56[133]},
      {stage0_58[126], stage0_58[127], stage0_58[128], stage0_58[129], stage0_58[130], stage0_58[131]},
      {stage1_60[21],stage1_59[33],stage1_58[33],stage1_57[63],stage1_56[90]}
   );
   gpc606_5 gpc1114 (
      {stage0_56[134], stage0_56[135], stage0_56[136], stage0_56[137], stage0_56[138], stage0_56[139]},
      {stage0_58[132], stage0_58[133], stage0_58[134], stage0_58[135], stage0_58[136], stage0_58[137]},
      {stage1_60[22],stage1_59[34],stage1_58[34],stage1_57[64],stage1_56[91]}
   );
   gpc606_5 gpc1115 (
      {stage0_56[140], stage0_56[141], stage0_56[142], stage0_56[143], stage0_56[144], stage0_56[145]},
      {stage0_58[138], stage0_58[139], stage0_58[140], stage0_58[141], stage0_58[142], stage0_58[143]},
      {stage1_60[23],stage1_59[35],stage1_58[35],stage1_57[65],stage1_56[92]}
   );
   gpc606_5 gpc1116 (
      {stage0_56[146], stage0_56[147], stage0_56[148], stage0_56[149], stage0_56[150], stage0_56[151]},
      {stage0_58[144], stage0_58[145], stage0_58[146], stage0_58[147], stage0_58[148], stage0_58[149]},
      {stage1_60[24],stage1_59[36],stage1_58[36],stage1_57[66],stage1_56[93]}
   );
   gpc606_5 gpc1117 (
      {stage0_56[152], stage0_56[153], stage0_56[154], stage0_56[155], stage0_56[156], stage0_56[157]},
      {stage0_58[150], stage0_58[151], stage0_58[152], stage0_58[153], stage0_58[154], stage0_58[155]},
      {stage1_60[25],stage1_59[37],stage1_58[37],stage1_57[67],stage1_56[94]}
   );
   gpc606_5 gpc1118 (
      {stage0_56[158], stage0_56[159], stage0_56[160], stage0_56[161], stage0_56[162], stage0_56[163]},
      {stage0_58[156], stage0_58[157], stage0_58[158], stage0_58[159], stage0_58[160], stage0_58[161]},
      {stage1_60[26],stage1_59[38],stage1_58[38],stage1_57[68],stage1_56[95]}
   );
   gpc606_5 gpc1119 (
      {stage0_56[164], stage0_56[165], stage0_56[166], stage0_56[167], stage0_56[168], stage0_56[169]},
      {stage0_58[162], stage0_58[163], stage0_58[164], stage0_58[165], stage0_58[166], stage0_58[167]},
      {stage1_60[27],stage1_59[39],stage1_58[39],stage1_57[69],stage1_56[96]}
   );
   gpc606_5 gpc1120 (
      {stage0_56[170], stage0_56[171], stage0_56[172], stage0_56[173], stage0_56[174], stage0_56[175]},
      {stage0_58[168], stage0_58[169], stage0_58[170], stage0_58[171], stage0_58[172], stage0_58[173]},
      {stage1_60[28],stage1_59[40],stage1_58[40],stage1_57[70],stage1_56[97]}
   );
   gpc606_5 gpc1121 (
      {stage0_57[72], stage0_57[73], stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[29],stage1_59[41],stage1_58[41],stage1_57[71]}
   );
   gpc606_5 gpc1122 (
      {stage0_57[78], stage0_57[79], stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[30],stage1_59[42],stage1_58[42],stage1_57[72]}
   );
   gpc606_5 gpc1123 (
      {stage0_57[84], stage0_57[85], stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[31],stage1_59[43],stage1_58[43],stage1_57[73]}
   );
   gpc606_5 gpc1124 (
      {stage0_57[90], stage0_57[91], stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[32],stage1_59[44],stage1_58[44],stage1_57[74]}
   );
   gpc606_5 gpc1125 (
      {stage0_57[96], stage0_57[97], stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[33],stage1_59[45],stage1_58[45],stage1_57[75]}
   );
   gpc606_5 gpc1126 (
      {stage0_57[102], stage0_57[103], stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[34],stage1_59[46],stage1_58[46],stage1_57[76]}
   );
   gpc606_5 gpc1127 (
      {stage0_57[108], stage0_57[109], stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[35],stage1_59[47],stage1_58[47],stage1_57[77]}
   );
   gpc606_5 gpc1128 (
      {stage0_57[114], stage0_57[115], stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[36],stage1_59[48],stage1_58[48],stage1_57[78]}
   );
   gpc606_5 gpc1129 (
      {stage0_57[120], stage0_57[121], stage0_57[122], stage0_57[123], stage0_57[124], stage0_57[125]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[37],stage1_59[49],stage1_58[49],stage1_57[79]}
   );
   gpc606_5 gpc1130 (
      {stage0_57[126], stage0_57[127], stage0_57[128], stage0_57[129], stage0_57[130], stage0_57[131]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[38],stage1_59[50],stage1_58[50],stage1_57[80]}
   );
   gpc606_5 gpc1131 (
      {stage0_57[132], stage0_57[133], stage0_57[134], stage0_57[135], stage0_57[136], stage0_57[137]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[39],stage1_59[51],stage1_58[51],stage1_57[81]}
   );
   gpc606_5 gpc1132 (
      {stage0_57[138], stage0_57[139], stage0_57[140], stage0_57[141], stage0_57[142], stage0_57[143]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[40],stage1_59[52],stage1_58[52],stage1_57[82]}
   );
   gpc606_5 gpc1133 (
      {stage0_57[144], stage0_57[145], stage0_57[146], stage0_57[147], stage0_57[148], stage0_57[149]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[41],stage1_59[53],stage1_58[53],stage1_57[83]}
   );
   gpc606_5 gpc1134 (
      {stage0_57[150], stage0_57[151], stage0_57[152], stage0_57[153], stage0_57[154], stage0_57[155]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[42],stage1_59[54],stage1_58[54],stage1_57[84]}
   );
   gpc606_5 gpc1135 (
      {stage0_57[156], stage0_57[157], stage0_57[158], stage0_57[159], stage0_57[160], stage0_57[161]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[43],stage1_59[55],stage1_58[55],stage1_57[85]}
   );
   gpc606_5 gpc1136 (
      {stage0_57[162], stage0_57[163], stage0_57[164], stage0_57[165], stage0_57[166], stage0_57[167]},
      {stage0_59[90], stage0_59[91], stage0_59[92], stage0_59[93], stage0_59[94], stage0_59[95]},
      {stage1_61[15],stage1_60[44],stage1_59[56],stage1_58[56],stage1_57[86]}
   );
   gpc606_5 gpc1137 (
      {stage0_57[168], stage0_57[169], stage0_57[170], stage0_57[171], stage0_57[172], stage0_57[173]},
      {stage0_59[96], stage0_59[97], stage0_59[98], stage0_59[99], stage0_59[100], stage0_59[101]},
      {stage1_61[16],stage1_60[45],stage1_59[57],stage1_58[57],stage1_57[87]}
   );
   gpc606_5 gpc1138 (
      {stage0_57[174], stage0_57[175], stage0_57[176], stage0_57[177], stage0_57[178], stage0_57[179]},
      {stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105], stage0_59[106], stage0_59[107]},
      {stage1_61[17],stage1_60[46],stage1_59[58],stage1_58[58],stage1_57[88]}
   );
   gpc606_5 gpc1139 (
      {stage0_57[180], stage0_57[181], stage0_57[182], stage0_57[183], stage0_57[184], stage0_57[185]},
      {stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111], stage0_59[112], stage0_59[113]},
      {stage1_61[18],stage1_60[47],stage1_59[59],stage1_58[59],stage1_57[89]}
   );
   gpc606_5 gpc1140 (
      {stage0_57[186], stage0_57[187], stage0_57[188], stage0_57[189], stage0_57[190], stage0_57[191]},
      {stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117], stage0_59[118], stage0_59[119]},
      {stage1_61[19],stage1_60[48],stage1_59[60],stage1_58[60],stage1_57[90]}
   );
   gpc606_5 gpc1141 (
      {stage0_57[192], stage0_57[193], stage0_57[194], stage0_57[195], stage0_57[196], stage0_57[197]},
      {stage0_59[120], stage0_59[121], stage0_59[122], stage0_59[123], stage0_59[124], stage0_59[125]},
      {stage1_61[20],stage1_60[49],stage1_59[61],stage1_58[61],stage1_57[91]}
   );
   gpc606_5 gpc1142 (
      {stage0_57[198], stage0_57[199], stage0_57[200], stage0_57[201], stage0_57[202], stage0_57[203]},
      {stage0_59[126], stage0_59[127], stage0_59[128], stage0_59[129], stage0_59[130], stage0_59[131]},
      {stage1_61[21],stage1_60[50],stage1_59[62],stage1_58[62],stage1_57[92]}
   );
   gpc606_5 gpc1143 (
      {stage0_57[204], stage0_57[205], stage0_57[206], stage0_57[207], stage0_57[208], stage0_57[209]},
      {stage0_59[132], stage0_59[133], stage0_59[134], stage0_59[135], stage0_59[136], stage0_59[137]},
      {stage1_61[22],stage1_60[51],stage1_59[63],stage1_58[63],stage1_57[93]}
   );
   gpc606_5 gpc1144 (
      {stage0_57[210], stage0_57[211], stage0_57[212], stage0_57[213], stage0_57[214], stage0_57[215]},
      {stage0_59[138], stage0_59[139], stage0_59[140], stage0_59[141], stage0_59[142], stage0_59[143]},
      {stage1_61[23],stage1_60[52],stage1_59[64],stage1_58[64],stage1_57[94]}
   );
   gpc606_5 gpc1145 (
      {stage0_57[216], stage0_57[217], stage0_57[218], stage0_57[219], stage0_57[220], stage0_57[221]},
      {stage0_59[144], stage0_59[145], stage0_59[146], stage0_59[147], stage0_59[148], stage0_59[149]},
      {stage1_61[24],stage1_60[53],stage1_59[65],stage1_58[65],stage1_57[95]}
   );
   gpc606_5 gpc1146 (
      {stage0_57[222], stage0_57[223], stage0_57[224], stage0_57[225], stage0_57[226], stage0_57[227]},
      {stage0_59[150], stage0_59[151], stage0_59[152], stage0_59[153], stage0_59[154], stage0_59[155]},
      {stage1_61[25],stage1_60[54],stage1_59[66],stage1_58[66],stage1_57[96]}
   );
   gpc615_5 gpc1147 (
      {stage0_57[228], stage0_57[229], stage0_57[230], stage0_57[231], stage0_57[232]},
      {stage0_58[174]},
      {stage0_59[156], stage0_59[157], stage0_59[158], stage0_59[159], stage0_59[160], stage0_59[161]},
      {stage1_61[26],stage1_60[55],stage1_59[67],stage1_58[67],stage1_57[97]}
   );
   gpc615_5 gpc1148 (
      {stage0_57[233], stage0_57[234], stage0_57[235], stage0_57[236], stage0_57[237]},
      {stage0_58[175]},
      {stage0_59[162], stage0_59[163], stage0_59[164], stage0_59[165], stage0_59[166], stage0_59[167]},
      {stage1_61[27],stage1_60[56],stage1_59[68],stage1_58[68],stage1_57[98]}
   );
   gpc615_5 gpc1149 (
      {stage0_57[238], stage0_57[239], stage0_57[240], stage0_57[241], stage0_57[242]},
      {stage0_58[176]},
      {stage0_59[168], stage0_59[169], stage0_59[170], stage0_59[171], stage0_59[172], stage0_59[173]},
      {stage1_61[28],stage1_60[57],stage1_59[69],stage1_58[69],stage1_57[99]}
   );
   gpc615_5 gpc1150 (
      {stage0_57[243], stage0_57[244], stage0_57[245], stage0_57[246], stage0_57[247]},
      {stage0_58[177]},
      {stage0_59[174], stage0_59[175], stage0_59[176], stage0_59[177], stage0_59[178], stage0_59[179]},
      {stage1_61[29],stage1_60[58],stage1_59[70],stage1_58[70],stage1_57[100]}
   );
   gpc615_5 gpc1151 (
      {stage0_57[248], stage0_57[249], stage0_57[250], stage0_57[251], stage0_57[252]},
      {stage0_58[178]},
      {stage0_59[180], stage0_59[181], stage0_59[182], stage0_59[183], stage0_59[184], stage0_59[185]},
      {stage1_61[30],stage1_60[59],stage1_59[71],stage1_58[71],stage1_57[101]}
   );
   gpc606_5 gpc1152 (
      {stage0_58[179], stage0_58[180], stage0_58[181], stage0_58[182], stage0_58[183], stage0_58[184]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[31],stage1_60[60],stage1_59[72],stage1_58[72]}
   );
   gpc606_5 gpc1153 (
      {stage0_58[185], stage0_58[186], stage0_58[187], stage0_58[188], stage0_58[189], stage0_58[190]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[32],stage1_60[61],stage1_59[73],stage1_58[73]}
   );
   gpc606_5 gpc1154 (
      {stage0_58[191], stage0_58[192], stage0_58[193], stage0_58[194], stage0_58[195], stage0_58[196]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[33],stage1_60[62],stage1_59[74],stage1_58[74]}
   );
   gpc606_5 gpc1155 (
      {stage0_58[197], stage0_58[198], stage0_58[199], stage0_58[200], stage0_58[201], stage0_58[202]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[34],stage1_60[63],stage1_59[75],stage1_58[75]}
   );
   gpc606_5 gpc1156 (
      {stage0_58[203], stage0_58[204], stage0_58[205], stage0_58[206], stage0_58[207], stage0_58[208]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[35],stage1_60[64],stage1_59[76],stage1_58[76]}
   );
   gpc606_5 gpc1157 (
      {stage0_58[209], stage0_58[210], stage0_58[211], stage0_58[212], stage0_58[213], stage0_58[214]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[36],stage1_60[65],stage1_59[77],stage1_58[77]}
   );
   gpc606_5 gpc1158 (
      {stage0_58[215], stage0_58[216], stage0_58[217], stage0_58[218], stage0_58[219], stage0_58[220]},
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage1_62[6],stage1_61[37],stage1_60[66],stage1_59[78],stage1_58[78]}
   );
   gpc606_5 gpc1159 (
      {stage0_58[221], stage0_58[222], stage0_58[223], stage0_58[224], stage0_58[225], stage0_58[226]},
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage1_62[7],stage1_61[38],stage1_60[67],stage1_59[79],stage1_58[79]}
   );
   gpc606_5 gpc1160 (
      {stage0_58[227], stage0_58[228], stage0_58[229], stage0_58[230], stage0_58[231], stage0_58[232]},
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage1_62[8],stage1_61[39],stage1_60[68],stage1_59[80],stage1_58[80]}
   );
   gpc606_5 gpc1161 (
      {stage0_58[233], stage0_58[234], stage0_58[235], stage0_58[236], stage0_58[237], stage0_58[238]},
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage1_62[9],stage1_61[40],stage1_60[69],stage1_59[81],stage1_58[81]}
   );
   gpc606_5 gpc1162 (
      {stage0_58[239], stage0_58[240], stage0_58[241], stage0_58[242], stage0_58[243], stage0_58[244]},
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage1_62[10],stage1_61[41],stage1_60[70],stage1_59[82],stage1_58[82]}
   );
   gpc615_5 gpc1163 (
      {stage0_58[245], stage0_58[246], stage0_58[247], stage0_58[248], stage0_58[249]},
      {stage0_59[186]},
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage1_62[11],stage1_61[42],stage1_60[71],stage1_59[83],stage1_58[83]}
   );
   gpc615_5 gpc1164 (
      {stage0_58[250], stage0_58[251], stage0_58[252], stage0_58[253], stage0_58[254]},
      {stage0_59[187]},
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage1_62[12],stage1_61[43],stage1_60[72],stage1_59[84],stage1_58[84]}
   );
   gpc1406_5 gpc1165 (
      {stage0_59[188], stage0_59[189], stage0_59[190], stage0_59[191], stage0_59[192], stage0_59[193]},
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3]},
      {stage0_62[0]},
      {stage1_63[0],stage1_62[13],stage1_61[44],stage1_60[73],stage1_59[85]}
   );
   gpc606_5 gpc1166 (
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5], stage0_62[6]},
      {stage1_64[0],stage1_63[1],stage1_62[14],stage1_61[45],stage1_60[74]}
   );
   gpc606_5 gpc1167 (
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11], stage0_62[12]},
      {stage1_64[1],stage1_63[2],stage1_62[15],stage1_61[46],stage1_60[75]}
   );
   gpc606_5 gpc1168 (
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17], stage0_62[18]},
      {stage1_64[2],stage1_63[3],stage1_62[16],stage1_61[47],stage1_60[76]}
   );
   gpc606_5 gpc1169 (
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23], stage0_62[24]},
      {stage1_64[3],stage1_63[4],stage1_62[17],stage1_61[48],stage1_60[77]}
   );
   gpc606_5 gpc1170 (
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29], stage0_62[30]},
      {stage1_64[4],stage1_63[5],stage1_62[18],stage1_61[49],stage1_60[78]}
   );
   gpc606_5 gpc1171 (
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35], stage0_62[36]},
      {stage1_64[5],stage1_63[6],stage1_62[19],stage1_61[50],stage1_60[79]}
   );
   gpc606_5 gpc1172 (
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41], stage0_62[42]},
      {stage1_64[6],stage1_63[7],stage1_62[20],stage1_61[51],stage1_60[80]}
   );
   gpc606_5 gpc1173 (
      {stage0_60[120], stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125]},
      {stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47], stage0_62[48]},
      {stage1_64[7],stage1_63[8],stage1_62[21],stage1_61[52],stage1_60[81]}
   );
   gpc606_5 gpc1174 (
      {stage0_60[126], stage0_60[127], stage0_60[128], stage0_60[129], stage0_60[130], stage0_60[131]},
      {stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53], stage0_62[54]},
      {stage1_64[8],stage1_63[9],stage1_62[22],stage1_61[53],stage1_60[82]}
   );
   gpc606_5 gpc1175 (
      {stage0_60[132], stage0_60[133], stage0_60[134], stage0_60[135], stage0_60[136], stage0_60[137]},
      {stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59], stage0_62[60]},
      {stage1_64[9],stage1_63[10],stage1_62[23],stage1_61[54],stage1_60[83]}
   );
   gpc606_5 gpc1176 (
      {stage0_60[138], stage0_60[139], stage0_60[140], stage0_60[141], stage0_60[142], stage0_60[143]},
      {stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65], stage0_62[66]},
      {stage1_64[10],stage1_63[11],stage1_62[24],stage1_61[55],stage1_60[84]}
   );
   gpc606_5 gpc1177 (
      {stage0_60[144], stage0_60[145], stage0_60[146], stage0_60[147], stage0_60[148], stage0_60[149]},
      {stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71], stage0_62[72]},
      {stage1_64[11],stage1_63[12],stage1_62[25],stage1_61[56],stage1_60[85]}
   );
   gpc606_5 gpc1178 (
      {stage0_60[150], stage0_60[151], stage0_60[152], stage0_60[153], stage0_60[154], stage0_60[155]},
      {stage0_62[73], stage0_62[74], stage0_62[75], stage0_62[76], stage0_62[77], stage0_62[78]},
      {stage1_64[12],stage1_63[13],stage1_62[26],stage1_61[57],stage1_60[86]}
   );
   gpc606_5 gpc1179 (
      {stage0_60[156], stage0_60[157], stage0_60[158], stage0_60[159], stage0_60[160], stage0_60[161]},
      {stage0_62[79], stage0_62[80], stage0_62[81], stage0_62[82], stage0_62[83], stage0_62[84]},
      {stage1_64[13],stage1_63[14],stage1_62[27],stage1_61[58],stage1_60[87]}
   );
   gpc606_5 gpc1180 (
      {stage0_60[162], stage0_60[163], stage0_60[164], stage0_60[165], stage0_60[166], stage0_60[167]},
      {stage0_62[85], stage0_62[86], stage0_62[87], stage0_62[88], stage0_62[89], stage0_62[90]},
      {stage1_64[14],stage1_63[15],stage1_62[28],stage1_61[59],stage1_60[88]}
   );
   gpc606_5 gpc1181 (
      {stage0_60[168], stage0_60[169], stage0_60[170], stage0_60[171], stage0_60[172], stage0_60[173]},
      {stage0_62[91], stage0_62[92], stage0_62[93], stage0_62[94], stage0_62[95], stage0_62[96]},
      {stage1_64[15],stage1_63[16],stage1_62[29],stage1_61[60],stage1_60[89]}
   );
   gpc606_5 gpc1182 (
      {stage0_60[174], stage0_60[175], stage0_60[176], stage0_60[177], stage0_60[178], stage0_60[179]},
      {stage0_62[97], stage0_62[98], stage0_62[99], stage0_62[100], stage0_62[101], stage0_62[102]},
      {stage1_64[16],stage1_63[17],stage1_62[30],stage1_61[61],stage1_60[90]}
   );
   gpc606_5 gpc1183 (
      {stage0_60[180], stage0_60[181], stage0_60[182], stage0_60[183], stage0_60[184], stage0_60[185]},
      {stage0_62[103], stage0_62[104], stage0_62[105], stage0_62[106], stage0_62[107], stage0_62[108]},
      {stage1_64[17],stage1_63[18],stage1_62[31],stage1_61[62],stage1_60[91]}
   );
   gpc606_5 gpc1184 (
      {stage0_60[186], stage0_60[187], stage0_60[188], stage0_60[189], stage0_60[190], stage0_60[191]},
      {stage0_62[109], stage0_62[110], stage0_62[111], stage0_62[112], stage0_62[113], stage0_62[114]},
      {stage1_64[18],stage1_63[19],stage1_62[32],stage1_61[63],stage1_60[92]}
   );
   gpc606_5 gpc1185 (
      {stage0_60[192], stage0_60[193], stage0_60[194], stage0_60[195], stage0_60[196], stage0_60[197]},
      {stage0_62[115], stage0_62[116], stage0_62[117], stage0_62[118], stage0_62[119], stage0_62[120]},
      {stage1_64[19],stage1_63[20],stage1_62[33],stage1_61[64],stage1_60[93]}
   );
   gpc606_5 gpc1186 (
      {stage0_60[198], stage0_60[199], stage0_60[200], stage0_60[201], stage0_60[202], stage0_60[203]},
      {stage0_62[121], stage0_62[122], stage0_62[123], stage0_62[124], stage0_62[125], stage0_62[126]},
      {stage1_64[20],stage1_63[21],stage1_62[34],stage1_61[65],stage1_60[94]}
   );
   gpc606_5 gpc1187 (
      {stage0_60[204], stage0_60[205], stage0_60[206], stage0_60[207], stage0_60[208], stage0_60[209]},
      {stage0_62[127], stage0_62[128], stage0_62[129], stage0_62[130], stage0_62[131], stage0_62[132]},
      {stage1_64[21],stage1_63[22],stage1_62[35],stage1_61[66],stage1_60[95]}
   );
   gpc606_5 gpc1188 (
      {stage0_61[4], stage0_61[5], stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[22],stage1_63[23],stage1_62[36],stage1_61[67]}
   );
   gpc606_5 gpc1189 (
      {stage0_61[10], stage0_61[11], stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[23],stage1_63[24],stage1_62[37],stage1_61[68]}
   );
   gpc606_5 gpc1190 (
      {stage0_61[16], stage0_61[17], stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[24],stage1_63[25],stage1_62[38],stage1_61[69]}
   );
   gpc606_5 gpc1191 (
      {stage0_61[22], stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[25],stage1_63[26],stage1_62[39],stage1_61[70]}
   );
   gpc606_5 gpc1192 (
      {stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[26],stage1_63[27],stage1_62[40],stage1_61[71]}
   );
   gpc606_5 gpc1193 (
      {stage0_61[34], stage0_61[35], stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[27],stage1_63[28],stage1_62[41],stage1_61[72]}
   );
   gpc606_5 gpc1194 (
      {stage0_61[40], stage0_61[41], stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[28],stage1_63[29],stage1_62[42],stage1_61[73]}
   );
   gpc606_5 gpc1195 (
      {stage0_61[46], stage0_61[47], stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[29],stage1_63[30],stage1_62[43],stage1_61[74]}
   );
   gpc606_5 gpc1196 (
      {stage0_61[52], stage0_61[53], stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[30],stage1_63[31],stage1_62[44],stage1_61[75]}
   );
   gpc606_5 gpc1197 (
      {stage0_61[58], stage0_61[59], stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[31],stage1_63[32],stage1_62[45],stage1_61[76]}
   );
   gpc606_5 gpc1198 (
      {stage0_61[64], stage0_61[65], stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[32],stage1_63[33],stage1_62[46],stage1_61[77]}
   );
   gpc606_5 gpc1199 (
      {stage0_61[70], stage0_61[71], stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[33],stage1_63[34],stage1_62[47],stage1_61[78]}
   );
   gpc606_5 gpc1200 (
      {stage0_61[76], stage0_61[77], stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[34],stage1_63[35],stage1_62[48],stage1_61[79]}
   );
   gpc606_5 gpc1201 (
      {stage0_61[82], stage0_61[83], stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[35],stage1_63[36],stage1_62[49],stage1_61[80]}
   );
   gpc606_5 gpc1202 (
      {stage0_61[88], stage0_61[89], stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[36],stage1_63[37],stage1_62[50],stage1_61[81]}
   );
   gpc606_5 gpc1203 (
      {stage0_61[94], stage0_61[95], stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[37],stage1_63[38],stage1_62[51],stage1_61[82]}
   );
   gpc606_5 gpc1204 (
      {stage0_61[100], stage0_61[101], stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[38],stage1_63[39],stage1_62[52],stage1_61[83]}
   );
   gpc606_5 gpc1205 (
      {stage0_61[106], stage0_61[107], stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[39],stage1_63[40],stage1_62[53],stage1_61[84]}
   );
   gpc606_5 gpc1206 (
      {stage0_61[112], stage0_61[113], stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117]},
      {stage0_63[108], stage0_63[109], stage0_63[110], stage0_63[111], stage0_63[112], stage0_63[113]},
      {stage1_65[18],stage1_64[40],stage1_63[41],stage1_62[54],stage1_61[85]}
   );
   gpc606_5 gpc1207 (
      {stage0_61[118], stage0_61[119], stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123]},
      {stage0_63[114], stage0_63[115], stage0_63[116], stage0_63[117], stage0_63[118], stage0_63[119]},
      {stage1_65[19],stage1_64[41],stage1_63[42],stage1_62[55],stage1_61[86]}
   );
   gpc606_5 gpc1208 (
      {stage0_61[124], stage0_61[125], stage0_61[126], stage0_61[127], stage0_61[128], stage0_61[129]},
      {stage0_63[120], stage0_63[121], stage0_63[122], stage0_63[123], stage0_63[124], stage0_63[125]},
      {stage1_65[20],stage1_64[42],stage1_63[43],stage1_62[56],stage1_61[87]}
   );
   gpc606_5 gpc1209 (
      {stage0_61[130], stage0_61[131], stage0_61[132], stage0_61[133], stage0_61[134], stage0_61[135]},
      {stage0_63[126], stage0_63[127], stage0_63[128], stage0_63[129], stage0_63[130], stage0_63[131]},
      {stage1_65[21],stage1_64[43],stage1_63[44],stage1_62[57],stage1_61[88]}
   );
   gpc606_5 gpc1210 (
      {stage0_61[136], stage0_61[137], stage0_61[138], stage0_61[139], stage0_61[140], stage0_61[141]},
      {stage0_63[132], stage0_63[133], stage0_63[134], stage0_63[135], stage0_63[136], stage0_63[137]},
      {stage1_65[22],stage1_64[44],stage1_63[45],stage1_62[58],stage1_61[89]}
   );
   gpc606_5 gpc1211 (
      {stage0_61[142], stage0_61[143], stage0_61[144], stage0_61[145], stage0_61[146], stage0_61[147]},
      {stage0_63[138], stage0_63[139], stage0_63[140], stage0_63[141], stage0_63[142], stage0_63[143]},
      {stage1_65[23],stage1_64[45],stage1_63[46],stage1_62[59],stage1_61[90]}
   );
   gpc606_5 gpc1212 (
      {stage0_61[148], stage0_61[149], stage0_61[150], stage0_61[151], stage0_61[152], stage0_61[153]},
      {stage0_63[144], stage0_63[145], stage0_63[146], stage0_63[147], stage0_63[148], stage0_63[149]},
      {stage1_65[24],stage1_64[46],stage1_63[47],stage1_62[60],stage1_61[91]}
   );
   gpc606_5 gpc1213 (
      {stage0_61[154], stage0_61[155], stage0_61[156], stage0_61[157], stage0_61[158], stage0_61[159]},
      {stage0_63[150], stage0_63[151], stage0_63[152], stage0_63[153], stage0_63[154], stage0_63[155]},
      {stage1_65[25],stage1_64[47],stage1_63[48],stage1_62[61],stage1_61[92]}
   );
   gpc606_5 gpc1214 (
      {stage0_61[160], stage0_61[161], stage0_61[162], stage0_61[163], stage0_61[164], stage0_61[165]},
      {stage0_63[156], stage0_63[157], stage0_63[158], stage0_63[159], stage0_63[160], stage0_63[161]},
      {stage1_65[26],stage1_64[48],stage1_63[49],stage1_62[62],stage1_61[93]}
   );
   gpc606_5 gpc1215 (
      {stage0_61[166], stage0_61[167], stage0_61[168], stage0_61[169], stage0_61[170], stage0_61[171]},
      {stage0_63[162], stage0_63[163], stage0_63[164], stage0_63[165], stage0_63[166], stage0_63[167]},
      {stage1_65[27],stage1_64[49],stage1_63[50],stage1_62[63],stage1_61[94]}
   );
   gpc606_5 gpc1216 (
      {stage0_61[172], stage0_61[173], stage0_61[174], stage0_61[175], stage0_61[176], stage0_61[177]},
      {stage0_63[168], stage0_63[169], stage0_63[170], stage0_63[171], stage0_63[172], stage0_63[173]},
      {stage1_65[28],stage1_64[50],stage1_63[51],stage1_62[64],stage1_61[95]}
   );
   gpc606_5 gpc1217 (
      {stage0_61[178], stage0_61[179], stage0_61[180], stage0_61[181], stage0_61[182], stage0_61[183]},
      {stage0_63[174], stage0_63[175], stage0_63[176], stage0_63[177], stage0_63[178], stage0_63[179]},
      {stage1_65[29],stage1_64[51],stage1_63[52],stage1_62[65],stage1_61[96]}
   );
   gpc606_5 gpc1218 (
      {stage0_61[184], stage0_61[185], stage0_61[186], stage0_61[187], stage0_61[188], stage0_61[189]},
      {stage0_63[180], stage0_63[181], stage0_63[182], stage0_63[183], stage0_63[184], stage0_63[185]},
      {stage1_65[30],stage1_64[52],stage1_63[53],stage1_62[66],stage1_61[97]}
   );
   gpc606_5 gpc1219 (
      {stage0_61[190], stage0_61[191], stage0_61[192], stage0_61[193], stage0_61[194], stage0_61[195]},
      {stage0_63[186], stage0_63[187], stage0_63[188], stage0_63[189], stage0_63[190], stage0_63[191]},
      {stage1_65[31],stage1_64[53],stage1_63[54],stage1_62[67],stage1_61[98]}
   );
   gpc606_5 gpc1220 (
      {stage0_61[196], stage0_61[197], stage0_61[198], stage0_61[199], stage0_61[200], stage0_61[201]},
      {stage0_63[192], stage0_63[193], stage0_63[194], stage0_63[195], stage0_63[196], stage0_63[197]},
      {stage1_65[32],stage1_64[54],stage1_63[55],stage1_62[68],stage1_61[99]}
   );
   gpc606_5 gpc1221 (
      {stage0_61[202], stage0_61[203], stage0_61[204], stage0_61[205], stage0_61[206], stage0_61[207]},
      {stage0_63[198], stage0_63[199], stage0_63[200], stage0_63[201], stage0_63[202], stage0_63[203]},
      {stage1_65[33],stage1_64[55],stage1_63[56],stage1_62[69],stage1_61[100]}
   );
   gpc606_5 gpc1222 (
      {stage0_61[208], stage0_61[209], stage0_61[210], stage0_61[211], stage0_61[212], stage0_61[213]},
      {stage0_63[204], stage0_63[205], stage0_63[206], stage0_63[207], stage0_63[208], stage0_63[209]},
      {stage1_65[34],stage1_64[56],stage1_63[57],stage1_62[70],stage1_61[101]}
   );
   gpc606_5 gpc1223 (
      {stage0_61[214], stage0_61[215], stage0_61[216], stage0_61[217], stage0_61[218], stage0_61[219]},
      {stage0_63[210], stage0_63[211], stage0_63[212], stage0_63[213], stage0_63[214], stage0_63[215]},
      {stage1_65[35],stage1_64[57],stage1_63[58],stage1_62[71],stage1_61[102]}
   );
   gpc606_5 gpc1224 (
      {stage0_61[220], stage0_61[221], stage0_61[222], stage0_61[223], stage0_61[224], stage0_61[225]},
      {stage0_63[216], stage0_63[217], stage0_63[218], stage0_63[219], stage0_63[220], stage0_63[221]},
      {stage1_65[36],stage1_64[58],stage1_63[59],stage1_62[72],stage1_61[103]}
   );
   gpc606_5 gpc1225 (
      {stage0_61[226], stage0_61[227], stage0_61[228], stage0_61[229], stage0_61[230], stage0_61[231]},
      {stage0_63[222], stage0_63[223], stage0_63[224], stage0_63[225], stage0_63[226], stage0_63[227]},
      {stage1_65[37],stage1_64[59],stage1_63[60],stage1_62[73],stage1_61[104]}
   );
   gpc606_5 gpc1226 (
      {stage0_61[232], stage0_61[233], stage0_61[234], stage0_61[235], stage0_61[236], stage0_61[237]},
      {stage0_63[228], stage0_63[229], stage0_63[230], stage0_63[231], stage0_63[232], stage0_63[233]},
      {stage1_65[38],stage1_64[60],stage1_63[61],stage1_62[74],stage1_61[105]}
   );
   gpc606_5 gpc1227 (
      {stage0_61[238], stage0_61[239], stage0_61[240], stage0_61[241], stage0_61[242], stage0_61[243]},
      {stage0_63[234], stage0_63[235], stage0_63[236], stage0_63[237], stage0_63[238], stage0_63[239]},
      {stage1_65[39],stage1_64[61],stage1_63[62],stage1_62[75],stage1_61[106]}
   );
   gpc606_5 gpc1228 (
      {stage0_61[244], stage0_61[245], stage0_61[246], stage0_61[247], stage0_61[248], stage0_61[249]},
      {stage0_63[240], stage0_63[241], stage0_63[242], stage0_63[243], stage0_63[244], stage0_63[245]},
      {stage1_65[40],stage1_64[62],stage1_63[63],stage1_62[76],stage1_61[107]}
   );
   gpc606_5 gpc1229 (
      {stage0_61[250], stage0_61[251], stage0_61[252], stage0_61[253], stage0_61[254], stage0_61[255]},
      {stage0_63[246], stage0_63[247], stage0_63[248], stage0_63[249], stage0_63[250], stage0_63[251]},
      {stage1_65[41],stage1_64[63],stage1_63[64],stage1_62[77],stage1_61[108]}
   );
   gpc1_1 gpc1230 (
      {stage0_0[212]},
      {stage1_0[47]}
   );
   gpc1_1 gpc1231 (
      {stage0_0[213]},
      {stage1_0[48]}
   );
   gpc1_1 gpc1232 (
      {stage0_0[214]},
      {stage1_0[49]}
   );
   gpc1_1 gpc1233 (
      {stage0_0[215]},
      {stage1_0[50]}
   );
   gpc1_1 gpc1234 (
      {stage0_0[216]},
      {stage1_0[51]}
   );
   gpc1_1 gpc1235 (
      {stage0_0[217]},
      {stage1_0[52]}
   );
   gpc1_1 gpc1236 (
      {stage0_0[218]},
      {stage1_0[53]}
   );
   gpc1_1 gpc1237 (
      {stage0_0[219]},
      {stage1_0[54]}
   );
   gpc1_1 gpc1238 (
      {stage0_0[220]},
      {stage1_0[55]}
   );
   gpc1_1 gpc1239 (
      {stage0_0[221]},
      {stage1_0[56]}
   );
   gpc1_1 gpc1240 (
      {stage0_0[222]},
      {stage1_0[57]}
   );
   gpc1_1 gpc1241 (
      {stage0_0[223]},
      {stage1_0[58]}
   );
   gpc1_1 gpc1242 (
      {stage0_0[224]},
      {stage1_0[59]}
   );
   gpc1_1 gpc1243 (
      {stage0_0[225]},
      {stage1_0[60]}
   );
   gpc1_1 gpc1244 (
      {stage0_0[226]},
      {stage1_0[61]}
   );
   gpc1_1 gpc1245 (
      {stage0_0[227]},
      {stage1_0[62]}
   );
   gpc1_1 gpc1246 (
      {stage0_0[228]},
      {stage1_0[63]}
   );
   gpc1_1 gpc1247 (
      {stage0_0[229]},
      {stage1_0[64]}
   );
   gpc1_1 gpc1248 (
      {stage0_0[230]},
      {stage1_0[65]}
   );
   gpc1_1 gpc1249 (
      {stage0_0[231]},
      {stage1_0[66]}
   );
   gpc1_1 gpc1250 (
      {stage0_0[232]},
      {stage1_0[67]}
   );
   gpc1_1 gpc1251 (
      {stage0_0[233]},
      {stage1_0[68]}
   );
   gpc1_1 gpc1252 (
      {stage0_0[234]},
      {stage1_0[69]}
   );
   gpc1_1 gpc1253 (
      {stage0_0[235]},
      {stage1_0[70]}
   );
   gpc1_1 gpc1254 (
      {stage0_0[236]},
      {stage1_0[71]}
   );
   gpc1_1 gpc1255 (
      {stage0_0[237]},
      {stage1_0[72]}
   );
   gpc1_1 gpc1256 (
      {stage0_0[238]},
      {stage1_0[73]}
   );
   gpc1_1 gpc1257 (
      {stage0_0[239]},
      {stage1_0[74]}
   );
   gpc1_1 gpc1258 (
      {stage0_0[240]},
      {stage1_0[75]}
   );
   gpc1_1 gpc1259 (
      {stage0_0[241]},
      {stage1_0[76]}
   );
   gpc1_1 gpc1260 (
      {stage0_0[242]},
      {stage1_0[77]}
   );
   gpc1_1 gpc1261 (
      {stage0_0[243]},
      {stage1_0[78]}
   );
   gpc1_1 gpc1262 (
      {stage0_0[244]},
      {stage1_0[79]}
   );
   gpc1_1 gpc1263 (
      {stage0_0[245]},
      {stage1_0[80]}
   );
   gpc1_1 gpc1264 (
      {stage0_0[246]},
      {stage1_0[81]}
   );
   gpc1_1 gpc1265 (
      {stage0_0[247]},
      {stage1_0[82]}
   );
   gpc1_1 gpc1266 (
      {stage0_0[248]},
      {stage1_0[83]}
   );
   gpc1_1 gpc1267 (
      {stage0_0[249]},
      {stage1_0[84]}
   );
   gpc1_1 gpc1268 (
      {stage0_0[250]},
      {stage1_0[85]}
   );
   gpc1_1 gpc1269 (
      {stage0_0[251]},
      {stage1_0[86]}
   );
   gpc1_1 gpc1270 (
      {stage0_0[252]},
      {stage1_0[87]}
   );
   gpc1_1 gpc1271 (
      {stage0_0[253]},
      {stage1_0[88]}
   );
   gpc1_1 gpc1272 (
      {stage0_0[254]},
      {stage1_0[89]}
   );
   gpc1_1 gpc1273 (
      {stage0_0[255]},
      {stage1_0[90]}
   );
   gpc1_1 gpc1274 (
      {stage0_1[234]},
      {stage1_1[61]}
   );
   gpc1_1 gpc1275 (
      {stage0_1[235]},
      {stage1_1[62]}
   );
   gpc1_1 gpc1276 (
      {stage0_1[236]},
      {stage1_1[63]}
   );
   gpc1_1 gpc1277 (
      {stage0_1[237]},
      {stage1_1[64]}
   );
   gpc1_1 gpc1278 (
      {stage0_1[238]},
      {stage1_1[65]}
   );
   gpc1_1 gpc1279 (
      {stage0_1[239]},
      {stage1_1[66]}
   );
   gpc1_1 gpc1280 (
      {stage0_1[240]},
      {stage1_1[67]}
   );
   gpc1_1 gpc1281 (
      {stage0_1[241]},
      {stage1_1[68]}
   );
   gpc1_1 gpc1282 (
      {stage0_1[242]},
      {stage1_1[69]}
   );
   gpc1_1 gpc1283 (
      {stage0_1[243]},
      {stage1_1[70]}
   );
   gpc1_1 gpc1284 (
      {stage0_1[244]},
      {stage1_1[71]}
   );
   gpc1_1 gpc1285 (
      {stage0_1[245]},
      {stage1_1[72]}
   );
   gpc1_1 gpc1286 (
      {stage0_1[246]},
      {stage1_1[73]}
   );
   gpc1_1 gpc1287 (
      {stage0_1[247]},
      {stage1_1[74]}
   );
   gpc1_1 gpc1288 (
      {stage0_1[248]},
      {stage1_1[75]}
   );
   gpc1_1 gpc1289 (
      {stage0_1[249]},
      {stage1_1[76]}
   );
   gpc1_1 gpc1290 (
      {stage0_1[250]},
      {stage1_1[77]}
   );
   gpc1_1 gpc1291 (
      {stage0_1[251]},
      {stage1_1[78]}
   );
   gpc1_1 gpc1292 (
      {stage0_1[252]},
      {stage1_1[79]}
   );
   gpc1_1 gpc1293 (
      {stage0_1[253]},
      {stage1_1[80]}
   );
   gpc1_1 gpc1294 (
      {stage0_1[254]},
      {stage1_1[81]}
   );
   gpc1_1 gpc1295 (
      {stage0_1[255]},
      {stage1_1[82]}
   );
   gpc1_1 gpc1296 (
      {stage0_2[199]},
      {stage1_2[74]}
   );
   gpc1_1 gpc1297 (
      {stage0_2[200]},
      {stage1_2[75]}
   );
   gpc1_1 gpc1298 (
      {stage0_2[201]},
      {stage1_2[76]}
   );
   gpc1_1 gpc1299 (
      {stage0_2[202]},
      {stage1_2[77]}
   );
   gpc1_1 gpc1300 (
      {stage0_2[203]},
      {stage1_2[78]}
   );
   gpc1_1 gpc1301 (
      {stage0_2[204]},
      {stage1_2[79]}
   );
   gpc1_1 gpc1302 (
      {stage0_2[205]},
      {stage1_2[80]}
   );
   gpc1_1 gpc1303 (
      {stage0_2[206]},
      {stage1_2[81]}
   );
   gpc1_1 gpc1304 (
      {stage0_2[207]},
      {stage1_2[82]}
   );
   gpc1_1 gpc1305 (
      {stage0_2[208]},
      {stage1_2[83]}
   );
   gpc1_1 gpc1306 (
      {stage0_2[209]},
      {stage1_2[84]}
   );
   gpc1_1 gpc1307 (
      {stage0_2[210]},
      {stage1_2[85]}
   );
   gpc1_1 gpc1308 (
      {stage0_2[211]},
      {stage1_2[86]}
   );
   gpc1_1 gpc1309 (
      {stage0_2[212]},
      {stage1_2[87]}
   );
   gpc1_1 gpc1310 (
      {stage0_2[213]},
      {stage1_2[88]}
   );
   gpc1_1 gpc1311 (
      {stage0_2[214]},
      {stage1_2[89]}
   );
   gpc1_1 gpc1312 (
      {stage0_2[215]},
      {stage1_2[90]}
   );
   gpc1_1 gpc1313 (
      {stage0_2[216]},
      {stage1_2[91]}
   );
   gpc1_1 gpc1314 (
      {stage0_2[217]},
      {stage1_2[92]}
   );
   gpc1_1 gpc1315 (
      {stage0_2[218]},
      {stage1_2[93]}
   );
   gpc1_1 gpc1316 (
      {stage0_2[219]},
      {stage1_2[94]}
   );
   gpc1_1 gpc1317 (
      {stage0_2[220]},
      {stage1_2[95]}
   );
   gpc1_1 gpc1318 (
      {stage0_2[221]},
      {stage1_2[96]}
   );
   gpc1_1 gpc1319 (
      {stage0_2[222]},
      {stage1_2[97]}
   );
   gpc1_1 gpc1320 (
      {stage0_2[223]},
      {stage1_2[98]}
   );
   gpc1_1 gpc1321 (
      {stage0_2[224]},
      {stage1_2[99]}
   );
   gpc1_1 gpc1322 (
      {stage0_2[225]},
      {stage1_2[100]}
   );
   gpc1_1 gpc1323 (
      {stage0_2[226]},
      {stage1_2[101]}
   );
   gpc1_1 gpc1324 (
      {stage0_2[227]},
      {stage1_2[102]}
   );
   gpc1_1 gpc1325 (
      {stage0_2[228]},
      {stage1_2[103]}
   );
   gpc1_1 gpc1326 (
      {stage0_2[229]},
      {stage1_2[104]}
   );
   gpc1_1 gpc1327 (
      {stage0_2[230]},
      {stage1_2[105]}
   );
   gpc1_1 gpc1328 (
      {stage0_2[231]},
      {stage1_2[106]}
   );
   gpc1_1 gpc1329 (
      {stage0_2[232]},
      {stage1_2[107]}
   );
   gpc1_1 gpc1330 (
      {stage0_2[233]},
      {stage1_2[108]}
   );
   gpc1_1 gpc1331 (
      {stage0_2[234]},
      {stage1_2[109]}
   );
   gpc1_1 gpc1332 (
      {stage0_2[235]},
      {stage1_2[110]}
   );
   gpc1_1 gpc1333 (
      {stage0_2[236]},
      {stage1_2[111]}
   );
   gpc1_1 gpc1334 (
      {stage0_2[237]},
      {stage1_2[112]}
   );
   gpc1_1 gpc1335 (
      {stage0_2[238]},
      {stage1_2[113]}
   );
   gpc1_1 gpc1336 (
      {stage0_2[239]},
      {stage1_2[114]}
   );
   gpc1_1 gpc1337 (
      {stage0_2[240]},
      {stage1_2[115]}
   );
   gpc1_1 gpc1338 (
      {stage0_2[241]},
      {stage1_2[116]}
   );
   gpc1_1 gpc1339 (
      {stage0_2[242]},
      {stage1_2[117]}
   );
   gpc1_1 gpc1340 (
      {stage0_2[243]},
      {stage1_2[118]}
   );
   gpc1_1 gpc1341 (
      {stage0_2[244]},
      {stage1_2[119]}
   );
   gpc1_1 gpc1342 (
      {stage0_2[245]},
      {stage1_2[120]}
   );
   gpc1_1 gpc1343 (
      {stage0_2[246]},
      {stage1_2[121]}
   );
   gpc1_1 gpc1344 (
      {stage0_2[247]},
      {stage1_2[122]}
   );
   gpc1_1 gpc1345 (
      {stage0_2[248]},
      {stage1_2[123]}
   );
   gpc1_1 gpc1346 (
      {stage0_2[249]},
      {stage1_2[124]}
   );
   gpc1_1 gpc1347 (
      {stage0_2[250]},
      {stage1_2[125]}
   );
   gpc1_1 gpc1348 (
      {stage0_2[251]},
      {stage1_2[126]}
   );
   gpc1_1 gpc1349 (
      {stage0_2[252]},
      {stage1_2[127]}
   );
   gpc1_1 gpc1350 (
      {stage0_2[253]},
      {stage1_2[128]}
   );
   gpc1_1 gpc1351 (
      {stage0_2[254]},
      {stage1_2[129]}
   );
   gpc1_1 gpc1352 (
      {stage0_2[255]},
      {stage1_2[130]}
   );
   gpc1_1 gpc1353 (
      {stage0_3[245]},
      {stage1_3[96]}
   );
   gpc1_1 gpc1354 (
      {stage0_3[246]},
      {stage1_3[97]}
   );
   gpc1_1 gpc1355 (
      {stage0_3[247]},
      {stage1_3[98]}
   );
   gpc1_1 gpc1356 (
      {stage0_3[248]},
      {stage1_3[99]}
   );
   gpc1_1 gpc1357 (
      {stage0_3[249]},
      {stage1_3[100]}
   );
   gpc1_1 gpc1358 (
      {stage0_3[250]},
      {stage1_3[101]}
   );
   gpc1_1 gpc1359 (
      {stage0_3[251]},
      {stage1_3[102]}
   );
   gpc1_1 gpc1360 (
      {stage0_3[252]},
      {stage1_3[103]}
   );
   gpc1_1 gpc1361 (
      {stage0_3[253]},
      {stage1_3[104]}
   );
   gpc1_1 gpc1362 (
      {stage0_3[254]},
      {stage1_3[105]}
   );
   gpc1_1 gpc1363 (
      {stage0_3[255]},
      {stage1_3[106]}
   );
   gpc1_1 gpc1364 (
      {stage0_6[236]},
      {stage1_6[96]}
   );
   gpc1_1 gpc1365 (
      {stage0_6[237]},
      {stage1_6[97]}
   );
   gpc1_1 gpc1366 (
      {stage0_6[238]},
      {stage1_6[98]}
   );
   gpc1_1 gpc1367 (
      {stage0_6[239]},
      {stage1_6[99]}
   );
   gpc1_1 gpc1368 (
      {stage0_6[240]},
      {stage1_6[100]}
   );
   gpc1_1 gpc1369 (
      {stage0_6[241]},
      {stage1_6[101]}
   );
   gpc1_1 gpc1370 (
      {stage0_6[242]},
      {stage1_6[102]}
   );
   gpc1_1 gpc1371 (
      {stage0_6[243]},
      {stage1_6[103]}
   );
   gpc1_1 gpc1372 (
      {stage0_6[244]},
      {stage1_6[104]}
   );
   gpc1_1 gpc1373 (
      {stage0_6[245]},
      {stage1_6[105]}
   );
   gpc1_1 gpc1374 (
      {stage0_6[246]},
      {stage1_6[106]}
   );
   gpc1_1 gpc1375 (
      {stage0_6[247]},
      {stage1_6[107]}
   );
   gpc1_1 gpc1376 (
      {stage0_6[248]},
      {stage1_6[108]}
   );
   gpc1_1 gpc1377 (
      {stage0_6[249]},
      {stage1_6[109]}
   );
   gpc1_1 gpc1378 (
      {stage0_6[250]},
      {stage1_6[110]}
   );
   gpc1_1 gpc1379 (
      {stage0_6[251]},
      {stage1_6[111]}
   );
   gpc1_1 gpc1380 (
      {stage0_6[252]},
      {stage1_6[112]}
   );
   gpc1_1 gpc1381 (
      {stage0_6[253]},
      {stage1_6[113]}
   );
   gpc1_1 gpc1382 (
      {stage0_6[254]},
      {stage1_6[114]}
   );
   gpc1_1 gpc1383 (
      {stage0_6[255]},
      {stage1_6[115]}
   );
   gpc1_1 gpc1384 (
      {stage0_7[251]},
      {stage1_7[105]}
   );
   gpc1_1 gpc1385 (
      {stage0_7[252]},
      {stage1_7[106]}
   );
   gpc1_1 gpc1386 (
      {stage0_7[253]},
      {stage1_7[107]}
   );
   gpc1_1 gpc1387 (
      {stage0_7[254]},
      {stage1_7[108]}
   );
   gpc1_1 gpc1388 (
      {stage0_7[255]},
      {stage1_7[109]}
   );
   gpc1_1 gpc1389 (
      {stage0_8[233]},
      {stage1_8[109]}
   );
   gpc1_1 gpc1390 (
      {stage0_8[234]},
      {stage1_8[110]}
   );
   gpc1_1 gpc1391 (
      {stage0_8[235]},
      {stage1_8[111]}
   );
   gpc1_1 gpc1392 (
      {stage0_8[236]},
      {stage1_8[112]}
   );
   gpc1_1 gpc1393 (
      {stage0_8[237]},
      {stage1_8[113]}
   );
   gpc1_1 gpc1394 (
      {stage0_8[238]},
      {stage1_8[114]}
   );
   gpc1_1 gpc1395 (
      {stage0_8[239]},
      {stage1_8[115]}
   );
   gpc1_1 gpc1396 (
      {stage0_8[240]},
      {stage1_8[116]}
   );
   gpc1_1 gpc1397 (
      {stage0_8[241]},
      {stage1_8[117]}
   );
   gpc1_1 gpc1398 (
      {stage0_8[242]},
      {stage1_8[118]}
   );
   gpc1_1 gpc1399 (
      {stage0_8[243]},
      {stage1_8[119]}
   );
   gpc1_1 gpc1400 (
      {stage0_8[244]},
      {stage1_8[120]}
   );
   gpc1_1 gpc1401 (
      {stage0_8[245]},
      {stage1_8[121]}
   );
   gpc1_1 gpc1402 (
      {stage0_8[246]},
      {stage1_8[122]}
   );
   gpc1_1 gpc1403 (
      {stage0_8[247]},
      {stage1_8[123]}
   );
   gpc1_1 gpc1404 (
      {stage0_8[248]},
      {stage1_8[124]}
   );
   gpc1_1 gpc1405 (
      {stage0_8[249]},
      {stage1_8[125]}
   );
   gpc1_1 gpc1406 (
      {stage0_8[250]},
      {stage1_8[126]}
   );
   gpc1_1 gpc1407 (
      {stage0_8[251]},
      {stage1_8[127]}
   );
   gpc1_1 gpc1408 (
      {stage0_8[252]},
      {stage1_8[128]}
   );
   gpc1_1 gpc1409 (
      {stage0_8[253]},
      {stage1_8[129]}
   );
   gpc1_1 gpc1410 (
      {stage0_8[254]},
      {stage1_8[130]}
   );
   gpc1_1 gpc1411 (
      {stage0_8[255]},
      {stage1_8[131]}
   );
   gpc1_1 gpc1412 (
      {stage0_9[235]},
      {stage1_9[99]}
   );
   gpc1_1 gpc1413 (
      {stage0_9[236]},
      {stage1_9[100]}
   );
   gpc1_1 gpc1414 (
      {stage0_9[237]},
      {stage1_9[101]}
   );
   gpc1_1 gpc1415 (
      {stage0_9[238]},
      {stage1_9[102]}
   );
   gpc1_1 gpc1416 (
      {stage0_9[239]},
      {stage1_9[103]}
   );
   gpc1_1 gpc1417 (
      {stage0_9[240]},
      {stage1_9[104]}
   );
   gpc1_1 gpc1418 (
      {stage0_9[241]},
      {stage1_9[105]}
   );
   gpc1_1 gpc1419 (
      {stage0_9[242]},
      {stage1_9[106]}
   );
   gpc1_1 gpc1420 (
      {stage0_9[243]},
      {stage1_9[107]}
   );
   gpc1_1 gpc1421 (
      {stage0_9[244]},
      {stage1_9[108]}
   );
   gpc1_1 gpc1422 (
      {stage0_9[245]},
      {stage1_9[109]}
   );
   gpc1_1 gpc1423 (
      {stage0_9[246]},
      {stage1_9[110]}
   );
   gpc1_1 gpc1424 (
      {stage0_9[247]},
      {stage1_9[111]}
   );
   gpc1_1 gpc1425 (
      {stage0_9[248]},
      {stage1_9[112]}
   );
   gpc1_1 gpc1426 (
      {stage0_9[249]},
      {stage1_9[113]}
   );
   gpc1_1 gpc1427 (
      {stage0_9[250]},
      {stage1_9[114]}
   );
   gpc1_1 gpc1428 (
      {stage0_9[251]},
      {stage1_9[115]}
   );
   gpc1_1 gpc1429 (
      {stage0_9[252]},
      {stage1_9[116]}
   );
   gpc1_1 gpc1430 (
      {stage0_9[253]},
      {stage1_9[117]}
   );
   gpc1_1 gpc1431 (
      {stage0_9[254]},
      {stage1_9[118]}
   );
   gpc1_1 gpc1432 (
      {stage0_9[255]},
      {stage1_9[119]}
   );
   gpc1_1 gpc1433 (
      {stage0_10[181]},
      {stage1_10[81]}
   );
   gpc1_1 gpc1434 (
      {stage0_10[182]},
      {stage1_10[82]}
   );
   gpc1_1 gpc1435 (
      {stage0_10[183]},
      {stage1_10[83]}
   );
   gpc1_1 gpc1436 (
      {stage0_10[184]},
      {stage1_10[84]}
   );
   gpc1_1 gpc1437 (
      {stage0_10[185]},
      {stage1_10[85]}
   );
   gpc1_1 gpc1438 (
      {stage0_10[186]},
      {stage1_10[86]}
   );
   gpc1_1 gpc1439 (
      {stage0_10[187]},
      {stage1_10[87]}
   );
   gpc1_1 gpc1440 (
      {stage0_10[188]},
      {stage1_10[88]}
   );
   gpc1_1 gpc1441 (
      {stage0_10[189]},
      {stage1_10[89]}
   );
   gpc1_1 gpc1442 (
      {stage0_10[190]},
      {stage1_10[90]}
   );
   gpc1_1 gpc1443 (
      {stage0_10[191]},
      {stage1_10[91]}
   );
   gpc1_1 gpc1444 (
      {stage0_10[192]},
      {stage1_10[92]}
   );
   gpc1_1 gpc1445 (
      {stage0_10[193]},
      {stage1_10[93]}
   );
   gpc1_1 gpc1446 (
      {stage0_10[194]},
      {stage1_10[94]}
   );
   gpc1_1 gpc1447 (
      {stage0_10[195]},
      {stage1_10[95]}
   );
   gpc1_1 gpc1448 (
      {stage0_10[196]},
      {stage1_10[96]}
   );
   gpc1_1 gpc1449 (
      {stage0_10[197]},
      {stage1_10[97]}
   );
   gpc1_1 gpc1450 (
      {stage0_10[198]},
      {stage1_10[98]}
   );
   gpc1_1 gpc1451 (
      {stage0_10[199]},
      {stage1_10[99]}
   );
   gpc1_1 gpc1452 (
      {stage0_10[200]},
      {stage1_10[100]}
   );
   gpc1_1 gpc1453 (
      {stage0_10[201]},
      {stage1_10[101]}
   );
   gpc1_1 gpc1454 (
      {stage0_10[202]},
      {stage1_10[102]}
   );
   gpc1_1 gpc1455 (
      {stage0_10[203]},
      {stage1_10[103]}
   );
   gpc1_1 gpc1456 (
      {stage0_10[204]},
      {stage1_10[104]}
   );
   gpc1_1 gpc1457 (
      {stage0_10[205]},
      {stage1_10[105]}
   );
   gpc1_1 gpc1458 (
      {stage0_10[206]},
      {stage1_10[106]}
   );
   gpc1_1 gpc1459 (
      {stage0_10[207]},
      {stage1_10[107]}
   );
   gpc1_1 gpc1460 (
      {stage0_10[208]},
      {stage1_10[108]}
   );
   gpc1_1 gpc1461 (
      {stage0_10[209]},
      {stage1_10[109]}
   );
   gpc1_1 gpc1462 (
      {stage0_10[210]},
      {stage1_10[110]}
   );
   gpc1_1 gpc1463 (
      {stage0_10[211]},
      {stage1_10[111]}
   );
   gpc1_1 gpc1464 (
      {stage0_10[212]},
      {stage1_10[112]}
   );
   gpc1_1 gpc1465 (
      {stage0_10[213]},
      {stage1_10[113]}
   );
   gpc1_1 gpc1466 (
      {stage0_10[214]},
      {stage1_10[114]}
   );
   gpc1_1 gpc1467 (
      {stage0_10[215]},
      {stage1_10[115]}
   );
   gpc1_1 gpc1468 (
      {stage0_10[216]},
      {stage1_10[116]}
   );
   gpc1_1 gpc1469 (
      {stage0_10[217]},
      {stage1_10[117]}
   );
   gpc1_1 gpc1470 (
      {stage0_10[218]},
      {stage1_10[118]}
   );
   gpc1_1 gpc1471 (
      {stage0_10[219]},
      {stage1_10[119]}
   );
   gpc1_1 gpc1472 (
      {stage0_10[220]},
      {stage1_10[120]}
   );
   gpc1_1 gpc1473 (
      {stage0_10[221]},
      {stage1_10[121]}
   );
   gpc1_1 gpc1474 (
      {stage0_10[222]},
      {stage1_10[122]}
   );
   gpc1_1 gpc1475 (
      {stage0_10[223]},
      {stage1_10[123]}
   );
   gpc1_1 gpc1476 (
      {stage0_10[224]},
      {stage1_10[124]}
   );
   gpc1_1 gpc1477 (
      {stage0_10[225]},
      {stage1_10[125]}
   );
   gpc1_1 gpc1478 (
      {stage0_10[226]},
      {stage1_10[126]}
   );
   gpc1_1 gpc1479 (
      {stage0_10[227]},
      {stage1_10[127]}
   );
   gpc1_1 gpc1480 (
      {stage0_10[228]},
      {stage1_10[128]}
   );
   gpc1_1 gpc1481 (
      {stage0_10[229]},
      {stage1_10[129]}
   );
   gpc1_1 gpc1482 (
      {stage0_10[230]},
      {stage1_10[130]}
   );
   gpc1_1 gpc1483 (
      {stage0_10[231]},
      {stage1_10[131]}
   );
   gpc1_1 gpc1484 (
      {stage0_10[232]},
      {stage1_10[132]}
   );
   gpc1_1 gpc1485 (
      {stage0_10[233]},
      {stage1_10[133]}
   );
   gpc1_1 gpc1486 (
      {stage0_10[234]},
      {stage1_10[134]}
   );
   gpc1_1 gpc1487 (
      {stage0_10[235]},
      {stage1_10[135]}
   );
   gpc1_1 gpc1488 (
      {stage0_10[236]},
      {stage1_10[136]}
   );
   gpc1_1 gpc1489 (
      {stage0_10[237]},
      {stage1_10[137]}
   );
   gpc1_1 gpc1490 (
      {stage0_10[238]},
      {stage1_10[138]}
   );
   gpc1_1 gpc1491 (
      {stage0_10[239]},
      {stage1_10[139]}
   );
   gpc1_1 gpc1492 (
      {stage0_10[240]},
      {stage1_10[140]}
   );
   gpc1_1 gpc1493 (
      {stage0_10[241]},
      {stage1_10[141]}
   );
   gpc1_1 gpc1494 (
      {stage0_10[242]},
      {stage1_10[142]}
   );
   gpc1_1 gpc1495 (
      {stage0_10[243]},
      {stage1_10[143]}
   );
   gpc1_1 gpc1496 (
      {stage0_10[244]},
      {stage1_10[144]}
   );
   gpc1_1 gpc1497 (
      {stage0_10[245]},
      {stage1_10[145]}
   );
   gpc1_1 gpc1498 (
      {stage0_10[246]},
      {stage1_10[146]}
   );
   gpc1_1 gpc1499 (
      {stage0_10[247]},
      {stage1_10[147]}
   );
   gpc1_1 gpc1500 (
      {stage0_10[248]},
      {stage1_10[148]}
   );
   gpc1_1 gpc1501 (
      {stage0_10[249]},
      {stage1_10[149]}
   );
   gpc1_1 gpc1502 (
      {stage0_10[250]},
      {stage1_10[150]}
   );
   gpc1_1 gpc1503 (
      {stage0_10[251]},
      {stage1_10[151]}
   );
   gpc1_1 gpc1504 (
      {stage0_10[252]},
      {stage1_10[152]}
   );
   gpc1_1 gpc1505 (
      {stage0_10[253]},
      {stage1_10[153]}
   );
   gpc1_1 gpc1506 (
      {stage0_10[254]},
      {stage1_10[154]}
   );
   gpc1_1 gpc1507 (
      {stage0_10[255]},
      {stage1_10[155]}
   );
   gpc1_1 gpc1508 (
      {stage0_11[183]},
      {stage1_11[81]}
   );
   gpc1_1 gpc1509 (
      {stage0_11[184]},
      {stage1_11[82]}
   );
   gpc1_1 gpc1510 (
      {stage0_11[185]},
      {stage1_11[83]}
   );
   gpc1_1 gpc1511 (
      {stage0_11[186]},
      {stage1_11[84]}
   );
   gpc1_1 gpc1512 (
      {stage0_11[187]},
      {stage1_11[85]}
   );
   gpc1_1 gpc1513 (
      {stage0_11[188]},
      {stage1_11[86]}
   );
   gpc1_1 gpc1514 (
      {stage0_11[189]},
      {stage1_11[87]}
   );
   gpc1_1 gpc1515 (
      {stage0_11[190]},
      {stage1_11[88]}
   );
   gpc1_1 gpc1516 (
      {stage0_11[191]},
      {stage1_11[89]}
   );
   gpc1_1 gpc1517 (
      {stage0_11[192]},
      {stage1_11[90]}
   );
   gpc1_1 gpc1518 (
      {stage0_11[193]},
      {stage1_11[91]}
   );
   gpc1_1 gpc1519 (
      {stage0_11[194]},
      {stage1_11[92]}
   );
   gpc1_1 gpc1520 (
      {stage0_11[195]},
      {stage1_11[93]}
   );
   gpc1_1 gpc1521 (
      {stage0_11[196]},
      {stage1_11[94]}
   );
   gpc1_1 gpc1522 (
      {stage0_11[197]},
      {stage1_11[95]}
   );
   gpc1_1 gpc1523 (
      {stage0_11[198]},
      {stage1_11[96]}
   );
   gpc1_1 gpc1524 (
      {stage0_11[199]},
      {stage1_11[97]}
   );
   gpc1_1 gpc1525 (
      {stage0_11[200]},
      {stage1_11[98]}
   );
   gpc1_1 gpc1526 (
      {stage0_11[201]},
      {stage1_11[99]}
   );
   gpc1_1 gpc1527 (
      {stage0_11[202]},
      {stage1_11[100]}
   );
   gpc1_1 gpc1528 (
      {stage0_11[203]},
      {stage1_11[101]}
   );
   gpc1_1 gpc1529 (
      {stage0_11[204]},
      {stage1_11[102]}
   );
   gpc1_1 gpc1530 (
      {stage0_11[205]},
      {stage1_11[103]}
   );
   gpc1_1 gpc1531 (
      {stage0_11[206]},
      {stage1_11[104]}
   );
   gpc1_1 gpc1532 (
      {stage0_11[207]},
      {stage1_11[105]}
   );
   gpc1_1 gpc1533 (
      {stage0_11[208]},
      {stage1_11[106]}
   );
   gpc1_1 gpc1534 (
      {stage0_11[209]},
      {stage1_11[107]}
   );
   gpc1_1 gpc1535 (
      {stage0_11[210]},
      {stage1_11[108]}
   );
   gpc1_1 gpc1536 (
      {stage0_11[211]},
      {stage1_11[109]}
   );
   gpc1_1 gpc1537 (
      {stage0_11[212]},
      {stage1_11[110]}
   );
   gpc1_1 gpc1538 (
      {stage0_11[213]},
      {stage1_11[111]}
   );
   gpc1_1 gpc1539 (
      {stage0_11[214]},
      {stage1_11[112]}
   );
   gpc1_1 gpc1540 (
      {stage0_11[215]},
      {stage1_11[113]}
   );
   gpc1_1 gpc1541 (
      {stage0_11[216]},
      {stage1_11[114]}
   );
   gpc1_1 gpc1542 (
      {stage0_11[217]},
      {stage1_11[115]}
   );
   gpc1_1 gpc1543 (
      {stage0_11[218]},
      {stage1_11[116]}
   );
   gpc1_1 gpc1544 (
      {stage0_11[219]},
      {stage1_11[117]}
   );
   gpc1_1 gpc1545 (
      {stage0_11[220]},
      {stage1_11[118]}
   );
   gpc1_1 gpc1546 (
      {stage0_11[221]},
      {stage1_11[119]}
   );
   gpc1_1 gpc1547 (
      {stage0_11[222]},
      {stage1_11[120]}
   );
   gpc1_1 gpc1548 (
      {stage0_11[223]},
      {stage1_11[121]}
   );
   gpc1_1 gpc1549 (
      {stage0_11[224]},
      {stage1_11[122]}
   );
   gpc1_1 gpc1550 (
      {stage0_11[225]},
      {stage1_11[123]}
   );
   gpc1_1 gpc1551 (
      {stage0_11[226]},
      {stage1_11[124]}
   );
   gpc1_1 gpc1552 (
      {stage0_11[227]},
      {stage1_11[125]}
   );
   gpc1_1 gpc1553 (
      {stage0_11[228]},
      {stage1_11[126]}
   );
   gpc1_1 gpc1554 (
      {stage0_11[229]},
      {stage1_11[127]}
   );
   gpc1_1 gpc1555 (
      {stage0_11[230]},
      {stage1_11[128]}
   );
   gpc1_1 gpc1556 (
      {stage0_11[231]},
      {stage1_11[129]}
   );
   gpc1_1 gpc1557 (
      {stage0_11[232]},
      {stage1_11[130]}
   );
   gpc1_1 gpc1558 (
      {stage0_11[233]},
      {stage1_11[131]}
   );
   gpc1_1 gpc1559 (
      {stage0_11[234]},
      {stage1_11[132]}
   );
   gpc1_1 gpc1560 (
      {stage0_11[235]},
      {stage1_11[133]}
   );
   gpc1_1 gpc1561 (
      {stage0_11[236]},
      {stage1_11[134]}
   );
   gpc1_1 gpc1562 (
      {stage0_11[237]},
      {stage1_11[135]}
   );
   gpc1_1 gpc1563 (
      {stage0_11[238]},
      {stage1_11[136]}
   );
   gpc1_1 gpc1564 (
      {stage0_11[239]},
      {stage1_11[137]}
   );
   gpc1_1 gpc1565 (
      {stage0_11[240]},
      {stage1_11[138]}
   );
   gpc1_1 gpc1566 (
      {stage0_11[241]},
      {stage1_11[139]}
   );
   gpc1_1 gpc1567 (
      {stage0_11[242]},
      {stage1_11[140]}
   );
   gpc1_1 gpc1568 (
      {stage0_11[243]},
      {stage1_11[141]}
   );
   gpc1_1 gpc1569 (
      {stage0_11[244]},
      {stage1_11[142]}
   );
   gpc1_1 gpc1570 (
      {stage0_11[245]},
      {stage1_11[143]}
   );
   gpc1_1 gpc1571 (
      {stage0_11[246]},
      {stage1_11[144]}
   );
   gpc1_1 gpc1572 (
      {stage0_11[247]},
      {stage1_11[145]}
   );
   gpc1_1 gpc1573 (
      {stage0_11[248]},
      {stage1_11[146]}
   );
   gpc1_1 gpc1574 (
      {stage0_11[249]},
      {stage1_11[147]}
   );
   gpc1_1 gpc1575 (
      {stage0_11[250]},
      {stage1_11[148]}
   );
   gpc1_1 gpc1576 (
      {stage0_11[251]},
      {stage1_11[149]}
   );
   gpc1_1 gpc1577 (
      {stage0_11[252]},
      {stage1_11[150]}
   );
   gpc1_1 gpc1578 (
      {stage0_11[253]},
      {stage1_11[151]}
   );
   gpc1_1 gpc1579 (
      {stage0_11[254]},
      {stage1_11[152]}
   );
   gpc1_1 gpc1580 (
      {stage0_11[255]},
      {stage1_11[153]}
   );
   gpc1_1 gpc1581 (
      {stage0_12[220]},
      {stage1_12[97]}
   );
   gpc1_1 gpc1582 (
      {stage0_12[221]},
      {stage1_12[98]}
   );
   gpc1_1 gpc1583 (
      {stage0_12[222]},
      {stage1_12[99]}
   );
   gpc1_1 gpc1584 (
      {stage0_12[223]},
      {stage1_12[100]}
   );
   gpc1_1 gpc1585 (
      {stage0_12[224]},
      {stage1_12[101]}
   );
   gpc1_1 gpc1586 (
      {stage0_12[225]},
      {stage1_12[102]}
   );
   gpc1_1 gpc1587 (
      {stage0_12[226]},
      {stage1_12[103]}
   );
   gpc1_1 gpc1588 (
      {stage0_12[227]},
      {stage1_12[104]}
   );
   gpc1_1 gpc1589 (
      {stage0_12[228]},
      {stage1_12[105]}
   );
   gpc1_1 gpc1590 (
      {stage0_12[229]},
      {stage1_12[106]}
   );
   gpc1_1 gpc1591 (
      {stage0_12[230]},
      {stage1_12[107]}
   );
   gpc1_1 gpc1592 (
      {stage0_12[231]},
      {stage1_12[108]}
   );
   gpc1_1 gpc1593 (
      {stage0_12[232]},
      {stage1_12[109]}
   );
   gpc1_1 gpc1594 (
      {stage0_12[233]},
      {stage1_12[110]}
   );
   gpc1_1 gpc1595 (
      {stage0_12[234]},
      {stage1_12[111]}
   );
   gpc1_1 gpc1596 (
      {stage0_12[235]},
      {stage1_12[112]}
   );
   gpc1_1 gpc1597 (
      {stage0_12[236]},
      {stage1_12[113]}
   );
   gpc1_1 gpc1598 (
      {stage0_12[237]},
      {stage1_12[114]}
   );
   gpc1_1 gpc1599 (
      {stage0_12[238]},
      {stage1_12[115]}
   );
   gpc1_1 gpc1600 (
      {stage0_12[239]},
      {stage1_12[116]}
   );
   gpc1_1 gpc1601 (
      {stage0_12[240]},
      {stage1_12[117]}
   );
   gpc1_1 gpc1602 (
      {stage0_12[241]},
      {stage1_12[118]}
   );
   gpc1_1 gpc1603 (
      {stage0_12[242]},
      {stage1_12[119]}
   );
   gpc1_1 gpc1604 (
      {stage0_12[243]},
      {stage1_12[120]}
   );
   gpc1_1 gpc1605 (
      {stage0_12[244]},
      {stage1_12[121]}
   );
   gpc1_1 gpc1606 (
      {stage0_12[245]},
      {stage1_12[122]}
   );
   gpc1_1 gpc1607 (
      {stage0_12[246]},
      {stage1_12[123]}
   );
   gpc1_1 gpc1608 (
      {stage0_12[247]},
      {stage1_12[124]}
   );
   gpc1_1 gpc1609 (
      {stage0_12[248]},
      {stage1_12[125]}
   );
   gpc1_1 gpc1610 (
      {stage0_12[249]},
      {stage1_12[126]}
   );
   gpc1_1 gpc1611 (
      {stage0_12[250]},
      {stage1_12[127]}
   );
   gpc1_1 gpc1612 (
      {stage0_12[251]},
      {stage1_12[128]}
   );
   gpc1_1 gpc1613 (
      {stage0_12[252]},
      {stage1_12[129]}
   );
   gpc1_1 gpc1614 (
      {stage0_12[253]},
      {stage1_12[130]}
   );
   gpc1_1 gpc1615 (
      {stage0_12[254]},
      {stage1_12[131]}
   );
   gpc1_1 gpc1616 (
      {stage0_12[255]},
      {stage1_12[132]}
   );
   gpc1_1 gpc1617 (
      {stage0_13[254]},
      {stage1_13[95]}
   );
   gpc1_1 gpc1618 (
      {stage0_13[255]},
      {stage1_13[96]}
   );
   gpc1_1 gpc1619 (
      {stage0_15[220]},
      {stage1_15[96]}
   );
   gpc1_1 gpc1620 (
      {stage0_15[221]},
      {stage1_15[97]}
   );
   gpc1_1 gpc1621 (
      {stage0_15[222]},
      {stage1_15[98]}
   );
   gpc1_1 gpc1622 (
      {stage0_15[223]},
      {stage1_15[99]}
   );
   gpc1_1 gpc1623 (
      {stage0_15[224]},
      {stage1_15[100]}
   );
   gpc1_1 gpc1624 (
      {stage0_15[225]},
      {stage1_15[101]}
   );
   gpc1_1 gpc1625 (
      {stage0_15[226]},
      {stage1_15[102]}
   );
   gpc1_1 gpc1626 (
      {stage0_15[227]},
      {stage1_15[103]}
   );
   gpc1_1 gpc1627 (
      {stage0_15[228]},
      {stage1_15[104]}
   );
   gpc1_1 gpc1628 (
      {stage0_15[229]},
      {stage1_15[105]}
   );
   gpc1_1 gpc1629 (
      {stage0_15[230]},
      {stage1_15[106]}
   );
   gpc1_1 gpc1630 (
      {stage0_15[231]},
      {stage1_15[107]}
   );
   gpc1_1 gpc1631 (
      {stage0_15[232]},
      {stage1_15[108]}
   );
   gpc1_1 gpc1632 (
      {stage0_15[233]},
      {stage1_15[109]}
   );
   gpc1_1 gpc1633 (
      {stage0_15[234]},
      {stage1_15[110]}
   );
   gpc1_1 gpc1634 (
      {stage0_15[235]},
      {stage1_15[111]}
   );
   gpc1_1 gpc1635 (
      {stage0_15[236]},
      {stage1_15[112]}
   );
   gpc1_1 gpc1636 (
      {stage0_15[237]},
      {stage1_15[113]}
   );
   gpc1_1 gpc1637 (
      {stage0_15[238]},
      {stage1_15[114]}
   );
   gpc1_1 gpc1638 (
      {stage0_15[239]},
      {stage1_15[115]}
   );
   gpc1_1 gpc1639 (
      {stage0_15[240]},
      {stage1_15[116]}
   );
   gpc1_1 gpc1640 (
      {stage0_15[241]},
      {stage1_15[117]}
   );
   gpc1_1 gpc1641 (
      {stage0_15[242]},
      {stage1_15[118]}
   );
   gpc1_1 gpc1642 (
      {stage0_15[243]},
      {stage1_15[119]}
   );
   gpc1_1 gpc1643 (
      {stage0_15[244]},
      {stage1_15[120]}
   );
   gpc1_1 gpc1644 (
      {stage0_15[245]},
      {stage1_15[121]}
   );
   gpc1_1 gpc1645 (
      {stage0_15[246]},
      {stage1_15[122]}
   );
   gpc1_1 gpc1646 (
      {stage0_15[247]},
      {stage1_15[123]}
   );
   gpc1_1 gpc1647 (
      {stage0_15[248]},
      {stage1_15[124]}
   );
   gpc1_1 gpc1648 (
      {stage0_15[249]},
      {stage1_15[125]}
   );
   gpc1_1 gpc1649 (
      {stage0_15[250]},
      {stage1_15[126]}
   );
   gpc1_1 gpc1650 (
      {stage0_15[251]},
      {stage1_15[127]}
   );
   gpc1_1 gpc1651 (
      {stage0_15[252]},
      {stage1_15[128]}
   );
   gpc1_1 gpc1652 (
      {stage0_15[253]},
      {stage1_15[129]}
   );
   gpc1_1 gpc1653 (
      {stage0_15[254]},
      {stage1_15[130]}
   );
   gpc1_1 gpc1654 (
      {stage0_15[255]},
      {stage1_15[131]}
   );
   gpc1_1 gpc1655 (
      {stage0_16[255]},
      {stage1_16[119]}
   );
   gpc1_1 gpc1656 (
      {stage0_17[251]},
      {stage1_17[106]}
   );
   gpc1_1 gpc1657 (
      {stage0_17[252]},
      {stage1_17[107]}
   );
   gpc1_1 gpc1658 (
      {stage0_17[253]},
      {stage1_17[108]}
   );
   gpc1_1 gpc1659 (
      {stage0_17[254]},
      {stage1_17[109]}
   );
   gpc1_1 gpc1660 (
      {stage0_17[255]},
      {stage1_17[110]}
   );
   gpc1_1 gpc1661 (
      {stage0_18[242]},
      {stage1_18[86]}
   );
   gpc1_1 gpc1662 (
      {stage0_18[243]},
      {stage1_18[87]}
   );
   gpc1_1 gpc1663 (
      {stage0_18[244]},
      {stage1_18[88]}
   );
   gpc1_1 gpc1664 (
      {stage0_18[245]},
      {stage1_18[89]}
   );
   gpc1_1 gpc1665 (
      {stage0_18[246]},
      {stage1_18[90]}
   );
   gpc1_1 gpc1666 (
      {stage0_18[247]},
      {stage1_18[91]}
   );
   gpc1_1 gpc1667 (
      {stage0_18[248]},
      {stage1_18[92]}
   );
   gpc1_1 gpc1668 (
      {stage0_18[249]},
      {stage1_18[93]}
   );
   gpc1_1 gpc1669 (
      {stage0_18[250]},
      {stage1_18[94]}
   );
   gpc1_1 gpc1670 (
      {stage0_18[251]},
      {stage1_18[95]}
   );
   gpc1_1 gpc1671 (
      {stage0_18[252]},
      {stage1_18[96]}
   );
   gpc1_1 gpc1672 (
      {stage0_18[253]},
      {stage1_18[97]}
   );
   gpc1_1 gpc1673 (
      {stage0_18[254]},
      {stage1_18[98]}
   );
   gpc1_1 gpc1674 (
      {stage0_18[255]},
      {stage1_18[99]}
   );
   gpc1_1 gpc1675 (
      {stage0_19[224]},
      {stage1_19[94]}
   );
   gpc1_1 gpc1676 (
      {stage0_19[225]},
      {stage1_19[95]}
   );
   gpc1_1 gpc1677 (
      {stage0_19[226]},
      {stage1_19[96]}
   );
   gpc1_1 gpc1678 (
      {stage0_19[227]},
      {stage1_19[97]}
   );
   gpc1_1 gpc1679 (
      {stage0_19[228]},
      {stage1_19[98]}
   );
   gpc1_1 gpc1680 (
      {stage0_19[229]},
      {stage1_19[99]}
   );
   gpc1_1 gpc1681 (
      {stage0_19[230]},
      {stage1_19[100]}
   );
   gpc1_1 gpc1682 (
      {stage0_19[231]},
      {stage1_19[101]}
   );
   gpc1_1 gpc1683 (
      {stage0_19[232]},
      {stage1_19[102]}
   );
   gpc1_1 gpc1684 (
      {stage0_19[233]},
      {stage1_19[103]}
   );
   gpc1_1 gpc1685 (
      {stage0_19[234]},
      {stage1_19[104]}
   );
   gpc1_1 gpc1686 (
      {stage0_19[235]},
      {stage1_19[105]}
   );
   gpc1_1 gpc1687 (
      {stage0_19[236]},
      {stage1_19[106]}
   );
   gpc1_1 gpc1688 (
      {stage0_19[237]},
      {stage1_19[107]}
   );
   gpc1_1 gpc1689 (
      {stage0_19[238]},
      {stage1_19[108]}
   );
   gpc1_1 gpc1690 (
      {stage0_19[239]},
      {stage1_19[109]}
   );
   gpc1_1 gpc1691 (
      {stage0_19[240]},
      {stage1_19[110]}
   );
   gpc1_1 gpc1692 (
      {stage0_19[241]},
      {stage1_19[111]}
   );
   gpc1_1 gpc1693 (
      {stage0_19[242]},
      {stage1_19[112]}
   );
   gpc1_1 gpc1694 (
      {stage0_19[243]},
      {stage1_19[113]}
   );
   gpc1_1 gpc1695 (
      {stage0_19[244]},
      {stage1_19[114]}
   );
   gpc1_1 gpc1696 (
      {stage0_19[245]},
      {stage1_19[115]}
   );
   gpc1_1 gpc1697 (
      {stage0_19[246]},
      {stage1_19[116]}
   );
   gpc1_1 gpc1698 (
      {stage0_19[247]},
      {stage1_19[117]}
   );
   gpc1_1 gpc1699 (
      {stage0_19[248]},
      {stage1_19[118]}
   );
   gpc1_1 gpc1700 (
      {stage0_19[249]},
      {stage1_19[119]}
   );
   gpc1_1 gpc1701 (
      {stage0_19[250]},
      {stage1_19[120]}
   );
   gpc1_1 gpc1702 (
      {stage0_19[251]},
      {stage1_19[121]}
   );
   gpc1_1 gpc1703 (
      {stage0_19[252]},
      {stage1_19[122]}
   );
   gpc1_1 gpc1704 (
      {stage0_19[253]},
      {stage1_19[123]}
   );
   gpc1_1 gpc1705 (
      {stage0_19[254]},
      {stage1_19[124]}
   );
   gpc1_1 gpc1706 (
      {stage0_19[255]},
      {stage1_19[125]}
   );
   gpc1_1 gpc1707 (
      {stage0_20[245]},
      {stage1_20[119]}
   );
   gpc1_1 gpc1708 (
      {stage0_20[246]},
      {stage1_20[120]}
   );
   gpc1_1 gpc1709 (
      {stage0_20[247]},
      {stage1_20[121]}
   );
   gpc1_1 gpc1710 (
      {stage0_20[248]},
      {stage1_20[122]}
   );
   gpc1_1 gpc1711 (
      {stage0_20[249]},
      {stage1_20[123]}
   );
   gpc1_1 gpc1712 (
      {stage0_20[250]},
      {stage1_20[124]}
   );
   gpc1_1 gpc1713 (
      {stage0_20[251]},
      {stage1_20[125]}
   );
   gpc1_1 gpc1714 (
      {stage0_20[252]},
      {stage1_20[126]}
   );
   gpc1_1 gpc1715 (
      {stage0_20[253]},
      {stage1_20[127]}
   );
   gpc1_1 gpc1716 (
      {stage0_20[254]},
      {stage1_20[128]}
   );
   gpc1_1 gpc1717 (
      {stage0_20[255]},
      {stage1_20[129]}
   );
   gpc1_1 gpc1718 (
      {stage0_21[252]},
      {stage1_21[104]}
   );
   gpc1_1 gpc1719 (
      {stage0_21[253]},
      {stage1_21[105]}
   );
   gpc1_1 gpc1720 (
      {stage0_21[254]},
      {stage1_21[106]}
   );
   gpc1_1 gpc1721 (
      {stage0_21[255]},
      {stage1_21[107]}
   );
   gpc1_1 gpc1722 (
      {stage0_22[252]},
      {stage1_22[88]}
   );
   gpc1_1 gpc1723 (
      {stage0_22[253]},
      {stage1_22[89]}
   );
   gpc1_1 gpc1724 (
      {stage0_22[254]},
      {stage1_22[90]}
   );
   gpc1_1 gpc1725 (
      {stage0_22[255]},
      {stage1_22[91]}
   );
   gpc1_1 gpc1726 (
      {stage0_23[226]},
      {stage1_23[99]}
   );
   gpc1_1 gpc1727 (
      {stage0_23[227]},
      {stage1_23[100]}
   );
   gpc1_1 gpc1728 (
      {stage0_23[228]},
      {stage1_23[101]}
   );
   gpc1_1 gpc1729 (
      {stage0_23[229]},
      {stage1_23[102]}
   );
   gpc1_1 gpc1730 (
      {stage0_23[230]},
      {stage1_23[103]}
   );
   gpc1_1 gpc1731 (
      {stage0_23[231]},
      {stage1_23[104]}
   );
   gpc1_1 gpc1732 (
      {stage0_23[232]},
      {stage1_23[105]}
   );
   gpc1_1 gpc1733 (
      {stage0_23[233]},
      {stage1_23[106]}
   );
   gpc1_1 gpc1734 (
      {stage0_23[234]},
      {stage1_23[107]}
   );
   gpc1_1 gpc1735 (
      {stage0_23[235]},
      {stage1_23[108]}
   );
   gpc1_1 gpc1736 (
      {stage0_23[236]},
      {stage1_23[109]}
   );
   gpc1_1 gpc1737 (
      {stage0_23[237]},
      {stage1_23[110]}
   );
   gpc1_1 gpc1738 (
      {stage0_23[238]},
      {stage1_23[111]}
   );
   gpc1_1 gpc1739 (
      {stage0_23[239]},
      {stage1_23[112]}
   );
   gpc1_1 gpc1740 (
      {stage0_23[240]},
      {stage1_23[113]}
   );
   gpc1_1 gpc1741 (
      {stage0_23[241]},
      {stage1_23[114]}
   );
   gpc1_1 gpc1742 (
      {stage0_23[242]},
      {stage1_23[115]}
   );
   gpc1_1 gpc1743 (
      {stage0_23[243]},
      {stage1_23[116]}
   );
   gpc1_1 gpc1744 (
      {stage0_23[244]},
      {stage1_23[117]}
   );
   gpc1_1 gpc1745 (
      {stage0_23[245]},
      {stage1_23[118]}
   );
   gpc1_1 gpc1746 (
      {stage0_23[246]},
      {stage1_23[119]}
   );
   gpc1_1 gpc1747 (
      {stage0_23[247]},
      {stage1_23[120]}
   );
   gpc1_1 gpc1748 (
      {stage0_23[248]},
      {stage1_23[121]}
   );
   gpc1_1 gpc1749 (
      {stage0_23[249]},
      {stage1_23[122]}
   );
   gpc1_1 gpc1750 (
      {stage0_23[250]},
      {stage1_23[123]}
   );
   gpc1_1 gpc1751 (
      {stage0_23[251]},
      {stage1_23[124]}
   );
   gpc1_1 gpc1752 (
      {stage0_23[252]},
      {stage1_23[125]}
   );
   gpc1_1 gpc1753 (
      {stage0_23[253]},
      {stage1_23[126]}
   );
   gpc1_1 gpc1754 (
      {stage0_23[254]},
      {stage1_23[127]}
   );
   gpc1_1 gpc1755 (
      {stage0_23[255]},
      {stage1_23[128]}
   );
   gpc1_1 gpc1756 (
      {stage0_24[231]},
      {stage1_24[115]}
   );
   gpc1_1 gpc1757 (
      {stage0_24[232]},
      {stage1_24[116]}
   );
   gpc1_1 gpc1758 (
      {stage0_24[233]},
      {stage1_24[117]}
   );
   gpc1_1 gpc1759 (
      {stage0_24[234]},
      {stage1_24[118]}
   );
   gpc1_1 gpc1760 (
      {stage0_24[235]},
      {stage1_24[119]}
   );
   gpc1_1 gpc1761 (
      {stage0_24[236]},
      {stage1_24[120]}
   );
   gpc1_1 gpc1762 (
      {stage0_24[237]},
      {stage1_24[121]}
   );
   gpc1_1 gpc1763 (
      {stage0_24[238]},
      {stage1_24[122]}
   );
   gpc1_1 gpc1764 (
      {stage0_24[239]},
      {stage1_24[123]}
   );
   gpc1_1 gpc1765 (
      {stage0_24[240]},
      {stage1_24[124]}
   );
   gpc1_1 gpc1766 (
      {stage0_24[241]},
      {stage1_24[125]}
   );
   gpc1_1 gpc1767 (
      {stage0_24[242]},
      {stage1_24[126]}
   );
   gpc1_1 gpc1768 (
      {stage0_24[243]},
      {stage1_24[127]}
   );
   gpc1_1 gpc1769 (
      {stage0_24[244]},
      {stage1_24[128]}
   );
   gpc1_1 gpc1770 (
      {stage0_24[245]},
      {stage1_24[129]}
   );
   gpc1_1 gpc1771 (
      {stage0_24[246]},
      {stage1_24[130]}
   );
   gpc1_1 gpc1772 (
      {stage0_24[247]},
      {stage1_24[131]}
   );
   gpc1_1 gpc1773 (
      {stage0_24[248]},
      {stage1_24[132]}
   );
   gpc1_1 gpc1774 (
      {stage0_24[249]},
      {stage1_24[133]}
   );
   gpc1_1 gpc1775 (
      {stage0_24[250]},
      {stage1_24[134]}
   );
   gpc1_1 gpc1776 (
      {stage0_24[251]},
      {stage1_24[135]}
   );
   gpc1_1 gpc1777 (
      {stage0_24[252]},
      {stage1_24[136]}
   );
   gpc1_1 gpc1778 (
      {stage0_24[253]},
      {stage1_24[137]}
   );
   gpc1_1 gpc1779 (
      {stage0_24[254]},
      {stage1_24[138]}
   );
   gpc1_1 gpc1780 (
      {stage0_24[255]},
      {stage1_24[139]}
   );
   gpc1_1 gpc1781 (
      {stage0_25[245]},
      {stage1_25[99]}
   );
   gpc1_1 gpc1782 (
      {stage0_25[246]},
      {stage1_25[100]}
   );
   gpc1_1 gpc1783 (
      {stage0_25[247]},
      {stage1_25[101]}
   );
   gpc1_1 gpc1784 (
      {stage0_25[248]},
      {stage1_25[102]}
   );
   gpc1_1 gpc1785 (
      {stage0_25[249]},
      {stage1_25[103]}
   );
   gpc1_1 gpc1786 (
      {stage0_25[250]},
      {stage1_25[104]}
   );
   gpc1_1 gpc1787 (
      {stage0_25[251]},
      {stage1_25[105]}
   );
   gpc1_1 gpc1788 (
      {stage0_25[252]},
      {stage1_25[106]}
   );
   gpc1_1 gpc1789 (
      {stage0_25[253]},
      {stage1_25[107]}
   );
   gpc1_1 gpc1790 (
      {stage0_25[254]},
      {stage1_25[108]}
   );
   gpc1_1 gpc1791 (
      {stage0_25[255]},
      {stage1_25[109]}
   );
   gpc1_1 gpc1792 (
      {stage0_26[195]},
      {stage1_26[80]}
   );
   gpc1_1 gpc1793 (
      {stage0_26[196]},
      {stage1_26[81]}
   );
   gpc1_1 gpc1794 (
      {stage0_26[197]},
      {stage1_26[82]}
   );
   gpc1_1 gpc1795 (
      {stage0_26[198]},
      {stage1_26[83]}
   );
   gpc1_1 gpc1796 (
      {stage0_26[199]},
      {stage1_26[84]}
   );
   gpc1_1 gpc1797 (
      {stage0_26[200]},
      {stage1_26[85]}
   );
   gpc1_1 gpc1798 (
      {stage0_26[201]},
      {stage1_26[86]}
   );
   gpc1_1 gpc1799 (
      {stage0_26[202]},
      {stage1_26[87]}
   );
   gpc1_1 gpc1800 (
      {stage0_26[203]},
      {stage1_26[88]}
   );
   gpc1_1 gpc1801 (
      {stage0_26[204]},
      {stage1_26[89]}
   );
   gpc1_1 gpc1802 (
      {stage0_26[205]},
      {stage1_26[90]}
   );
   gpc1_1 gpc1803 (
      {stage0_26[206]},
      {stage1_26[91]}
   );
   gpc1_1 gpc1804 (
      {stage0_26[207]},
      {stage1_26[92]}
   );
   gpc1_1 gpc1805 (
      {stage0_26[208]},
      {stage1_26[93]}
   );
   gpc1_1 gpc1806 (
      {stage0_26[209]},
      {stage1_26[94]}
   );
   gpc1_1 gpc1807 (
      {stage0_26[210]},
      {stage1_26[95]}
   );
   gpc1_1 gpc1808 (
      {stage0_26[211]},
      {stage1_26[96]}
   );
   gpc1_1 gpc1809 (
      {stage0_26[212]},
      {stage1_26[97]}
   );
   gpc1_1 gpc1810 (
      {stage0_26[213]},
      {stage1_26[98]}
   );
   gpc1_1 gpc1811 (
      {stage0_26[214]},
      {stage1_26[99]}
   );
   gpc1_1 gpc1812 (
      {stage0_26[215]},
      {stage1_26[100]}
   );
   gpc1_1 gpc1813 (
      {stage0_26[216]},
      {stage1_26[101]}
   );
   gpc1_1 gpc1814 (
      {stage0_26[217]},
      {stage1_26[102]}
   );
   gpc1_1 gpc1815 (
      {stage0_26[218]},
      {stage1_26[103]}
   );
   gpc1_1 gpc1816 (
      {stage0_26[219]},
      {stage1_26[104]}
   );
   gpc1_1 gpc1817 (
      {stage0_26[220]},
      {stage1_26[105]}
   );
   gpc1_1 gpc1818 (
      {stage0_26[221]},
      {stage1_26[106]}
   );
   gpc1_1 gpc1819 (
      {stage0_26[222]},
      {stage1_26[107]}
   );
   gpc1_1 gpc1820 (
      {stage0_26[223]},
      {stage1_26[108]}
   );
   gpc1_1 gpc1821 (
      {stage0_26[224]},
      {stage1_26[109]}
   );
   gpc1_1 gpc1822 (
      {stage0_26[225]},
      {stage1_26[110]}
   );
   gpc1_1 gpc1823 (
      {stage0_26[226]},
      {stage1_26[111]}
   );
   gpc1_1 gpc1824 (
      {stage0_26[227]},
      {stage1_26[112]}
   );
   gpc1_1 gpc1825 (
      {stage0_26[228]},
      {stage1_26[113]}
   );
   gpc1_1 gpc1826 (
      {stage0_26[229]},
      {stage1_26[114]}
   );
   gpc1_1 gpc1827 (
      {stage0_26[230]},
      {stage1_26[115]}
   );
   gpc1_1 gpc1828 (
      {stage0_26[231]},
      {stage1_26[116]}
   );
   gpc1_1 gpc1829 (
      {stage0_26[232]},
      {stage1_26[117]}
   );
   gpc1_1 gpc1830 (
      {stage0_26[233]},
      {stage1_26[118]}
   );
   gpc1_1 gpc1831 (
      {stage0_26[234]},
      {stage1_26[119]}
   );
   gpc1_1 gpc1832 (
      {stage0_26[235]},
      {stage1_26[120]}
   );
   gpc1_1 gpc1833 (
      {stage0_26[236]},
      {stage1_26[121]}
   );
   gpc1_1 gpc1834 (
      {stage0_26[237]},
      {stage1_26[122]}
   );
   gpc1_1 gpc1835 (
      {stage0_26[238]},
      {stage1_26[123]}
   );
   gpc1_1 gpc1836 (
      {stage0_26[239]},
      {stage1_26[124]}
   );
   gpc1_1 gpc1837 (
      {stage0_26[240]},
      {stage1_26[125]}
   );
   gpc1_1 gpc1838 (
      {stage0_26[241]},
      {stage1_26[126]}
   );
   gpc1_1 gpc1839 (
      {stage0_26[242]},
      {stage1_26[127]}
   );
   gpc1_1 gpc1840 (
      {stage0_26[243]},
      {stage1_26[128]}
   );
   gpc1_1 gpc1841 (
      {stage0_26[244]},
      {stage1_26[129]}
   );
   gpc1_1 gpc1842 (
      {stage0_26[245]},
      {stage1_26[130]}
   );
   gpc1_1 gpc1843 (
      {stage0_26[246]},
      {stage1_26[131]}
   );
   gpc1_1 gpc1844 (
      {stage0_26[247]},
      {stage1_26[132]}
   );
   gpc1_1 gpc1845 (
      {stage0_26[248]},
      {stage1_26[133]}
   );
   gpc1_1 gpc1846 (
      {stage0_26[249]},
      {stage1_26[134]}
   );
   gpc1_1 gpc1847 (
      {stage0_26[250]},
      {stage1_26[135]}
   );
   gpc1_1 gpc1848 (
      {stage0_26[251]},
      {stage1_26[136]}
   );
   gpc1_1 gpc1849 (
      {stage0_26[252]},
      {stage1_26[137]}
   );
   gpc1_1 gpc1850 (
      {stage0_26[253]},
      {stage1_26[138]}
   );
   gpc1_1 gpc1851 (
      {stage0_26[254]},
      {stage1_26[139]}
   );
   gpc1_1 gpc1852 (
      {stage0_26[255]},
      {stage1_26[140]}
   );
   gpc1_1 gpc1853 (
      {stage0_27[224]},
      {stage1_27[87]}
   );
   gpc1_1 gpc1854 (
      {stage0_27[225]},
      {stage1_27[88]}
   );
   gpc1_1 gpc1855 (
      {stage0_27[226]},
      {stage1_27[89]}
   );
   gpc1_1 gpc1856 (
      {stage0_27[227]},
      {stage1_27[90]}
   );
   gpc1_1 gpc1857 (
      {stage0_27[228]},
      {stage1_27[91]}
   );
   gpc1_1 gpc1858 (
      {stage0_27[229]},
      {stage1_27[92]}
   );
   gpc1_1 gpc1859 (
      {stage0_27[230]},
      {stage1_27[93]}
   );
   gpc1_1 gpc1860 (
      {stage0_27[231]},
      {stage1_27[94]}
   );
   gpc1_1 gpc1861 (
      {stage0_27[232]},
      {stage1_27[95]}
   );
   gpc1_1 gpc1862 (
      {stage0_27[233]},
      {stage1_27[96]}
   );
   gpc1_1 gpc1863 (
      {stage0_27[234]},
      {stage1_27[97]}
   );
   gpc1_1 gpc1864 (
      {stage0_27[235]},
      {stage1_27[98]}
   );
   gpc1_1 gpc1865 (
      {stage0_27[236]},
      {stage1_27[99]}
   );
   gpc1_1 gpc1866 (
      {stage0_27[237]},
      {stage1_27[100]}
   );
   gpc1_1 gpc1867 (
      {stage0_27[238]},
      {stage1_27[101]}
   );
   gpc1_1 gpc1868 (
      {stage0_27[239]},
      {stage1_27[102]}
   );
   gpc1_1 gpc1869 (
      {stage0_27[240]},
      {stage1_27[103]}
   );
   gpc1_1 gpc1870 (
      {stage0_27[241]},
      {stage1_27[104]}
   );
   gpc1_1 gpc1871 (
      {stage0_27[242]},
      {stage1_27[105]}
   );
   gpc1_1 gpc1872 (
      {stage0_27[243]},
      {stage1_27[106]}
   );
   gpc1_1 gpc1873 (
      {stage0_27[244]},
      {stage1_27[107]}
   );
   gpc1_1 gpc1874 (
      {stage0_27[245]},
      {stage1_27[108]}
   );
   gpc1_1 gpc1875 (
      {stage0_27[246]},
      {stage1_27[109]}
   );
   gpc1_1 gpc1876 (
      {stage0_27[247]},
      {stage1_27[110]}
   );
   gpc1_1 gpc1877 (
      {stage0_27[248]},
      {stage1_27[111]}
   );
   gpc1_1 gpc1878 (
      {stage0_27[249]},
      {stage1_27[112]}
   );
   gpc1_1 gpc1879 (
      {stage0_27[250]},
      {stage1_27[113]}
   );
   gpc1_1 gpc1880 (
      {stage0_27[251]},
      {stage1_27[114]}
   );
   gpc1_1 gpc1881 (
      {stage0_27[252]},
      {stage1_27[115]}
   );
   gpc1_1 gpc1882 (
      {stage0_27[253]},
      {stage1_27[116]}
   );
   gpc1_1 gpc1883 (
      {stage0_27[254]},
      {stage1_27[117]}
   );
   gpc1_1 gpc1884 (
      {stage0_27[255]},
      {stage1_27[118]}
   );
   gpc1_1 gpc1885 (
      {stage0_28[235]},
      {stage1_28[106]}
   );
   gpc1_1 gpc1886 (
      {stage0_28[236]},
      {stage1_28[107]}
   );
   gpc1_1 gpc1887 (
      {stage0_28[237]},
      {stage1_28[108]}
   );
   gpc1_1 gpc1888 (
      {stage0_28[238]},
      {stage1_28[109]}
   );
   gpc1_1 gpc1889 (
      {stage0_28[239]},
      {stage1_28[110]}
   );
   gpc1_1 gpc1890 (
      {stage0_28[240]},
      {stage1_28[111]}
   );
   gpc1_1 gpc1891 (
      {stage0_28[241]},
      {stage1_28[112]}
   );
   gpc1_1 gpc1892 (
      {stage0_28[242]},
      {stage1_28[113]}
   );
   gpc1_1 gpc1893 (
      {stage0_28[243]},
      {stage1_28[114]}
   );
   gpc1_1 gpc1894 (
      {stage0_28[244]},
      {stage1_28[115]}
   );
   gpc1_1 gpc1895 (
      {stage0_28[245]},
      {stage1_28[116]}
   );
   gpc1_1 gpc1896 (
      {stage0_28[246]},
      {stage1_28[117]}
   );
   gpc1_1 gpc1897 (
      {stage0_28[247]},
      {stage1_28[118]}
   );
   gpc1_1 gpc1898 (
      {stage0_28[248]},
      {stage1_28[119]}
   );
   gpc1_1 gpc1899 (
      {stage0_28[249]},
      {stage1_28[120]}
   );
   gpc1_1 gpc1900 (
      {stage0_28[250]},
      {stage1_28[121]}
   );
   gpc1_1 gpc1901 (
      {stage0_28[251]},
      {stage1_28[122]}
   );
   gpc1_1 gpc1902 (
      {stage0_28[252]},
      {stage1_28[123]}
   );
   gpc1_1 gpc1903 (
      {stage0_28[253]},
      {stage1_28[124]}
   );
   gpc1_1 gpc1904 (
      {stage0_28[254]},
      {stage1_28[125]}
   );
   gpc1_1 gpc1905 (
      {stage0_28[255]},
      {stage1_28[126]}
   );
   gpc1_1 gpc1906 (
      {stage0_29[247]},
      {stage1_29[101]}
   );
   gpc1_1 gpc1907 (
      {stage0_29[248]},
      {stage1_29[102]}
   );
   gpc1_1 gpc1908 (
      {stage0_29[249]},
      {stage1_29[103]}
   );
   gpc1_1 gpc1909 (
      {stage0_29[250]},
      {stage1_29[104]}
   );
   gpc1_1 gpc1910 (
      {stage0_29[251]},
      {stage1_29[105]}
   );
   gpc1_1 gpc1911 (
      {stage0_29[252]},
      {stage1_29[106]}
   );
   gpc1_1 gpc1912 (
      {stage0_29[253]},
      {stage1_29[107]}
   );
   gpc1_1 gpc1913 (
      {stage0_29[254]},
      {stage1_29[108]}
   );
   gpc1_1 gpc1914 (
      {stage0_29[255]},
      {stage1_29[109]}
   );
   gpc1_1 gpc1915 (
      {stage0_30[254]},
      {stage1_30[89]}
   );
   gpc1_1 gpc1916 (
      {stage0_30[255]},
      {stage1_30[90]}
   );
   gpc1_1 gpc1917 (
      {stage0_31[243]},
      {stage1_31[102]}
   );
   gpc1_1 gpc1918 (
      {stage0_31[244]},
      {stage1_31[103]}
   );
   gpc1_1 gpc1919 (
      {stage0_31[245]},
      {stage1_31[104]}
   );
   gpc1_1 gpc1920 (
      {stage0_31[246]},
      {stage1_31[105]}
   );
   gpc1_1 gpc1921 (
      {stage0_31[247]},
      {stage1_31[106]}
   );
   gpc1_1 gpc1922 (
      {stage0_31[248]},
      {stage1_31[107]}
   );
   gpc1_1 gpc1923 (
      {stage0_31[249]},
      {stage1_31[108]}
   );
   gpc1_1 gpc1924 (
      {stage0_31[250]},
      {stage1_31[109]}
   );
   gpc1_1 gpc1925 (
      {stage0_31[251]},
      {stage1_31[110]}
   );
   gpc1_1 gpc1926 (
      {stage0_31[252]},
      {stage1_31[111]}
   );
   gpc1_1 gpc1927 (
      {stage0_31[253]},
      {stage1_31[112]}
   );
   gpc1_1 gpc1928 (
      {stage0_31[254]},
      {stage1_31[113]}
   );
   gpc1_1 gpc1929 (
      {stage0_31[255]},
      {stage1_31[114]}
   );
   gpc1_1 gpc1930 (
      {stage0_33[252]},
      {stage1_33[107]}
   );
   gpc1_1 gpc1931 (
      {stage0_33[253]},
      {stage1_33[108]}
   );
   gpc1_1 gpc1932 (
      {stage0_33[254]},
      {stage1_33[109]}
   );
   gpc1_1 gpc1933 (
      {stage0_33[255]},
      {stage1_33[110]}
   );
   gpc1_1 gpc1934 (
      {stage0_34[249]},
      {stage1_34[97]}
   );
   gpc1_1 gpc1935 (
      {stage0_34[250]},
      {stage1_34[98]}
   );
   gpc1_1 gpc1936 (
      {stage0_34[251]},
      {stage1_34[99]}
   );
   gpc1_1 gpc1937 (
      {stage0_34[252]},
      {stage1_34[100]}
   );
   gpc1_1 gpc1938 (
      {stage0_34[253]},
      {stage1_34[101]}
   );
   gpc1_1 gpc1939 (
      {stage0_34[254]},
      {stage1_34[102]}
   );
   gpc1_1 gpc1940 (
      {stage0_34[255]},
      {stage1_34[103]}
   );
   gpc1_1 gpc1941 (
      {stage0_35[236]},
      {stage1_35[99]}
   );
   gpc1_1 gpc1942 (
      {stage0_35[237]},
      {stage1_35[100]}
   );
   gpc1_1 gpc1943 (
      {stage0_35[238]},
      {stage1_35[101]}
   );
   gpc1_1 gpc1944 (
      {stage0_35[239]},
      {stage1_35[102]}
   );
   gpc1_1 gpc1945 (
      {stage0_35[240]},
      {stage1_35[103]}
   );
   gpc1_1 gpc1946 (
      {stage0_35[241]},
      {stage1_35[104]}
   );
   gpc1_1 gpc1947 (
      {stage0_35[242]},
      {stage1_35[105]}
   );
   gpc1_1 gpc1948 (
      {stage0_35[243]},
      {stage1_35[106]}
   );
   gpc1_1 gpc1949 (
      {stage0_35[244]},
      {stage1_35[107]}
   );
   gpc1_1 gpc1950 (
      {stage0_35[245]},
      {stage1_35[108]}
   );
   gpc1_1 gpc1951 (
      {stage0_35[246]},
      {stage1_35[109]}
   );
   gpc1_1 gpc1952 (
      {stage0_35[247]},
      {stage1_35[110]}
   );
   gpc1_1 gpc1953 (
      {stage0_35[248]},
      {stage1_35[111]}
   );
   gpc1_1 gpc1954 (
      {stage0_35[249]},
      {stage1_35[112]}
   );
   gpc1_1 gpc1955 (
      {stage0_35[250]},
      {stage1_35[113]}
   );
   gpc1_1 gpc1956 (
      {stage0_35[251]},
      {stage1_35[114]}
   );
   gpc1_1 gpc1957 (
      {stage0_35[252]},
      {stage1_35[115]}
   );
   gpc1_1 gpc1958 (
      {stage0_35[253]},
      {stage1_35[116]}
   );
   gpc1_1 gpc1959 (
      {stage0_35[254]},
      {stage1_35[117]}
   );
   gpc1_1 gpc1960 (
      {stage0_35[255]},
      {stage1_35[118]}
   );
   gpc1_1 gpc1961 (
      {stage0_36[212]},
      {stage1_36[101]}
   );
   gpc1_1 gpc1962 (
      {stage0_36[213]},
      {stage1_36[102]}
   );
   gpc1_1 gpc1963 (
      {stage0_36[214]},
      {stage1_36[103]}
   );
   gpc1_1 gpc1964 (
      {stage0_36[215]},
      {stage1_36[104]}
   );
   gpc1_1 gpc1965 (
      {stage0_36[216]},
      {stage1_36[105]}
   );
   gpc1_1 gpc1966 (
      {stage0_36[217]},
      {stage1_36[106]}
   );
   gpc1_1 gpc1967 (
      {stage0_36[218]},
      {stage1_36[107]}
   );
   gpc1_1 gpc1968 (
      {stage0_36[219]},
      {stage1_36[108]}
   );
   gpc1_1 gpc1969 (
      {stage0_36[220]},
      {stage1_36[109]}
   );
   gpc1_1 gpc1970 (
      {stage0_36[221]},
      {stage1_36[110]}
   );
   gpc1_1 gpc1971 (
      {stage0_36[222]},
      {stage1_36[111]}
   );
   gpc1_1 gpc1972 (
      {stage0_36[223]},
      {stage1_36[112]}
   );
   gpc1_1 gpc1973 (
      {stage0_36[224]},
      {stage1_36[113]}
   );
   gpc1_1 gpc1974 (
      {stage0_36[225]},
      {stage1_36[114]}
   );
   gpc1_1 gpc1975 (
      {stage0_36[226]},
      {stage1_36[115]}
   );
   gpc1_1 gpc1976 (
      {stage0_36[227]},
      {stage1_36[116]}
   );
   gpc1_1 gpc1977 (
      {stage0_36[228]},
      {stage1_36[117]}
   );
   gpc1_1 gpc1978 (
      {stage0_36[229]},
      {stage1_36[118]}
   );
   gpc1_1 gpc1979 (
      {stage0_36[230]},
      {stage1_36[119]}
   );
   gpc1_1 gpc1980 (
      {stage0_36[231]},
      {stage1_36[120]}
   );
   gpc1_1 gpc1981 (
      {stage0_36[232]},
      {stage1_36[121]}
   );
   gpc1_1 gpc1982 (
      {stage0_36[233]},
      {stage1_36[122]}
   );
   gpc1_1 gpc1983 (
      {stage0_36[234]},
      {stage1_36[123]}
   );
   gpc1_1 gpc1984 (
      {stage0_36[235]},
      {stage1_36[124]}
   );
   gpc1_1 gpc1985 (
      {stage0_36[236]},
      {stage1_36[125]}
   );
   gpc1_1 gpc1986 (
      {stage0_36[237]},
      {stage1_36[126]}
   );
   gpc1_1 gpc1987 (
      {stage0_36[238]},
      {stage1_36[127]}
   );
   gpc1_1 gpc1988 (
      {stage0_36[239]},
      {stage1_36[128]}
   );
   gpc1_1 gpc1989 (
      {stage0_36[240]},
      {stage1_36[129]}
   );
   gpc1_1 gpc1990 (
      {stage0_36[241]},
      {stage1_36[130]}
   );
   gpc1_1 gpc1991 (
      {stage0_36[242]},
      {stage1_36[131]}
   );
   gpc1_1 gpc1992 (
      {stage0_36[243]},
      {stage1_36[132]}
   );
   gpc1_1 gpc1993 (
      {stage0_36[244]},
      {stage1_36[133]}
   );
   gpc1_1 gpc1994 (
      {stage0_36[245]},
      {stage1_36[134]}
   );
   gpc1_1 gpc1995 (
      {stage0_36[246]},
      {stage1_36[135]}
   );
   gpc1_1 gpc1996 (
      {stage0_36[247]},
      {stage1_36[136]}
   );
   gpc1_1 gpc1997 (
      {stage0_36[248]},
      {stage1_36[137]}
   );
   gpc1_1 gpc1998 (
      {stage0_36[249]},
      {stage1_36[138]}
   );
   gpc1_1 gpc1999 (
      {stage0_36[250]},
      {stage1_36[139]}
   );
   gpc1_1 gpc2000 (
      {stage0_36[251]},
      {stage1_36[140]}
   );
   gpc1_1 gpc2001 (
      {stage0_36[252]},
      {stage1_36[141]}
   );
   gpc1_1 gpc2002 (
      {stage0_36[253]},
      {stage1_36[142]}
   );
   gpc1_1 gpc2003 (
      {stage0_36[254]},
      {stage1_36[143]}
   );
   gpc1_1 gpc2004 (
      {stage0_36[255]},
      {stage1_36[144]}
   );
   gpc1_1 gpc2005 (
      {stage0_37[252]},
      {stage1_37[101]}
   );
   gpc1_1 gpc2006 (
      {stage0_37[253]},
      {stage1_37[102]}
   );
   gpc1_1 gpc2007 (
      {stage0_37[254]},
      {stage1_37[103]}
   );
   gpc1_1 gpc2008 (
      {stage0_37[255]},
      {stage1_37[104]}
   );
   gpc1_1 gpc2009 (
      {stage0_38[217]},
      {stage1_38[98]}
   );
   gpc1_1 gpc2010 (
      {stage0_38[218]},
      {stage1_38[99]}
   );
   gpc1_1 gpc2011 (
      {stage0_38[219]},
      {stage1_38[100]}
   );
   gpc1_1 gpc2012 (
      {stage0_38[220]},
      {stage1_38[101]}
   );
   gpc1_1 gpc2013 (
      {stage0_38[221]},
      {stage1_38[102]}
   );
   gpc1_1 gpc2014 (
      {stage0_38[222]},
      {stage1_38[103]}
   );
   gpc1_1 gpc2015 (
      {stage0_38[223]},
      {stage1_38[104]}
   );
   gpc1_1 gpc2016 (
      {stage0_38[224]},
      {stage1_38[105]}
   );
   gpc1_1 gpc2017 (
      {stage0_38[225]},
      {stage1_38[106]}
   );
   gpc1_1 gpc2018 (
      {stage0_38[226]},
      {stage1_38[107]}
   );
   gpc1_1 gpc2019 (
      {stage0_38[227]},
      {stage1_38[108]}
   );
   gpc1_1 gpc2020 (
      {stage0_38[228]},
      {stage1_38[109]}
   );
   gpc1_1 gpc2021 (
      {stage0_38[229]},
      {stage1_38[110]}
   );
   gpc1_1 gpc2022 (
      {stage0_38[230]},
      {stage1_38[111]}
   );
   gpc1_1 gpc2023 (
      {stage0_38[231]},
      {stage1_38[112]}
   );
   gpc1_1 gpc2024 (
      {stage0_38[232]},
      {stage1_38[113]}
   );
   gpc1_1 gpc2025 (
      {stage0_38[233]},
      {stage1_38[114]}
   );
   gpc1_1 gpc2026 (
      {stage0_38[234]},
      {stage1_38[115]}
   );
   gpc1_1 gpc2027 (
      {stage0_38[235]},
      {stage1_38[116]}
   );
   gpc1_1 gpc2028 (
      {stage0_38[236]},
      {stage1_38[117]}
   );
   gpc1_1 gpc2029 (
      {stage0_38[237]},
      {stage1_38[118]}
   );
   gpc1_1 gpc2030 (
      {stage0_38[238]},
      {stage1_38[119]}
   );
   gpc1_1 gpc2031 (
      {stage0_38[239]},
      {stage1_38[120]}
   );
   gpc1_1 gpc2032 (
      {stage0_38[240]},
      {stage1_38[121]}
   );
   gpc1_1 gpc2033 (
      {stage0_38[241]},
      {stage1_38[122]}
   );
   gpc1_1 gpc2034 (
      {stage0_38[242]},
      {stage1_38[123]}
   );
   gpc1_1 gpc2035 (
      {stage0_38[243]},
      {stage1_38[124]}
   );
   gpc1_1 gpc2036 (
      {stage0_38[244]},
      {stage1_38[125]}
   );
   gpc1_1 gpc2037 (
      {stage0_38[245]},
      {stage1_38[126]}
   );
   gpc1_1 gpc2038 (
      {stage0_38[246]},
      {stage1_38[127]}
   );
   gpc1_1 gpc2039 (
      {stage0_38[247]},
      {stage1_38[128]}
   );
   gpc1_1 gpc2040 (
      {stage0_38[248]},
      {stage1_38[129]}
   );
   gpc1_1 gpc2041 (
      {stage0_38[249]},
      {stage1_38[130]}
   );
   gpc1_1 gpc2042 (
      {stage0_38[250]},
      {stage1_38[131]}
   );
   gpc1_1 gpc2043 (
      {stage0_38[251]},
      {stage1_38[132]}
   );
   gpc1_1 gpc2044 (
      {stage0_38[252]},
      {stage1_38[133]}
   );
   gpc1_1 gpc2045 (
      {stage0_38[253]},
      {stage1_38[134]}
   );
   gpc1_1 gpc2046 (
      {stage0_38[254]},
      {stage1_38[135]}
   );
   gpc1_1 gpc2047 (
      {stage0_38[255]},
      {stage1_38[136]}
   );
   gpc1_1 gpc2048 (
      {stage0_39[218]},
      {stage1_39[87]}
   );
   gpc1_1 gpc2049 (
      {stage0_39[219]},
      {stage1_39[88]}
   );
   gpc1_1 gpc2050 (
      {stage0_39[220]},
      {stage1_39[89]}
   );
   gpc1_1 gpc2051 (
      {stage0_39[221]},
      {stage1_39[90]}
   );
   gpc1_1 gpc2052 (
      {stage0_39[222]},
      {stage1_39[91]}
   );
   gpc1_1 gpc2053 (
      {stage0_39[223]},
      {stage1_39[92]}
   );
   gpc1_1 gpc2054 (
      {stage0_39[224]},
      {stage1_39[93]}
   );
   gpc1_1 gpc2055 (
      {stage0_39[225]},
      {stage1_39[94]}
   );
   gpc1_1 gpc2056 (
      {stage0_39[226]},
      {stage1_39[95]}
   );
   gpc1_1 gpc2057 (
      {stage0_39[227]},
      {stage1_39[96]}
   );
   gpc1_1 gpc2058 (
      {stage0_39[228]},
      {stage1_39[97]}
   );
   gpc1_1 gpc2059 (
      {stage0_39[229]},
      {stage1_39[98]}
   );
   gpc1_1 gpc2060 (
      {stage0_39[230]},
      {stage1_39[99]}
   );
   gpc1_1 gpc2061 (
      {stage0_39[231]},
      {stage1_39[100]}
   );
   gpc1_1 gpc2062 (
      {stage0_39[232]},
      {stage1_39[101]}
   );
   gpc1_1 gpc2063 (
      {stage0_39[233]},
      {stage1_39[102]}
   );
   gpc1_1 gpc2064 (
      {stage0_39[234]},
      {stage1_39[103]}
   );
   gpc1_1 gpc2065 (
      {stage0_39[235]},
      {stage1_39[104]}
   );
   gpc1_1 gpc2066 (
      {stage0_39[236]},
      {stage1_39[105]}
   );
   gpc1_1 gpc2067 (
      {stage0_39[237]},
      {stage1_39[106]}
   );
   gpc1_1 gpc2068 (
      {stage0_39[238]},
      {stage1_39[107]}
   );
   gpc1_1 gpc2069 (
      {stage0_39[239]},
      {stage1_39[108]}
   );
   gpc1_1 gpc2070 (
      {stage0_39[240]},
      {stage1_39[109]}
   );
   gpc1_1 gpc2071 (
      {stage0_39[241]},
      {stage1_39[110]}
   );
   gpc1_1 gpc2072 (
      {stage0_39[242]},
      {stage1_39[111]}
   );
   gpc1_1 gpc2073 (
      {stage0_39[243]},
      {stage1_39[112]}
   );
   gpc1_1 gpc2074 (
      {stage0_39[244]},
      {stage1_39[113]}
   );
   gpc1_1 gpc2075 (
      {stage0_39[245]},
      {stage1_39[114]}
   );
   gpc1_1 gpc2076 (
      {stage0_39[246]},
      {stage1_39[115]}
   );
   gpc1_1 gpc2077 (
      {stage0_39[247]},
      {stage1_39[116]}
   );
   gpc1_1 gpc2078 (
      {stage0_39[248]},
      {stage1_39[117]}
   );
   gpc1_1 gpc2079 (
      {stage0_39[249]},
      {stage1_39[118]}
   );
   gpc1_1 gpc2080 (
      {stage0_39[250]},
      {stage1_39[119]}
   );
   gpc1_1 gpc2081 (
      {stage0_39[251]},
      {stage1_39[120]}
   );
   gpc1_1 gpc2082 (
      {stage0_39[252]},
      {stage1_39[121]}
   );
   gpc1_1 gpc2083 (
      {stage0_39[253]},
      {stage1_39[122]}
   );
   gpc1_1 gpc2084 (
      {stage0_39[254]},
      {stage1_39[123]}
   );
   gpc1_1 gpc2085 (
      {stage0_39[255]},
      {stage1_39[124]}
   );
   gpc1_1 gpc2086 (
      {stage0_41[224]},
      {stage1_41[111]}
   );
   gpc1_1 gpc2087 (
      {stage0_41[225]},
      {stage1_41[112]}
   );
   gpc1_1 gpc2088 (
      {stage0_41[226]},
      {stage1_41[113]}
   );
   gpc1_1 gpc2089 (
      {stage0_41[227]},
      {stage1_41[114]}
   );
   gpc1_1 gpc2090 (
      {stage0_41[228]},
      {stage1_41[115]}
   );
   gpc1_1 gpc2091 (
      {stage0_41[229]},
      {stage1_41[116]}
   );
   gpc1_1 gpc2092 (
      {stage0_41[230]},
      {stage1_41[117]}
   );
   gpc1_1 gpc2093 (
      {stage0_41[231]},
      {stage1_41[118]}
   );
   gpc1_1 gpc2094 (
      {stage0_41[232]},
      {stage1_41[119]}
   );
   gpc1_1 gpc2095 (
      {stage0_41[233]},
      {stage1_41[120]}
   );
   gpc1_1 gpc2096 (
      {stage0_41[234]},
      {stage1_41[121]}
   );
   gpc1_1 gpc2097 (
      {stage0_41[235]},
      {stage1_41[122]}
   );
   gpc1_1 gpc2098 (
      {stage0_41[236]},
      {stage1_41[123]}
   );
   gpc1_1 gpc2099 (
      {stage0_41[237]},
      {stage1_41[124]}
   );
   gpc1_1 gpc2100 (
      {stage0_41[238]},
      {stage1_41[125]}
   );
   gpc1_1 gpc2101 (
      {stage0_41[239]},
      {stage1_41[126]}
   );
   gpc1_1 gpc2102 (
      {stage0_41[240]},
      {stage1_41[127]}
   );
   gpc1_1 gpc2103 (
      {stage0_41[241]},
      {stage1_41[128]}
   );
   gpc1_1 gpc2104 (
      {stage0_41[242]},
      {stage1_41[129]}
   );
   gpc1_1 gpc2105 (
      {stage0_41[243]},
      {stage1_41[130]}
   );
   gpc1_1 gpc2106 (
      {stage0_41[244]},
      {stage1_41[131]}
   );
   gpc1_1 gpc2107 (
      {stage0_41[245]},
      {stage1_41[132]}
   );
   gpc1_1 gpc2108 (
      {stage0_41[246]},
      {stage1_41[133]}
   );
   gpc1_1 gpc2109 (
      {stage0_41[247]},
      {stage1_41[134]}
   );
   gpc1_1 gpc2110 (
      {stage0_41[248]},
      {stage1_41[135]}
   );
   gpc1_1 gpc2111 (
      {stage0_41[249]},
      {stage1_41[136]}
   );
   gpc1_1 gpc2112 (
      {stage0_41[250]},
      {stage1_41[137]}
   );
   gpc1_1 gpc2113 (
      {stage0_41[251]},
      {stage1_41[138]}
   );
   gpc1_1 gpc2114 (
      {stage0_41[252]},
      {stage1_41[139]}
   );
   gpc1_1 gpc2115 (
      {stage0_41[253]},
      {stage1_41[140]}
   );
   gpc1_1 gpc2116 (
      {stage0_41[254]},
      {stage1_41[141]}
   );
   gpc1_1 gpc2117 (
      {stage0_41[255]},
      {stage1_41[142]}
   );
   gpc1_1 gpc2118 (
      {stage0_42[175]},
      {stage1_42[91]}
   );
   gpc1_1 gpc2119 (
      {stage0_42[176]},
      {stage1_42[92]}
   );
   gpc1_1 gpc2120 (
      {stage0_42[177]},
      {stage1_42[93]}
   );
   gpc1_1 gpc2121 (
      {stage0_42[178]},
      {stage1_42[94]}
   );
   gpc1_1 gpc2122 (
      {stage0_42[179]},
      {stage1_42[95]}
   );
   gpc1_1 gpc2123 (
      {stage0_42[180]},
      {stage1_42[96]}
   );
   gpc1_1 gpc2124 (
      {stage0_42[181]},
      {stage1_42[97]}
   );
   gpc1_1 gpc2125 (
      {stage0_42[182]},
      {stage1_42[98]}
   );
   gpc1_1 gpc2126 (
      {stage0_42[183]},
      {stage1_42[99]}
   );
   gpc1_1 gpc2127 (
      {stage0_42[184]},
      {stage1_42[100]}
   );
   gpc1_1 gpc2128 (
      {stage0_42[185]},
      {stage1_42[101]}
   );
   gpc1_1 gpc2129 (
      {stage0_42[186]},
      {stage1_42[102]}
   );
   gpc1_1 gpc2130 (
      {stage0_42[187]},
      {stage1_42[103]}
   );
   gpc1_1 gpc2131 (
      {stage0_42[188]},
      {stage1_42[104]}
   );
   gpc1_1 gpc2132 (
      {stage0_42[189]},
      {stage1_42[105]}
   );
   gpc1_1 gpc2133 (
      {stage0_42[190]},
      {stage1_42[106]}
   );
   gpc1_1 gpc2134 (
      {stage0_42[191]},
      {stage1_42[107]}
   );
   gpc1_1 gpc2135 (
      {stage0_42[192]},
      {stage1_42[108]}
   );
   gpc1_1 gpc2136 (
      {stage0_42[193]},
      {stage1_42[109]}
   );
   gpc1_1 gpc2137 (
      {stage0_42[194]},
      {stage1_42[110]}
   );
   gpc1_1 gpc2138 (
      {stage0_42[195]},
      {stage1_42[111]}
   );
   gpc1_1 gpc2139 (
      {stage0_42[196]},
      {stage1_42[112]}
   );
   gpc1_1 gpc2140 (
      {stage0_42[197]},
      {stage1_42[113]}
   );
   gpc1_1 gpc2141 (
      {stage0_42[198]},
      {stage1_42[114]}
   );
   gpc1_1 gpc2142 (
      {stage0_42[199]},
      {stage1_42[115]}
   );
   gpc1_1 gpc2143 (
      {stage0_42[200]},
      {stage1_42[116]}
   );
   gpc1_1 gpc2144 (
      {stage0_42[201]},
      {stage1_42[117]}
   );
   gpc1_1 gpc2145 (
      {stage0_42[202]},
      {stage1_42[118]}
   );
   gpc1_1 gpc2146 (
      {stage0_42[203]},
      {stage1_42[119]}
   );
   gpc1_1 gpc2147 (
      {stage0_42[204]},
      {stage1_42[120]}
   );
   gpc1_1 gpc2148 (
      {stage0_42[205]},
      {stage1_42[121]}
   );
   gpc1_1 gpc2149 (
      {stage0_42[206]},
      {stage1_42[122]}
   );
   gpc1_1 gpc2150 (
      {stage0_42[207]},
      {stage1_42[123]}
   );
   gpc1_1 gpc2151 (
      {stage0_42[208]},
      {stage1_42[124]}
   );
   gpc1_1 gpc2152 (
      {stage0_42[209]},
      {stage1_42[125]}
   );
   gpc1_1 gpc2153 (
      {stage0_42[210]},
      {stage1_42[126]}
   );
   gpc1_1 gpc2154 (
      {stage0_42[211]},
      {stage1_42[127]}
   );
   gpc1_1 gpc2155 (
      {stage0_42[212]},
      {stage1_42[128]}
   );
   gpc1_1 gpc2156 (
      {stage0_42[213]},
      {stage1_42[129]}
   );
   gpc1_1 gpc2157 (
      {stage0_42[214]},
      {stage1_42[130]}
   );
   gpc1_1 gpc2158 (
      {stage0_42[215]},
      {stage1_42[131]}
   );
   gpc1_1 gpc2159 (
      {stage0_42[216]},
      {stage1_42[132]}
   );
   gpc1_1 gpc2160 (
      {stage0_42[217]},
      {stage1_42[133]}
   );
   gpc1_1 gpc2161 (
      {stage0_42[218]},
      {stage1_42[134]}
   );
   gpc1_1 gpc2162 (
      {stage0_42[219]},
      {stage1_42[135]}
   );
   gpc1_1 gpc2163 (
      {stage0_42[220]},
      {stage1_42[136]}
   );
   gpc1_1 gpc2164 (
      {stage0_42[221]},
      {stage1_42[137]}
   );
   gpc1_1 gpc2165 (
      {stage0_42[222]},
      {stage1_42[138]}
   );
   gpc1_1 gpc2166 (
      {stage0_42[223]},
      {stage1_42[139]}
   );
   gpc1_1 gpc2167 (
      {stage0_42[224]},
      {stage1_42[140]}
   );
   gpc1_1 gpc2168 (
      {stage0_42[225]},
      {stage1_42[141]}
   );
   gpc1_1 gpc2169 (
      {stage0_42[226]},
      {stage1_42[142]}
   );
   gpc1_1 gpc2170 (
      {stage0_42[227]},
      {stage1_42[143]}
   );
   gpc1_1 gpc2171 (
      {stage0_42[228]},
      {stage1_42[144]}
   );
   gpc1_1 gpc2172 (
      {stage0_42[229]},
      {stage1_42[145]}
   );
   gpc1_1 gpc2173 (
      {stage0_42[230]},
      {stage1_42[146]}
   );
   gpc1_1 gpc2174 (
      {stage0_42[231]},
      {stage1_42[147]}
   );
   gpc1_1 gpc2175 (
      {stage0_42[232]},
      {stage1_42[148]}
   );
   gpc1_1 gpc2176 (
      {stage0_42[233]},
      {stage1_42[149]}
   );
   gpc1_1 gpc2177 (
      {stage0_42[234]},
      {stage1_42[150]}
   );
   gpc1_1 gpc2178 (
      {stage0_42[235]},
      {stage1_42[151]}
   );
   gpc1_1 gpc2179 (
      {stage0_42[236]},
      {stage1_42[152]}
   );
   gpc1_1 gpc2180 (
      {stage0_42[237]},
      {stage1_42[153]}
   );
   gpc1_1 gpc2181 (
      {stage0_42[238]},
      {stage1_42[154]}
   );
   gpc1_1 gpc2182 (
      {stage0_42[239]},
      {stage1_42[155]}
   );
   gpc1_1 gpc2183 (
      {stage0_42[240]},
      {stage1_42[156]}
   );
   gpc1_1 gpc2184 (
      {stage0_42[241]},
      {stage1_42[157]}
   );
   gpc1_1 gpc2185 (
      {stage0_42[242]},
      {stage1_42[158]}
   );
   gpc1_1 gpc2186 (
      {stage0_42[243]},
      {stage1_42[159]}
   );
   gpc1_1 gpc2187 (
      {stage0_42[244]},
      {stage1_42[160]}
   );
   gpc1_1 gpc2188 (
      {stage0_42[245]},
      {stage1_42[161]}
   );
   gpc1_1 gpc2189 (
      {stage0_42[246]},
      {stage1_42[162]}
   );
   gpc1_1 gpc2190 (
      {stage0_42[247]},
      {stage1_42[163]}
   );
   gpc1_1 gpc2191 (
      {stage0_42[248]},
      {stage1_42[164]}
   );
   gpc1_1 gpc2192 (
      {stage0_42[249]},
      {stage1_42[165]}
   );
   gpc1_1 gpc2193 (
      {stage0_42[250]},
      {stage1_42[166]}
   );
   gpc1_1 gpc2194 (
      {stage0_42[251]},
      {stage1_42[167]}
   );
   gpc1_1 gpc2195 (
      {stage0_42[252]},
      {stage1_42[168]}
   );
   gpc1_1 gpc2196 (
      {stage0_42[253]},
      {stage1_42[169]}
   );
   gpc1_1 gpc2197 (
      {stage0_42[254]},
      {stage1_42[170]}
   );
   gpc1_1 gpc2198 (
      {stage0_42[255]},
      {stage1_42[171]}
   );
   gpc1_1 gpc2199 (
      {stage0_43[250]},
      {stage1_43[73]}
   );
   gpc1_1 gpc2200 (
      {stage0_43[251]},
      {stage1_43[74]}
   );
   gpc1_1 gpc2201 (
      {stage0_43[252]},
      {stage1_43[75]}
   );
   gpc1_1 gpc2202 (
      {stage0_43[253]},
      {stage1_43[76]}
   );
   gpc1_1 gpc2203 (
      {stage0_43[254]},
      {stage1_43[77]}
   );
   gpc1_1 gpc2204 (
      {stage0_43[255]},
      {stage1_43[78]}
   );
   gpc1_1 gpc2205 (
      {stage0_44[203]},
      {stage1_44[93]}
   );
   gpc1_1 gpc2206 (
      {stage0_44[204]},
      {stage1_44[94]}
   );
   gpc1_1 gpc2207 (
      {stage0_44[205]},
      {stage1_44[95]}
   );
   gpc1_1 gpc2208 (
      {stage0_44[206]},
      {stage1_44[96]}
   );
   gpc1_1 gpc2209 (
      {stage0_44[207]},
      {stage1_44[97]}
   );
   gpc1_1 gpc2210 (
      {stage0_44[208]},
      {stage1_44[98]}
   );
   gpc1_1 gpc2211 (
      {stage0_44[209]},
      {stage1_44[99]}
   );
   gpc1_1 gpc2212 (
      {stage0_44[210]},
      {stage1_44[100]}
   );
   gpc1_1 gpc2213 (
      {stage0_44[211]},
      {stage1_44[101]}
   );
   gpc1_1 gpc2214 (
      {stage0_44[212]},
      {stage1_44[102]}
   );
   gpc1_1 gpc2215 (
      {stage0_44[213]},
      {stage1_44[103]}
   );
   gpc1_1 gpc2216 (
      {stage0_44[214]},
      {stage1_44[104]}
   );
   gpc1_1 gpc2217 (
      {stage0_44[215]},
      {stage1_44[105]}
   );
   gpc1_1 gpc2218 (
      {stage0_44[216]},
      {stage1_44[106]}
   );
   gpc1_1 gpc2219 (
      {stage0_44[217]},
      {stage1_44[107]}
   );
   gpc1_1 gpc2220 (
      {stage0_44[218]},
      {stage1_44[108]}
   );
   gpc1_1 gpc2221 (
      {stage0_44[219]},
      {stage1_44[109]}
   );
   gpc1_1 gpc2222 (
      {stage0_44[220]},
      {stage1_44[110]}
   );
   gpc1_1 gpc2223 (
      {stage0_44[221]},
      {stage1_44[111]}
   );
   gpc1_1 gpc2224 (
      {stage0_44[222]},
      {stage1_44[112]}
   );
   gpc1_1 gpc2225 (
      {stage0_44[223]},
      {stage1_44[113]}
   );
   gpc1_1 gpc2226 (
      {stage0_44[224]},
      {stage1_44[114]}
   );
   gpc1_1 gpc2227 (
      {stage0_44[225]},
      {stage1_44[115]}
   );
   gpc1_1 gpc2228 (
      {stage0_44[226]},
      {stage1_44[116]}
   );
   gpc1_1 gpc2229 (
      {stage0_44[227]},
      {stage1_44[117]}
   );
   gpc1_1 gpc2230 (
      {stage0_44[228]},
      {stage1_44[118]}
   );
   gpc1_1 gpc2231 (
      {stage0_44[229]},
      {stage1_44[119]}
   );
   gpc1_1 gpc2232 (
      {stage0_44[230]},
      {stage1_44[120]}
   );
   gpc1_1 gpc2233 (
      {stage0_44[231]},
      {stage1_44[121]}
   );
   gpc1_1 gpc2234 (
      {stage0_44[232]},
      {stage1_44[122]}
   );
   gpc1_1 gpc2235 (
      {stage0_44[233]},
      {stage1_44[123]}
   );
   gpc1_1 gpc2236 (
      {stage0_44[234]},
      {stage1_44[124]}
   );
   gpc1_1 gpc2237 (
      {stage0_44[235]},
      {stage1_44[125]}
   );
   gpc1_1 gpc2238 (
      {stage0_44[236]},
      {stage1_44[126]}
   );
   gpc1_1 gpc2239 (
      {stage0_44[237]},
      {stage1_44[127]}
   );
   gpc1_1 gpc2240 (
      {stage0_44[238]},
      {stage1_44[128]}
   );
   gpc1_1 gpc2241 (
      {stage0_44[239]},
      {stage1_44[129]}
   );
   gpc1_1 gpc2242 (
      {stage0_44[240]},
      {stage1_44[130]}
   );
   gpc1_1 gpc2243 (
      {stage0_44[241]},
      {stage1_44[131]}
   );
   gpc1_1 gpc2244 (
      {stage0_44[242]},
      {stage1_44[132]}
   );
   gpc1_1 gpc2245 (
      {stage0_44[243]},
      {stage1_44[133]}
   );
   gpc1_1 gpc2246 (
      {stage0_44[244]},
      {stage1_44[134]}
   );
   gpc1_1 gpc2247 (
      {stage0_44[245]},
      {stage1_44[135]}
   );
   gpc1_1 gpc2248 (
      {stage0_44[246]},
      {stage1_44[136]}
   );
   gpc1_1 gpc2249 (
      {stage0_44[247]},
      {stage1_44[137]}
   );
   gpc1_1 gpc2250 (
      {stage0_44[248]},
      {stage1_44[138]}
   );
   gpc1_1 gpc2251 (
      {stage0_44[249]},
      {stage1_44[139]}
   );
   gpc1_1 gpc2252 (
      {stage0_44[250]},
      {stage1_44[140]}
   );
   gpc1_1 gpc2253 (
      {stage0_44[251]},
      {stage1_44[141]}
   );
   gpc1_1 gpc2254 (
      {stage0_44[252]},
      {stage1_44[142]}
   );
   gpc1_1 gpc2255 (
      {stage0_44[253]},
      {stage1_44[143]}
   );
   gpc1_1 gpc2256 (
      {stage0_44[254]},
      {stage1_44[144]}
   );
   gpc1_1 gpc2257 (
      {stage0_44[255]},
      {stage1_44[145]}
   );
   gpc1_1 gpc2258 (
      {stage0_45[200]},
      {stage1_45[103]}
   );
   gpc1_1 gpc2259 (
      {stage0_45[201]},
      {stage1_45[104]}
   );
   gpc1_1 gpc2260 (
      {stage0_45[202]},
      {stage1_45[105]}
   );
   gpc1_1 gpc2261 (
      {stage0_45[203]},
      {stage1_45[106]}
   );
   gpc1_1 gpc2262 (
      {stage0_45[204]},
      {stage1_45[107]}
   );
   gpc1_1 gpc2263 (
      {stage0_45[205]},
      {stage1_45[108]}
   );
   gpc1_1 gpc2264 (
      {stage0_45[206]},
      {stage1_45[109]}
   );
   gpc1_1 gpc2265 (
      {stage0_45[207]},
      {stage1_45[110]}
   );
   gpc1_1 gpc2266 (
      {stage0_45[208]},
      {stage1_45[111]}
   );
   gpc1_1 gpc2267 (
      {stage0_45[209]},
      {stage1_45[112]}
   );
   gpc1_1 gpc2268 (
      {stage0_45[210]},
      {stage1_45[113]}
   );
   gpc1_1 gpc2269 (
      {stage0_45[211]},
      {stage1_45[114]}
   );
   gpc1_1 gpc2270 (
      {stage0_45[212]},
      {stage1_45[115]}
   );
   gpc1_1 gpc2271 (
      {stage0_45[213]},
      {stage1_45[116]}
   );
   gpc1_1 gpc2272 (
      {stage0_45[214]},
      {stage1_45[117]}
   );
   gpc1_1 gpc2273 (
      {stage0_45[215]},
      {stage1_45[118]}
   );
   gpc1_1 gpc2274 (
      {stage0_45[216]},
      {stage1_45[119]}
   );
   gpc1_1 gpc2275 (
      {stage0_45[217]},
      {stage1_45[120]}
   );
   gpc1_1 gpc2276 (
      {stage0_45[218]},
      {stage1_45[121]}
   );
   gpc1_1 gpc2277 (
      {stage0_45[219]},
      {stage1_45[122]}
   );
   gpc1_1 gpc2278 (
      {stage0_45[220]},
      {stage1_45[123]}
   );
   gpc1_1 gpc2279 (
      {stage0_45[221]},
      {stage1_45[124]}
   );
   gpc1_1 gpc2280 (
      {stage0_45[222]},
      {stage1_45[125]}
   );
   gpc1_1 gpc2281 (
      {stage0_45[223]},
      {stage1_45[126]}
   );
   gpc1_1 gpc2282 (
      {stage0_45[224]},
      {stage1_45[127]}
   );
   gpc1_1 gpc2283 (
      {stage0_45[225]},
      {stage1_45[128]}
   );
   gpc1_1 gpc2284 (
      {stage0_45[226]},
      {stage1_45[129]}
   );
   gpc1_1 gpc2285 (
      {stage0_45[227]},
      {stage1_45[130]}
   );
   gpc1_1 gpc2286 (
      {stage0_45[228]},
      {stage1_45[131]}
   );
   gpc1_1 gpc2287 (
      {stage0_45[229]},
      {stage1_45[132]}
   );
   gpc1_1 gpc2288 (
      {stage0_45[230]},
      {stage1_45[133]}
   );
   gpc1_1 gpc2289 (
      {stage0_45[231]},
      {stage1_45[134]}
   );
   gpc1_1 gpc2290 (
      {stage0_45[232]},
      {stage1_45[135]}
   );
   gpc1_1 gpc2291 (
      {stage0_45[233]},
      {stage1_45[136]}
   );
   gpc1_1 gpc2292 (
      {stage0_45[234]},
      {stage1_45[137]}
   );
   gpc1_1 gpc2293 (
      {stage0_45[235]},
      {stage1_45[138]}
   );
   gpc1_1 gpc2294 (
      {stage0_45[236]},
      {stage1_45[139]}
   );
   gpc1_1 gpc2295 (
      {stage0_45[237]},
      {stage1_45[140]}
   );
   gpc1_1 gpc2296 (
      {stage0_45[238]},
      {stage1_45[141]}
   );
   gpc1_1 gpc2297 (
      {stage0_45[239]},
      {stage1_45[142]}
   );
   gpc1_1 gpc2298 (
      {stage0_45[240]},
      {stage1_45[143]}
   );
   gpc1_1 gpc2299 (
      {stage0_45[241]},
      {stage1_45[144]}
   );
   gpc1_1 gpc2300 (
      {stage0_45[242]},
      {stage1_45[145]}
   );
   gpc1_1 gpc2301 (
      {stage0_45[243]},
      {stage1_45[146]}
   );
   gpc1_1 gpc2302 (
      {stage0_45[244]},
      {stage1_45[147]}
   );
   gpc1_1 gpc2303 (
      {stage0_45[245]},
      {stage1_45[148]}
   );
   gpc1_1 gpc2304 (
      {stage0_45[246]},
      {stage1_45[149]}
   );
   gpc1_1 gpc2305 (
      {stage0_45[247]},
      {stage1_45[150]}
   );
   gpc1_1 gpc2306 (
      {stage0_45[248]},
      {stage1_45[151]}
   );
   gpc1_1 gpc2307 (
      {stage0_45[249]},
      {stage1_45[152]}
   );
   gpc1_1 gpc2308 (
      {stage0_45[250]},
      {stage1_45[153]}
   );
   gpc1_1 gpc2309 (
      {stage0_45[251]},
      {stage1_45[154]}
   );
   gpc1_1 gpc2310 (
      {stage0_45[252]},
      {stage1_45[155]}
   );
   gpc1_1 gpc2311 (
      {stage0_45[253]},
      {stage1_45[156]}
   );
   gpc1_1 gpc2312 (
      {stage0_45[254]},
      {stage1_45[157]}
   );
   gpc1_1 gpc2313 (
      {stage0_45[255]},
      {stage1_45[158]}
   );
   gpc1_1 gpc2314 (
      {stage0_46[237]},
      {stage1_46[82]}
   );
   gpc1_1 gpc2315 (
      {stage0_46[238]},
      {stage1_46[83]}
   );
   gpc1_1 gpc2316 (
      {stage0_46[239]},
      {stage1_46[84]}
   );
   gpc1_1 gpc2317 (
      {stage0_46[240]},
      {stage1_46[85]}
   );
   gpc1_1 gpc2318 (
      {stage0_46[241]},
      {stage1_46[86]}
   );
   gpc1_1 gpc2319 (
      {stage0_46[242]},
      {stage1_46[87]}
   );
   gpc1_1 gpc2320 (
      {stage0_46[243]},
      {stage1_46[88]}
   );
   gpc1_1 gpc2321 (
      {stage0_46[244]},
      {stage1_46[89]}
   );
   gpc1_1 gpc2322 (
      {stage0_46[245]},
      {stage1_46[90]}
   );
   gpc1_1 gpc2323 (
      {stage0_46[246]},
      {stage1_46[91]}
   );
   gpc1_1 gpc2324 (
      {stage0_46[247]},
      {stage1_46[92]}
   );
   gpc1_1 gpc2325 (
      {stage0_46[248]},
      {stage1_46[93]}
   );
   gpc1_1 gpc2326 (
      {stage0_46[249]},
      {stage1_46[94]}
   );
   gpc1_1 gpc2327 (
      {stage0_46[250]},
      {stage1_46[95]}
   );
   gpc1_1 gpc2328 (
      {stage0_46[251]},
      {stage1_46[96]}
   );
   gpc1_1 gpc2329 (
      {stage0_46[252]},
      {stage1_46[97]}
   );
   gpc1_1 gpc2330 (
      {stage0_46[253]},
      {stage1_46[98]}
   );
   gpc1_1 gpc2331 (
      {stage0_46[254]},
      {stage1_46[99]}
   );
   gpc1_1 gpc2332 (
      {stage0_46[255]},
      {stage1_46[100]}
   );
   gpc1_1 gpc2333 (
      {stage0_47[205]},
      {stage1_47[79]}
   );
   gpc1_1 gpc2334 (
      {stage0_47[206]},
      {stage1_47[80]}
   );
   gpc1_1 gpc2335 (
      {stage0_47[207]},
      {stage1_47[81]}
   );
   gpc1_1 gpc2336 (
      {stage0_47[208]},
      {stage1_47[82]}
   );
   gpc1_1 gpc2337 (
      {stage0_47[209]},
      {stage1_47[83]}
   );
   gpc1_1 gpc2338 (
      {stage0_47[210]},
      {stage1_47[84]}
   );
   gpc1_1 gpc2339 (
      {stage0_47[211]},
      {stage1_47[85]}
   );
   gpc1_1 gpc2340 (
      {stage0_47[212]},
      {stage1_47[86]}
   );
   gpc1_1 gpc2341 (
      {stage0_47[213]},
      {stage1_47[87]}
   );
   gpc1_1 gpc2342 (
      {stage0_47[214]},
      {stage1_47[88]}
   );
   gpc1_1 gpc2343 (
      {stage0_47[215]},
      {stage1_47[89]}
   );
   gpc1_1 gpc2344 (
      {stage0_47[216]},
      {stage1_47[90]}
   );
   gpc1_1 gpc2345 (
      {stage0_47[217]},
      {stage1_47[91]}
   );
   gpc1_1 gpc2346 (
      {stage0_47[218]},
      {stage1_47[92]}
   );
   gpc1_1 gpc2347 (
      {stage0_47[219]},
      {stage1_47[93]}
   );
   gpc1_1 gpc2348 (
      {stage0_47[220]},
      {stage1_47[94]}
   );
   gpc1_1 gpc2349 (
      {stage0_47[221]},
      {stage1_47[95]}
   );
   gpc1_1 gpc2350 (
      {stage0_47[222]},
      {stage1_47[96]}
   );
   gpc1_1 gpc2351 (
      {stage0_47[223]},
      {stage1_47[97]}
   );
   gpc1_1 gpc2352 (
      {stage0_47[224]},
      {stage1_47[98]}
   );
   gpc1_1 gpc2353 (
      {stage0_47[225]},
      {stage1_47[99]}
   );
   gpc1_1 gpc2354 (
      {stage0_47[226]},
      {stage1_47[100]}
   );
   gpc1_1 gpc2355 (
      {stage0_47[227]},
      {stage1_47[101]}
   );
   gpc1_1 gpc2356 (
      {stage0_47[228]},
      {stage1_47[102]}
   );
   gpc1_1 gpc2357 (
      {stage0_47[229]},
      {stage1_47[103]}
   );
   gpc1_1 gpc2358 (
      {stage0_47[230]},
      {stage1_47[104]}
   );
   gpc1_1 gpc2359 (
      {stage0_47[231]},
      {stage1_47[105]}
   );
   gpc1_1 gpc2360 (
      {stage0_47[232]},
      {stage1_47[106]}
   );
   gpc1_1 gpc2361 (
      {stage0_47[233]},
      {stage1_47[107]}
   );
   gpc1_1 gpc2362 (
      {stage0_47[234]},
      {stage1_47[108]}
   );
   gpc1_1 gpc2363 (
      {stage0_47[235]},
      {stage1_47[109]}
   );
   gpc1_1 gpc2364 (
      {stage0_47[236]},
      {stage1_47[110]}
   );
   gpc1_1 gpc2365 (
      {stage0_47[237]},
      {stage1_47[111]}
   );
   gpc1_1 gpc2366 (
      {stage0_47[238]},
      {stage1_47[112]}
   );
   gpc1_1 gpc2367 (
      {stage0_47[239]},
      {stage1_47[113]}
   );
   gpc1_1 gpc2368 (
      {stage0_47[240]},
      {stage1_47[114]}
   );
   gpc1_1 gpc2369 (
      {stage0_47[241]},
      {stage1_47[115]}
   );
   gpc1_1 gpc2370 (
      {stage0_47[242]},
      {stage1_47[116]}
   );
   gpc1_1 gpc2371 (
      {stage0_47[243]},
      {stage1_47[117]}
   );
   gpc1_1 gpc2372 (
      {stage0_47[244]},
      {stage1_47[118]}
   );
   gpc1_1 gpc2373 (
      {stage0_47[245]},
      {stage1_47[119]}
   );
   gpc1_1 gpc2374 (
      {stage0_47[246]},
      {stage1_47[120]}
   );
   gpc1_1 gpc2375 (
      {stage0_47[247]},
      {stage1_47[121]}
   );
   gpc1_1 gpc2376 (
      {stage0_47[248]},
      {stage1_47[122]}
   );
   gpc1_1 gpc2377 (
      {stage0_47[249]},
      {stage1_47[123]}
   );
   gpc1_1 gpc2378 (
      {stage0_47[250]},
      {stage1_47[124]}
   );
   gpc1_1 gpc2379 (
      {stage0_47[251]},
      {stage1_47[125]}
   );
   gpc1_1 gpc2380 (
      {stage0_47[252]},
      {stage1_47[126]}
   );
   gpc1_1 gpc2381 (
      {stage0_47[253]},
      {stage1_47[127]}
   );
   gpc1_1 gpc2382 (
      {stage0_47[254]},
      {stage1_47[128]}
   );
   gpc1_1 gpc2383 (
      {stage0_47[255]},
      {stage1_47[129]}
   );
   gpc1_1 gpc2384 (
      {stage0_48[253]},
      {stage1_48[105]}
   );
   gpc1_1 gpc2385 (
      {stage0_48[254]},
      {stage1_48[106]}
   );
   gpc1_1 gpc2386 (
      {stage0_48[255]},
      {stage1_48[107]}
   );
   gpc1_1 gpc2387 (
      {stage0_49[209]},
      {stage1_49[105]}
   );
   gpc1_1 gpc2388 (
      {stage0_49[210]},
      {stage1_49[106]}
   );
   gpc1_1 gpc2389 (
      {stage0_49[211]},
      {stage1_49[107]}
   );
   gpc1_1 gpc2390 (
      {stage0_49[212]},
      {stage1_49[108]}
   );
   gpc1_1 gpc2391 (
      {stage0_49[213]},
      {stage1_49[109]}
   );
   gpc1_1 gpc2392 (
      {stage0_49[214]},
      {stage1_49[110]}
   );
   gpc1_1 gpc2393 (
      {stage0_49[215]},
      {stage1_49[111]}
   );
   gpc1_1 gpc2394 (
      {stage0_49[216]},
      {stage1_49[112]}
   );
   gpc1_1 gpc2395 (
      {stage0_49[217]},
      {stage1_49[113]}
   );
   gpc1_1 gpc2396 (
      {stage0_49[218]},
      {stage1_49[114]}
   );
   gpc1_1 gpc2397 (
      {stage0_49[219]},
      {stage1_49[115]}
   );
   gpc1_1 gpc2398 (
      {stage0_49[220]},
      {stage1_49[116]}
   );
   gpc1_1 gpc2399 (
      {stage0_49[221]},
      {stage1_49[117]}
   );
   gpc1_1 gpc2400 (
      {stage0_49[222]},
      {stage1_49[118]}
   );
   gpc1_1 gpc2401 (
      {stage0_49[223]},
      {stage1_49[119]}
   );
   gpc1_1 gpc2402 (
      {stage0_49[224]},
      {stage1_49[120]}
   );
   gpc1_1 gpc2403 (
      {stage0_49[225]},
      {stage1_49[121]}
   );
   gpc1_1 gpc2404 (
      {stage0_49[226]},
      {stage1_49[122]}
   );
   gpc1_1 gpc2405 (
      {stage0_49[227]},
      {stage1_49[123]}
   );
   gpc1_1 gpc2406 (
      {stage0_49[228]},
      {stage1_49[124]}
   );
   gpc1_1 gpc2407 (
      {stage0_49[229]},
      {stage1_49[125]}
   );
   gpc1_1 gpc2408 (
      {stage0_49[230]},
      {stage1_49[126]}
   );
   gpc1_1 gpc2409 (
      {stage0_49[231]},
      {stage1_49[127]}
   );
   gpc1_1 gpc2410 (
      {stage0_49[232]},
      {stage1_49[128]}
   );
   gpc1_1 gpc2411 (
      {stage0_49[233]},
      {stage1_49[129]}
   );
   gpc1_1 gpc2412 (
      {stage0_49[234]},
      {stage1_49[130]}
   );
   gpc1_1 gpc2413 (
      {stage0_49[235]},
      {stage1_49[131]}
   );
   gpc1_1 gpc2414 (
      {stage0_49[236]},
      {stage1_49[132]}
   );
   gpc1_1 gpc2415 (
      {stage0_49[237]},
      {stage1_49[133]}
   );
   gpc1_1 gpc2416 (
      {stage0_49[238]},
      {stage1_49[134]}
   );
   gpc1_1 gpc2417 (
      {stage0_49[239]},
      {stage1_49[135]}
   );
   gpc1_1 gpc2418 (
      {stage0_49[240]},
      {stage1_49[136]}
   );
   gpc1_1 gpc2419 (
      {stage0_49[241]},
      {stage1_49[137]}
   );
   gpc1_1 gpc2420 (
      {stage0_49[242]},
      {stage1_49[138]}
   );
   gpc1_1 gpc2421 (
      {stage0_49[243]},
      {stage1_49[139]}
   );
   gpc1_1 gpc2422 (
      {stage0_49[244]},
      {stage1_49[140]}
   );
   gpc1_1 gpc2423 (
      {stage0_49[245]},
      {stage1_49[141]}
   );
   gpc1_1 gpc2424 (
      {stage0_49[246]},
      {stage1_49[142]}
   );
   gpc1_1 gpc2425 (
      {stage0_49[247]},
      {stage1_49[143]}
   );
   gpc1_1 gpc2426 (
      {stage0_49[248]},
      {stage1_49[144]}
   );
   gpc1_1 gpc2427 (
      {stage0_49[249]},
      {stage1_49[145]}
   );
   gpc1_1 gpc2428 (
      {stage0_49[250]},
      {stage1_49[146]}
   );
   gpc1_1 gpc2429 (
      {stage0_49[251]},
      {stage1_49[147]}
   );
   gpc1_1 gpc2430 (
      {stage0_49[252]},
      {stage1_49[148]}
   );
   gpc1_1 gpc2431 (
      {stage0_49[253]},
      {stage1_49[149]}
   );
   gpc1_1 gpc2432 (
      {stage0_49[254]},
      {stage1_49[150]}
   );
   gpc1_1 gpc2433 (
      {stage0_49[255]},
      {stage1_49[151]}
   );
   gpc1_1 gpc2434 (
      {stage0_50[243]},
      {stage1_50[86]}
   );
   gpc1_1 gpc2435 (
      {stage0_50[244]},
      {stage1_50[87]}
   );
   gpc1_1 gpc2436 (
      {stage0_50[245]},
      {stage1_50[88]}
   );
   gpc1_1 gpc2437 (
      {stage0_50[246]},
      {stage1_50[89]}
   );
   gpc1_1 gpc2438 (
      {stage0_50[247]},
      {stage1_50[90]}
   );
   gpc1_1 gpc2439 (
      {stage0_50[248]},
      {stage1_50[91]}
   );
   gpc1_1 gpc2440 (
      {stage0_50[249]},
      {stage1_50[92]}
   );
   gpc1_1 gpc2441 (
      {stage0_50[250]},
      {stage1_50[93]}
   );
   gpc1_1 gpc2442 (
      {stage0_50[251]},
      {stage1_50[94]}
   );
   gpc1_1 gpc2443 (
      {stage0_50[252]},
      {stage1_50[95]}
   );
   gpc1_1 gpc2444 (
      {stage0_50[253]},
      {stage1_50[96]}
   );
   gpc1_1 gpc2445 (
      {stage0_50[254]},
      {stage1_50[97]}
   );
   gpc1_1 gpc2446 (
      {stage0_50[255]},
      {stage1_50[98]}
   );
   gpc1_1 gpc2447 (
      {stage0_51[236]},
      {stage1_51[86]}
   );
   gpc1_1 gpc2448 (
      {stage0_51[237]},
      {stage1_51[87]}
   );
   gpc1_1 gpc2449 (
      {stage0_51[238]},
      {stage1_51[88]}
   );
   gpc1_1 gpc2450 (
      {stage0_51[239]},
      {stage1_51[89]}
   );
   gpc1_1 gpc2451 (
      {stage0_51[240]},
      {stage1_51[90]}
   );
   gpc1_1 gpc2452 (
      {stage0_51[241]},
      {stage1_51[91]}
   );
   gpc1_1 gpc2453 (
      {stage0_51[242]},
      {stage1_51[92]}
   );
   gpc1_1 gpc2454 (
      {stage0_51[243]},
      {stage1_51[93]}
   );
   gpc1_1 gpc2455 (
      {stage0_51[244]},
      {stage1_51[94]}
   );
   gpc1_1 gpc2456 (
      {stage0_51[245]},
      {stage1_51[95]}
   );
   gpc1_1 gpc2457 (
      {stage0_51[246]},
      {stage1_51[96]}
   );
   gpc1_1 gpc2458 (
      {stage0_51[247]},
      {stage1_51[97]}
   );
   gpc1_1 gpc2459 (
      {stage0_51[248]},
      {stage1_51[98]}
   );
   gpc1_1 gpc2460 (
      {stage0_51[249]},
      {stage1_51[99]}
   );
   gpc1_1 gpc2461 (
      {stage0_51[250]},
      {stage1_51[100]}
   );
   gpc1_1 gpc2462 (
      {stage0_51[251]},
      {stage1_51[101]}
   );
   gpc1_1 gpc2463 (
      {stage0_51[252]},
      {stage1_51[102]}
   );
   gpc1_1 gpc2464 (
      {stage0_51[253]},
      {stage1_51[103]}
   );
   gpc1_1 gpc2465 (
      {stage0_51[254]},
      {stage1_51[104]}
   );
   gpc1_1 gpc2466 (
      {stage0_51[255]},
      {stage1_51[105]}
   );
   gpc1_1 gpc2467 (
      {stage0_52[223]},
      {stage1_52[107]}
   );
   gpc1_1 gpc2468 (
      {stage0_52[224]},
      {stage1_52[108]}
   );
   gpc1_1 gpc2469 (
      {stage0_52[225]},
      {stage1_52[109]}
   );
   gpc1_1 gpc2470 (
      {stage0_52[226]},
      {stage1_52[110]}
   );
   gpc1_1 gpc2471 (
      {stage0_52[227]},
      {stage1_52[111]}
   );
   gpc1_1 gpc2472 (
      {stage0_52[228]},
      {stage1_52[112]}
   );
   gpc1_1 gpc2473 (
      {stage0_52[229]},
      {stage1_52[113]}
   );
   gpc1_1 gpc2474 (
      {stage0_52[230]},
      {stage1_52[114]}
   );
   gpc1_1 gpc2475 (
      {stage0_52[231]},
      {stage1_52[115]}
   );
   gpc1_1 gpc2476 (
      {stage0_52[232]},
      {stage1_52[116]}
   );
   gpc1_1 gpc2477 (
      {stage0_52[233]},
      {stage1_52[117]}
   );
   gpc1_1 gpc2478 (
      {stage0_52[234]},
      {stage1_52[118]}
   );
   gpc1_1 gpc2479 (
      {stage0_52[235]},
      {stage1_52[119]}
   );
   gpc1_1 gpc2480 (
      {stage0_52[236]},
      {stage1_52[120]}
   );
   gpc1_1 gpc2481 (
      {stage0_52[237]},
      {stage1_52[121]}
   );
   gpc1_1 gpc2482 (
      {stage0_52[238]},
      {stage1_52[122]}
   );
   gpc1_1 gpc2483 (
      {stage0_52[239]},
      {stage1_52[123]}
   );
   gpc1_1 gpc2484 (
      {stage0_52[240]},
      {stage1_52[124]}
   );
   gpc1_1 gpc2485 (
      {stage0_52[241]},
      {stage1_52[125]}
   );
   gpc1_1 gpc2486 (
      {stage0_52[242]},
      {stage1_52[126]}
   );
   gpc1_1 gpc2487 (
      {stage0_52[243]},
      {stage1_52[127]}
   );
   gpc1_1 gpc2488 (
      {stage0_52[244]},
      {stage1_52[128]}
   );
   gpc1_1 gpc2489 (
      {stage0_52[245]},
      {stage1_52[129]}
   );
   gpc1_1 gpc2490 (
      {stage0_52[246]},
      {stage1_52[130]}
   );
   gpc1_1 gpc2491 (
      {stage0_52[247]},
      {stage1_52[131]}
   );
   gpc1_1 gpc2492 (
      {stage0_52[248]},
      {stage1_52[132]}
   );
   gpc1_1 gpc2493 (
      {stage0_52[249]},
      {stage1_52[133]}
   );
   gpc1_1 gpc2494 (
      {stage0_52[250]},
      {stage1_52[134]}
   );
   gpc1_1 gpc2495 (
      {stage0_52[251]},
      {stage1_52[135]}
   );
   gpc1_1 gpc2496 (
      {stage0_52[252]},
      {stage1_52[136]}
   );
   gpc1_1 gpc2497 (
      {stage0_52[253]},
      {stage1_52[137]}
   );
   gpc1_1 gpc2498 (
      {stage0_52[254]},
      {stage1_52[138]}
   );
   gpc1_1 gpc2499 (
      {stage0_52[255]},
      {stage1_52[139]}
   );
   gpc1_1 gpc2500 (
      {stage0_53[254]},
      {stage1_53[106]}
   );
   gpc1_1 gpc2501 (
      {stage0_53[255]},
      {stage1_53[107]}
   );
   gpc1_1 gpc2502 (
      {stage0_54[178]},
      {stage1_54[82]}
   );
   gpc1_1 gpc2503 (
      {stage0_54[179]},
      {stage1_54[83]}
   );
   gpc1_1 gpc2504 (
      {stage0_54[180]},
      {stage1_54[84]}
   );
   gpc1_1 gpc2505 (
      {stage0_54[181]},
      {stage1_54[85]}
   );
   gpc1_1 gpc2506 (
      {stage0_54[182]},
      {stage1_54[86]}
   );
   gpc1_1 gpc2507 (
      {stage0_54[183]},
      {stage1_54[87]}
   );
   gpc1_1 gpc2508 (
      {stage0_54[184]},
      {stage1_54[88]}
   );
   gpc1_1 gpc2509 (
      {stage0_54[185]},
      {stage1_54[89]}
   );
   gpc1_1 gpc2510 (
      {stage0_54[186]},
      {stage1_54[90]}
   );
   gpc1_1 gpc2511 (
      {stage0_54[187]},
      {stage1_54[91]}
   );
   gpc1_1 gpc2512 (
      {stage0_54[188]},
      {stage1_54[92]}
   );
   gpc1_1 gpc2513 (
      {stage0_54[189]},
      {stage1_54[93]}
   );
   gpc1_1 gpc2514 (
      {stage0_54[190]},
      {stage1_54[94]}
   );
   gpc1_1 gpc2515 (
      {stage0_54[191]},
      {stage1_54[95]}
   );
   gpc1_1 gpc2516 (
      {stage0_54[192]},
      {stage1_54[96]}
   );
   gpc1_1 gpc2517 (
      {stage0_54[193]},
      {stage1_54[97]}
   );
   gpc1_1 gpc2518 (
      {stage0_54[194]},
      {stage1_54[98]}
   );
   gpc1_1 gpc2519 (
      {stage0_54[195]},
      {stage1_54[99]}
   );
   gpc1_1 gpc2520 (
      {stage0_54[196]},
      {stage1_54[100]}
   );
   gpc1_1 gpc2521 (
      {stage0_54[197]},
      {stage1_54[101]}
   );
   gpc1_1 gpc2522 (
      {stage0_54[198]},
      {stage1_54[102]}
   );
   gpc1_1 gpc2523 (
      {stage0_54[199]},
      {stage1_54[103]}
   );
   gpc1_1 gpc2524 (
      {stage0_54[200]},
      {stage1_54[104]}
   );
   gpc1_1 gpc2525 (
      {stage0_54[201]},
      {stage1_54[105]}
   );
   gpc1_1 gpc2526 (
      {stage0_54[202]},
      {stage1_54[106]}
   );
   gpc1_1 gpc2527 (
      {stage0_54[203]},
      {stage1_54[107]}
   );
   gpc1_1 gpc2528 (
      {stage0_54[204]},
      {stage1_54[108]}
   );
   gpc1_1 gpc2529 (
      {stage0_54[205]},
      {stage1_54[109]}
   );
   gpc1_1 gpc2530 (
      {stage0_54[206]},
      {stage1_54[110]}
   );
   gpc1_1 gpc2531 (
      {stage0_54[207]},
      {stage1_54[111]}
   );
   gpc1_1 gpc2532 (
      {stage0_54[208]},
      {stage1_54[112]}
   );
   gpc1_1 gpc2533 (
      {stage0_54[209]},
      {stage1_54[113]}
   );
   gpc1_1 gpc2534 (
      {stage0_54[210]},
      {stage1_54[114]}
   );
   gpc1_1 gpc2535 (
      {stage0_54[211]},
      {stage1_54[115]}
   );
   gpc1_1 gpc2536 (
      {stage0_54[212]},
      {stage1_54[116]}
   );
   gpc1_1 gpc2537 (
      {stage0_54[213]},
      {stage1_54[117]}
   );
   gpc1_1 gpc2538 (
      {stage0_54[214]},
      {stage1_54[118]}
   );
   gpc1_1 gpc2539 (
      {stage0_54[215]},
      {stage1_54[119]}
   );
   gpc1_1 gpc2540 (
      {stage0_54[216]},
      {stage1_54[120]}
   );
   gpc1_1 gpc2541 (
      {stage0_54[217]},
      {stage1_54[121]}
   );
   gpc1_1 gpc2542 (
      {stage0_54[218]},
      {stage1_54[122]}
   );
   gpc1_1 gpc2543 (
      {stage0_54[219]},
      {stage1_54[123]}
   );
   gpc1_1 gpc2544 (
      {stage0_54[220]},
      {stage1_54[124]}
   );
   gpc1_1 gpc2545 (
      {stage0_54[221]},
      {stage1_54[125]}
   );
   gpc1_1 gpc2546 (
      {stage0_54[222]},
      {stage1_54[126]}
   );
   gpc1_1 gpc2547 (
      {stage0_54[223]},
      {stage1_54[127]}
   );
   gpc1_1 gpc2548 (
      {stage0_54[224]},
      {stage1_54[128]}
   );
   gpc1_1 gpc2549 (
      {stage0_54[225]},
      {stage1_54[129]}
   );
   gpc1_1 gpc2550 (
      {stage0_54[226]},
      {stage1_54[130]}
   );
   gpc1_1 gpc2551 (
      {stage0_54[227]},
      {stage1_54[131]}
   );
   gpc1_1 gpc2552 (
      {stage0_54[228]},
      {stage1_54[132]}
   );
   gpc1_1 gpc2553 (
      {stage0_54[229]},
      {stage1_54[133]}
   );
   gpc1_1 gpc2554 (
      {stage0_54[230]},
      {stage1_54[134]}
   );
   gpc1_1 gpc2555 (
      {stage0_54[231]},
      {stage1_54[135]}
   );
   gpc1_1 gpc2556 (
      {stage0_54[232]},
      {stage1_54[136]}
   );
   gpc1_1 gpc2557 (
      {stage0_54[233]},
      {stage1_54[137]}
   );
   gpc1_1 gpc2558 (
      {stage0_54[234]},
      {stage1_54[138]}
   );
   gpc1_1 gpc2559 (
      {stage0_54[235]},
      {stage1_54[139]}
   );
   gpc1_1 gpc2560 (
      {stage0_54[236]},
      {stage1_54[140]}
   );
   gpc1_1 gpc2561 (
      {stage0_54[237]},
      {stage1_54[141]}
   );
   gpc1_1 gpc2562 (
      {stage0_54[238]},
      {stage1_54[142]}
   );
   gpc1_1 gpc2563 (
      {stage0_54[239]},
      {stage1_54[143]}
   );
   gpc1_1 gpc2564 (
      {stage0_54[240]},
      {stage1_54[144]}
   );
   gpc1_1 gpc2565 (
      {stage0_54[241]},
      {stage1_54[145]}
   );
   gpc1_1 gpc2566 (
      {stage0_54[242]},
      {stage1_54[146]}
   );
   gpc1_1 gpc2567 (
      {stage0_54[243]},
      {stage1_54[147]}
   );
   gpc1_1 gpc2568 (
      {stage0_54[244]},
      {stage1_54[148]}
   );
   gpc1_1 gpc2569 (
      {stage0_54[245]},
      {stage1_54[149]}
   );
   gpc1_1 gpc2570 (
      {stage0_54[246]},
      {stage1_54[150]}
   );
   gpc1_1 gpc2571 (
      {stage0_54[247]},
      {stage1_54[151]}
   );
   gpc1_1 gpc2572 (
      {stage0_54[248]},
      {stage1_54[152]}
   );
   gpc1_1 gpc2573 (
      {stage0_54[249]},
      {stage1_54[153]}
   );
   gpc1_1 gpc2574 (
      {stage0_54[250]},
      {stage1_54[154]}
   );
   gpc1_1 gpc2575 (
      {stage0_54[251]},
      {stage1_54[155]}
   );
   gpc1_1 gpc2576 (
      {stage0_54[252]},
      {stage1_54[156]}
   );
   gpc1_1 gpc2577 (
      {stage0_54[253]},
      {stage1_54[157]}
   );
   gpc1_1 gpc2578 (
      {stage0_54[254]},
      {stage1_54[158]}
   );
   gpc1_1 gpc2579 (
      {stage0_54[255]},
      {stage1_54[159]}
   );
   gpc1_1 gpc2580 (
      {stage0_55[250]},
      {stage1_55[84]}
   );
   gpc1_1 gpc2581 (
      {stage0_55[251]},
      {stage1_55[85]}
   );
   gpc1_1 gpc2582 (
      {stage0_55[252]},
      {stage1_55[86]}
   );
   gpc1_1 gpc2583 (
      {stage0_55[253]},
      {stage1_55[87]}
   );
   gpc1_1 gpc2584 (
      {stage0_55[254]},
      {stage1_55[88]}
   );
   gpc1_1 gpc2585 (
      {stage0_55[255]},
      {stage1_55[89]}
   );
   gpc1_1 gpc2586 (
      {stage0_56[176]},
      {stage1_56[98]}
   );
   gpc1_1 gpc2587 (
      {stage0_56[177]},
      {stage1_56[99]}
   );
   gpc1_1 gpc2588 (
      {stage0_56[178]},
      {stage1_56[100]}
   );
   gpc1_1 gpc2589 (
      {stage0_56[179]},
      {stage1_56[101]}
   );
   gpc1_1 gpc2590 (
      {stage0_56[180]},
      {stage1_56[102]}
   );
   gpc1_1 gpc2591 (
      {stage0_56[181]},
      {stage1_56[103]}
   );
   gpc1_1 gpc2592 (
      {stage0_56[182]},
      {stage1_56[104]}
   );
   gpc1_1 gpc2593 (
      {stage0_56[183]},
      {stage1_56[105]}
   );
   gpc1_1 gpc2594 (
      {stage0_56[184]},
      {stage1_56[106]}
   );
   gpc1_1 gpc2595 (
      {stage0_56[185]},
      {stage1_56[107]}
   );
   gpc1_1 gpc2596 (
      {stage0_56[186]},
      {stage1_56[108]}
   );
   gpc1_1 gpc2597 (
      {stage0_56[187]},
      {stage1_56[109]}
   );
   gpc1_1 gpc2598 (
      {stage0_56[188]},
      {stage1_56[110]}
   );
   gpc1_1 gpc2599 (
      {stage0_56[189]},
      {stage1_56[111]}
   );
   gpc1_1 gpc2600 (
      {stage0_56[190]},
      {stage1_56[112]}
   );
   gpc1_1 gpc2601 (
      {stage0_56[191]},
      {stage1_56[113]}
   );
   gpc1_1 gpc2602 (
      {stage0_56[192]},
      {stage1_56[114]}
   );
   gpc1_1 gpc2603 (
      {stage0_56[193]},
      {stage1_56[115]}
   );
   gpc1_1 gpc2604 (
      {stage0_56[194]},
      {stage1_56[116]}
   );
   gpc1_1 gpc2605 (
      {stage0_56[195]},
      {stage1_56[117]}
   );
   gpc1_1 gpc2606 (
      {stage0_56[196]},
      {stage1_56[118]}
   );
   gpc1_1 gpc2607 (
      {stage0_56[197]},
      {stage1_56[119]}
   );
   gpc1_1 gpc2608 (
      {stage0_56[198]},
      {stage1_56[120]}
   );
   gpc1_1 gpc2609 (
      {stage0_56[199]},
      {stage1_56[121]}
   );
   gpc1_1 gpc2610 (
      {stage0_56[200]},
      {stage1_56[122]}
   );
   gpc1_1 gpc2611 (
      {stage0_56[201]},
      {stage1_56[123]}
   );
   gpc1_1 gpc2612 (
      {stage0_56[202]},
      {stage1_56[124]}
   );
   gpc1_1 gpc2613 (
      {stage0_56[203]},
      {stage1_56[125]}
   );
   gpc1_1 gpc2614 (
      {stage0_56[204]},
      {stage1_56[126]}
   );
   gpc1_1 gpc2615 (
      {stage0_56[205]},
      {stage1_56[127]}
   );
   gpc1_1 gpc2616 (
      {stage0_56[206]},
      {stage1_56[128]}
   );
   gpc1_1 gpc2617 (
      {stage0_56[207]},
      {stage1_56[129]}
   );
   gpc1_1 gpc2618 (
      {stage0_56[208]},
      {stage1_56[130]}
   );
   gpc1_1 gpc2619 (
      {stage0_56[209]},
      {stage1_56[131]}
   );
   gpc1_1 gpc2620 (
      {stage0_56[210]},
      {stage1_56[132]}
   );
   gpc1_1 gpc2621 (
      {stage0_56[211]},
      {stage1_56[133]}
   );
   gpc1_1 gpc2622 (
      {stage0_56[212]},
      {stage1_56[134]}
   );
   gpc1_1 gpc2623 (
      {stage0_56[213]},
      {stage1_56[135]}
   );
   gpc1_1 gpc2624 (
      {stage0_56[214]},
      {stage1_56[136]}
   );
   gpc1_1 gpc2625 (
      {stage0_56[215]},
      {stage1_56[137]}
   );
   gpc1_1 gpc2626 (
      {stage0_56[216]},
      {stage1_56[138]}
   );
   gpc1_1 gpc2627 (
      {stage0_56[217]},
      {stage1_56[139]}
   );
   gpc1_1 gpc2628 (
      {stage0_56[218]},
      {stage1_56[140]}
   );
   gpc1_1 gpc2629 (
      {stage0_56[219]},
      {stage1_56[141]}
   );
   gpc1_1 gpc2630 (
      {stage0_56[220]},
      {stage1_56[142]}
   );
   gpc1_1 gpc2631 (
      {stage0_56[221]},
      {stage1_56[143]}
   );
   gpc1_1 gpc2632 (
      {stage0_56[222]},
      {stage1_56[144]}
   );
   gpc1_1 gpc2633 (
      {stage0_56[223]},
      {stage1_56[145]}
   );
   gpc1_1 gpc2634 (
      {stage0_56[224]},
      {stage1_56[146]}
   );
   gpc1_1 gpc2635 (
      {stage0_56[225]},
      {stage1_56[147]}
   );
   gpc1_1 gpc2636 (
      {stage0_56[226]},
      {stage1_56[148]}
   );
   gpc1_1 gpc2637 (
      {stage0_56[227]},
      {stage1_56[149]}
   );
   gpc1_1 gpc2638 (
      {stage0_56[228]},
      {stage1_56[150]}
   );
   gpc1_1 gpc2639 (
      {stage0_56[229]},
      {stage1_56[151]}
   );
   gpc1_1 gpc2640 (
      {stage0_56[230]},
      {stage1_56[152]}
   );
   gpc1_1 gpc2641 (
      {stage0_56[231]},
      {stage1_56[153]}
   );
   gpc1_1 gpc2642 (
      {stage0_56[232]},
      {stage1_56[154]}
   );
   gpc1_1 gpc2643 (
      {stage0_56[233]},
      {stage1_56[155]}
   );
   gpc1_1 gpc2644 (
      {stage0_56[234]},
      {stage1_56[156]}
   );
   gpc1_1 gpc2645 (
      {stage0_56[235]},
      {stage1_56[157]}
   );
   gpc1_1 gpc2646 (
      {stage0_56[236]},
      {stage1_56[158]}
   );
   gpc1_1 gpc2647 (
      {stage0_56[237]},
      {stage1_56[159]}
   );
   gpc1_1 gpc2648 (
      {stage0_56[238]},
      {stage1_56[160]}
   );
   gpc1_1 gpc2649 (
      {stage0_56[239]},
      {stage1_56[161]}
   );
   gpc1_1 gpc2650 (
      {stage0_56[240]},
      {stage1_56[162]}
   );
   gpc1_1 gpc2651 (
      {stage0_56[241]},
      {stage1_56[163]}
   );
   gpc1_1 gpc2652 (
      {stage0_56[242]},
      {stage1_56[164]}
   );
   gpc1_1 gpc2653 (
      {stage0_56[243]},
      {stage1_56[165]}
   );
   gpc1_1 gpc2654 (
      {stage0_56[244]},
      {stage1_56[166]}
   );
   gpc1_1 gpc2655 (
      {stage0_56[245]},
      {stage1_56[167]}
   );
   gpc1_1 gpc2656 (
      {stage0_56[246]},
      {stage1_56[168]}
   );
   gpc1_1 gpc2657 (
      {stage0_56[247]},
      {stage1_56[169]}
   );
   gpc1_1 gpc2658 (
      {stage0_56[248]},
      {stage1_56[170]}
   );
   gpc1_1 gpc2659 (
      {stage0_56[249]},
      {stage1_56[171]}
   );
   gpc1_1 gpc2660 (
      {stage0_56[250]},
      {stage1_56[172]}
   );
   gpc1_1 gpc2661 (
      {stage0_56[251]},
      {stage1_56[173]}
   );
   gpc1_1 gpc2662 (
      {stage0_56[252]},
      {stage1_56[174]}
   );
   gpc1_1 gpc2663 (
      {stage0_56[253]},
      {stage1_56[175]}
   );
   gpc1_1 gpc2664 (
      {stage0_56[254]},
      {stage1_56[176]}
   );
   gpc1_1 gpc2665 (
      {stage0_56[255]},
      {stage1_56[177]}
   );
   gpc1_1 gpc2666 (
      {stage0_57[253]},
      {stage1_57[102]}
   );
   gpc1_1 gpc2667 (
      {stage0_57[254]},
      {stage1_57[103]}
   );
   gpc1_1 gpc2668 (
      {stage0_57[255]},
      {stage1_57[104]}
   );
   gpc1_1 gpc2669 (
      {stage0_58[255]},
      {stage1_58[85]}
   );
   gpc1_1 gpc2670 (
      {stage0_59[194]},
      {stage1_59[86]}
   );
   gpc1_1 gpc2671 (
      {stage0_59[195]},
      {stage1_59[87]}
   );
   gpc1_1 gpc2672 (
      {stage0_59[196]},
      {stage1_59[88]}
   );
   gpc1_1 gpc2673 (
      {stage0_59[197]},
      {stage1_59[89]}
   );
   gpc1_1 gpc2674 (
      {stage0_59[198]},
      {stage1_59[90]}
   );
   gpc1_1 gpc2675 (
      {stage0_59[199]},
      {stage1_59[91]}
   );
   gpc1_1 gpc2676 (
      {stage0_59[200]},
      {stage1_59[92]}
   );
   gpc1_1 gpc2677 (
      {stage0_59[201]},
      {stage1_59[93]}
   );
   gpc1_1 gpc2678 (
      {stage0_59[202]},
      {stage1_59[94]}
   );
   gpc1_1 gpc2679 (
      {stage0_59[203]},
      {stage1_59[95]}
   );
   gpc1_1 gpc2680 (
      {stage0_59[204]},
      {stage1_59[96]}
   );
   gpc1_1 gpc2681 (
      {stage0_59[205]},
      {stage1_59[97]}
   );
   gpc1_1 gpc2682 (
      {stage0_59[206]},
      {stage1_59[98]}
   );
   gpc1_1 gpc2683 (
      {stage0_59[207]},
      {stage1_59[99]}
   );
   gpc1_1 gpc2684 (
      {stage0_59[208]},
      {stage1_59[100]}
   );
   gpc1_1 gpc2685 (
      {stage0_59[209]},
      {stage1_59[101]}
   );
   gpc1_1 gpc2686 (
      {stage0_59[210]},
      {stage1_59[102]}
   );
   gpc1_1 gpc2687 (
      {stage0_59[211]},
      {stage1_59[103]}
   );
   gpc1_1 gpc2688 (
      {stage0_59[212]},
      {stage1_59[104]}
   );
   gpc1_1 gpc2689 (
      {stage0_59[213]},
      {stage1_59[105]}
   );
   gpc1_1 gpc2690 (
      {stage0_59[214]},
      {stage1_59[106]}
   );
   gpc1_1 gpc2691 (
      {stage0_59[215]},
      {stage1_59[107]}
   );
   gpc1_1 gpc2692 (
      {stage0_59[216]},
      {stage1_59[108]}
   );
   gpc1_1 gpc2693 (
      {stage0_59[217]},
      {stage1_59[109]}
   );
   gpc1_1 gpc2694 (
      {stage0_59[218]},
      {stage1_59[110]}
   );
   gpc1_1 gpc2695 (
      {stage0_59[219]},
      {stage1_59[111]}
   );
   gpc1_1 gpc2696 (
      {stage0_59[220]},
      {stage1_59[112]}
   );
   gpc1_1 gpc2697 (
      {stage0_59[221]},
      {stage1_59[113]}
   );
   gpc1_1 gpc2698 (
      {stage0_59[222]},
      {stage1_59[114]}
   );
   gpc1_1 gpc2699 (
      {stage0_59[223]},
      {stage1_59[115]}
   );
   gpc1_1 gpc2700 (
      {stage0_59[224]},
      {stage1_59[116]}
   );
   gpc1_1 gpc2701 (
      {stage0_59[225]},
      {stage1_59[117]}
   );
   gpc1_1 gpc2702 (
      {stage0_59[226]},
      {stage1_59[118]}
   );
   gpc1_1 gpc2703 (
      {stage0_59[227]},
      {stage1_59[119]}
   );
   gpc1_1 gpc2704 (
      {stage0_59[228]},
      {stage1_59[120]}
   );
   gpc1_1 gpc2705 (
      {stage0_59[229]},
      {stage1_59[121]}
   );
   gpc1_1 gpc2706 (
      {stage0_59[230]},
      {stage1_59[122]}
   );
   gpc1_1 gpc2707 (
      {stage0_59[231]},
      {stage1_59[123]}
   );
   gpc1_1 gpc2708 (
      {stage0_59[232]},
      {stage1_59[124]}
   );
   gpc1_1 gpc2709 (
      {stage0_59[233]},
      {stage1_59[125]}
   );
   gpc1_1 gpc2710 (
      {stage0_59[234]},
      {stage1_59[126]}
   );
   gpc1_1 gpc2711 (
      {stage0_59[235]},
      {stage1_59[127]}
   );
   gpc1_1 gpc2712 (
      {stage0_59[236]},
      {stage1_59[128]}
   );
   gpc1_1 gpc2713 (
      {stage0_59[237]},
      {stage1_59[129]}
   );
   gpc1_1 gpc2714 (
      {stage0_59[238]},
      {stage1_59[130]}
   );
   gpc1_1 gpc2715 (
      {stage0_59[239]},
      {stage1_59[131]}
   );
   gpc1_1 gpc2716 (
      {stage0_59[240]},
      {stage1_59[132]}
   );
   gpc1_1 gpc2717 (
      {stage0_59[241]},
      {stage1_59[133]}
   );
   gpc1_1 gpc2718 (
      {stage0_59[242]},
      {stage1_59[134]}
   );
   gpc1_1 gpc2719 (
      {stage0_59[243]},
      {stage1_59[135]}
   );
   gpc1_1 gpc2720 (
      {stage0_59[244]},
      {stage1_59[136]}
   );
   gpc1_1 gpc2721 (
      {stage0_59[245]},
      {stage1_59[137]}
   );
   gpc1_1 gpc2722 (
      {stage0_59[246]},
      {stage1_59[138]}
   );
   gpc1_1 gpc2723 (
      {stage0_59[247]},
      {stage1_59[139]}
   );
   gpc1_1 gpc2724 (
      {stage0_59[248]},
      {stage1_59[140]}
   );
   gpc1_1 gpc2725 (
      {stage0_59[249]},
      {stage1_59[141]}
   );
   gpc1_1 gpc2726 (
      {stage0_59[250]},
      {stage1_59[142]}
   );
   gpc1_1 gpc2727 (
      {stage0_59[251]},
      {stage1_59[143]}
   );
   gpc1_1 gpc2728 (
      {stage0_59[252]},
      {stage1_59[144]}
   );
   gpc1_1 gpc2729 (
      {stage0_59[253]},
      {stage1_59[145]}
   );
   gpc1_1 gpc2730 (
      {stage0_59[254]},
      {stage1_59[146]}
   );
   gpc1_1 gpc2731 (
      {stage0_59[255]},
      {stage1_59[147]}
   );
   gpc1_1 gpc2732 (
      {stage0_60[210]},
      {stage1_60[96]}
   );
   gpc1_1 gpc2733 (
      {stage0_60[211]},
      {stage1_60[97]}
   );
   gpc1_1 gpc2734 (
      {stage0_60[212]},
      {stage1_60[98]}
   );
   gpc1_1 gpc2735 (
      {stage0_60[213]},
      {stage1_60[99]}
   );
   gpc1_1 gpc2736 (
      {stage0_60[214]},
      {stage1_60[100]}
   );
   gpc1_1 gpc2737 (
      {stage0_60[215]},
      {stage1_60[101]}
   );
   gpc1_1 gpc2738 (
      {stage0_60[216]},
      {stage1_60[102]}
   );
   gpc1_1 gpc2739 (
      {stage0_60[217]},
      {stage1_60[103]}
   );
   gpc1_1 gpc2740 (
      {stage0_60[218]},
      {stage1_60[104]}
   );
   gpc1_1 gpc2741 (
      {stage0_60[219]},
      {stage1_60[105]}
   );
   gpc1_1 gpc2742 (
      {stage0_60[220]},
      {stage1_60[106]}
   );
   gpc1_1 gpc2743 (
      {stage0_60[221]},
      {stage1_60[107]}
   );
   gpc1_1 gpc2744 (
      {stage0_60[222]},
      {stage1_60[108]}
   );
   gpc1_1 gpc2745 (
      {stage0_60[223]},
      {stage1_60[109]}
   );
   gpc1_1 gpc2746 (
      {stage0_60[224]},
      {stage1_60[110]}
   );
   gpc1_1 gpc2747 (
      {stage0_60[225]},
      {stage1_60[111]}
   );
   gpc1_1 gpc2748 (
      {stage0_60[226]},
      {stage1_60[112]}
   );
   gpc1_1 gpc2749 (
      {stage0_60[227]},
      {stage1_60[113]}
   );
   gpc1_1 gpc2750 (
      {stage0_60[228]},
      {stage1_60[114]}
   );
   gpc1_1 gpc2751 (
      {stage0_60[229]},
      {stage1_60[115]}
   );
   gpc1_1 gpc2752 (
      {stage0_60[230]},
      {stage1_60[116]}
   );
   gpc1_1 gpc2753 (
      {stage0_60[231]},
      {stage1_60[117]}
   );
   gpc1_1 gpc2754 (
      {stage0_60[232]},
      {stage1_60[118]}
   );
   gpc1_1 gpc2755 (
      {stage0_60[233]},
      {stage1_60[119]}
   );
   gpc1_1 gpc2756 (
      {stage0_60[234]},
      {stage1_60[120]}
   );
   gpc1_1 gpc2757 (
      {stage0_60[235]},
      {stage1_60[121]}
   );
   gpc1_1 gpc2758 (
      {stage0_60[236]},
      {stage1_60[122]}
   );
   gpc1_1 gpc2759 (
      {stage0_60[237]},
      {stage1_60[123]}
   );
   gpc1_1 gpc2760 (
      {stage0_60[238]},
      {stage1_60[124]}
   );
   gpc1_1 gpc2761 (
      {stage0_60[239]},
      {stage1_60[125]}
   );
   gpc1_1 gpc2762 (
      {stage0_60[240]},
      {stage1_60[126]}
   );
   gpc1_1 gpc2763 (
      {stage0_60[241]},
      {stage1_60[127]}
   );
   gpc1_1 gpc2764 (
      {stage0_60[242]},
      {stage1_60[128]}
   );
   gpc1_1 gpc2765 (
      {stage0_60[243]},
      {stage1_60[129]}
   );
   gpc1_1 gpc2766 (
      {stage0_60[244]},
      {stage1_60[130]}
   );
   gpc1_1 gpc2767 (
      {stage0_60[245]},
      {stage1_60[131]}
   );
   gpc1_1 gpc2768 (
      {stage0_60[246]},
      {stage1_60[132]}
   );
   gpc1_1 gpc2769 (
      {stage0_60[247]},
      {stage1_60[133]}
   );
   gpc1_1 gpc2770 (
      {stage0_60[248]},
      {stage1_60[134]}
   );
   gpc1_1 gpc2771 (
      {stage0_60[249]},
      {stage1_60[135]}
   );
   gpc1_1 gpc2772 (
      {stage0_60[250]},
      {stage1_60[136]}
   );
   gpc1_1 gpc2773 (
      {stage0_60[251]},
      {stage1_60[137]}
   );
   gpc1_1 gpc2774 (
      {stage0_60[252]},
      {stage1_60[138]}
   );
   gpc1_1 gpc2775 (
      {stage0_60[253]},
      {stage1_60[139]}
   );
   gpc1_1 gpc2776 (
      {stage0_60[254]},
      {stage1_60[140]}
   );
   gpc1_1 gpc2777 (
      {stage0_60[255]},
      {stage1_60[141]}
   );
   gpc1_1 gpc2778 (
      {stage0_62[133]},
      {stage1_62[78]}
   );
   gpc1_1 gpc2779 (
      {stage0_62[134]},
      {stage1_62[79]}
   );
   gpc1_1 gpc2780 (
      {stage0_62[135]},
      {stage1_62[80]}
   );
   gpc1_1 gpc2781 (
      {stage0_62[136]},
      {stage1_62[81]}
   );
   gpc1_1 gpc2782 (
      {stage0_62[137]},
      {stage1_62[82]}
   );
   gpc1_1 gpc2783 (
      {stage0_62[138]},
      {stage1_62[83]}
   );
   gpc1_1 gpc2784 (
      {stage0_62[139]},
      {stage1_62[84]}
   );
   gpc1_1 gpc2785 (
      {stage0_62[140]},
      {stage1_62[85]}
   );
   gpc1_1 gpc2786 (
      {stage0_62[141]},
      {stage1_62[86]}
   );
   gpc1_1 gpc2787 (
      {stage0_62[142]},
      {stage1_62[87]}
   );
   gpc1_1 gpc2788 (
      {stage0_62[143]},
      {stage1_62[88]}
   );
   gpc1_1 gpc2789 (
      {stage0_62[144]},
      {stage1_62[89]}
   );
   gpc1_1 gpc2790 (
      {stage0_62[145]},
      {stage1_62[90]}
   );
   gpc1_1 gpc2791 (
      {stage0_62[146]},
      {stage1_62[91]}
   );
   gpc1_1 gpc2792 (
      {stage0_62[147]},
      {stage1_62[92]}
   );
   gpc1_1 gpc2793 (
      {stage0_62[148]},
      {stage1_62[93]}
   );
   gpc1_1 gpc2794 (
      {stage0_62[149]},
      {stage1_62[94]}
   );
   gpc1_1 gpc2795 (
      {stage0_62[150]},
      {stage1_62[95]}
   );
   gpc1_1 gpc2796 (
      {stage0_62[151]},
      {stage1_62[96]}
   );
   gpc1_1 gpc2797 (
      {stage0_62[152]},
      {stage1_62[97]}
   );
   gpc1_1 gpc2798 (
      {stage0_62[153]},
      {stage1_62[98]}
   );
   gpc1_1 gpc2799 (
      {stage0_62[154]},
      {stage1_62[99]}
   );
   gpc1_1 gpc2800 (
      {stage0_62[155]},
      {stage1_62[100]}
   );
   gpc1_1 gpc2801 (
      {stage0_62[156]},
      {stage1_62[101]}
   );
   gpc1_1 gpc2802 (
      {stage0_62[157]},
      {stage1_62[102]}
   );
   gpc1_1 gpc2803 (
      {stage0_62[158]},
      {stage1_62[103]}
   );
   gpc1_1 gpc2804 (
      {stage0_62[159]},
      {stage1_62[104]}
   );
   gpc1_1 gpc2805 (
      {stage0_62[160]},
      {stage1_62[105]}
   );
   gpc1_1 gpc2806 (
      {stage0_62[161]},
      {stage1_62[106]}
   );
   gpc1_1 gpc2807 (
      {stage0_62[162]},
      {stage1_62[107]}
   );
   gpc1_1 gpc2808 (
      {stage0_62[163]},
      {stage1_62[108]}
   );
   gpc1_1 gpc2809 (
      {stage0_62[164]},
      {stage1_62[109]}
   );
   gpc1_1 gpc2810 (
      {stage0_62[165]},
      {stage1_62[110]}
   );
   gpc1_1 gpc2811 (
      {stage0_62[166]},
      {stage1_62[111]}
   );
   gpc1_1 gpc2812 (
      {stage0_62[167]},
      {stage1_62[112]}
   );
   gpc1_1 gpc2813 (
      {stage0_62[168]},
      {stage1_62[113]}
   );
   gpc1_1 gpc2814 (
      {stage0_62[169]},
      {stage1_62[114]}
   );
   gpc1_1 gpc2815 (
      {stage0_62[170]},
      {stage1_62[115]}
   );
   gpc1_1 gpc2816 (
      {stage0_62[171]},
      {stage1_62[116]}
   );
   gpc1_1 gpc2817 (
      {stage0_62[172]},
      {stage1_62[117]}
   );
   gpc1_1 gpc2818 (
      {stage0_62[173]},
      {stage1_62[118]}
   );
   gpc1_1 gpc2819 (
      {stage0_62[174]},
      {stage1_62[119]}
   );
   gpc1_1 gpc2820 (
      {stage0_62[175]},
      {stage1_62[120]}
   );
   gpc1_1 gpc2821 (
      {stage0_62[176]},
      {stage1_62[121]}
   );
   gpc1_1 gpc2822 (
      {stage0_62[177]},
      {stage1_62[122]}
   );
   gpc1_1 gpc2823 (
      {stage0_62[178]},
      {stage1_62[123]}
   );
   gpc1_1 gpc2824 (
      {stage0_62[179]},
      {stage1_62[124]}
   );
   gpc1_1 gpc2825 (
      {stage0_62[180]},
      {stage1_62[125]}
   );
   gpc1_1 gpc2826 (
      {stage0_62[181]},
      {stage1_62[126]}
   );
   gpc1_1 gpc2827 (
      {stage0_62[182]},
      {stage1_62[127]}
   );
   gpc1_1 gpc2828 (
      {stage0_62[183]},
      {stage1_62[128]}
   );
   gpc1_1 gpc2829 (
      {stage0_62[184]},
      {stage1_62[129]}
   );
   gpc1_1 gpc2830 (
      {stage0_62[185]},
      {stage1_62[130]}
   );
   gpc1_1 gpc2831 (
      {stage0_62[186]},
      {stage1_62[131]}
   );
   gpc1_1 gpc2832 (
      {stage0_62[187]},
      {stage1_62[132]}
   );
   gpc1_1 gpc2833 (
      {stage0_62[188]},
      {stage1_62[133]}
   );
   gpc1_1 gpc2834 (
      {stage0_62[189]},
      {stage1_62[134]}
   );
   gpc1_1 gpc2835 (
      {stage0_62[190]},
      {stage1_62[135]}
   );
   gpc1_1 gpc2836 (
      {stage0_62[191]},
      {stage1_62[136]}
   );
   gpc1_1 gpc2837 (
      {stage0_62[192]},
      {stage1_62[137]}
   );
   gpc1_1 gpc2838 (
      {stage0_62[193]},
      {stage1_62[138]}
   );
   gpc1_1 gpc2839 (
      {stage0_62[194]},
      {stage1_62[139]}
   );
   gpc1_1 gpc2840 (
      {stage0_62[195]},
      {stage1_62[140]}
   );
   gpc1_1 gpc2841 (
      {stage0_62[196]},
      {stage1_62[141]}
   );
   gpc1_1 gpc2842 (
      {stage0_62[197]},
      {stage1_62[142]}
   );
   gpc1_1 gpc2843 (
      {stage0_62[198]},
      {stage1_62[143]}
   );
   gpc1_1 gpc2844 (
      {stage0_62[199]},
      {stage1_62[144]}
   );
   gpc1_1 gpc2845 (
      {stage0_62[200]},
      {stage1_62[145]}
   );
   gpc1_1 gpc2846 (
      {stage0_62[201]},
      {stage1_62[146]}
   );
   gpc1_1 gpc2847 (
      {stage0_62[202]},
      {stage1_62[147]}
   );
   gpc1_1 gpc2848 (
      {stage0_62[203]},
      {stage1_62[148]}
   );
   gpc1_1 gpc2849 (
      {stage0_62[204]},
      {stage1_62[149]}
   );
   gpc1_1 gpc2850 (
      {stage0_62[205]},
      {stage1_62[150]}
   );
   gpc1_1 gpc2851 (
      {stage0_62[206]},
      {stage1_62[151]}
   );
   gpc1_1 gpc2852 (
      {stage0_62[207]},
      {stage1_62[152]}
   );
   gpc1_1 gpc2853 (
      {stage0_62[208]},
      {stage1_62[153]}
   );
   gpc1_1 gpc2854 (
      {stage0_62[209]},
      {stage1_62[154]}
   );
   gpc1_1 gpc2855 (
      {stage0_62[210]},
      {stage1_62[155]}
   );
   gpc1_1 gpc2856 (
      {stage0_62[211]},
      {stage1_62[156]}
   );
   gpc1_1 gpc2857 (
      {stage0_62[212]},
      {stage1_62[157]}
   );
   gpc1_1 gpc2858 (
      {stage0_62[213]},
      {stage1_62[158]}
   );
   gpc1_1 gpc2859 (
      {stage0_62[214]},
      {stage1_62[159]}
   );
   gpc1_1 gpc2860 (
      {stage0_62[215]},
      {stage1_62[160]}
   );
   gpc1_1 gpc2861 (
      {stage0_62[216]},
      {stage1_62[161]}
   );
   gpc1_1 gpc2862 (
      {stage0_62[217]},
      {stage1_62[162]}
   );
   gpc1_1 gpc2863 (
      {stage0_62[218]},
      {stage1_62[163]}
   );
   gpc1_1 gpc2864 (
      {stage0_62[219]},
      {stage1_62[164]}
   );
   gpc1_1 gpc2865 (
      {stage0_62[220]},
      {stage1_62[165]}
   );
   gpc1_1 gpc2866 (
      {stage0_62[221]},
      {stage1_62[166]}
   );
   gpc1_1 gpc2867 (
      {stage0_62[222]},
      {stage1_62[167]}
   );
   gpc1_1 gpc2868 (
      {stage0_62[223]},
      {stage1_62[168]}
   );
   gpc1_1 gpc2869 (
      {stage0_62[224]},
      {stage1_62[169]}
   );
   gpc1_1 gpc2870 (
      {stage0_62[225]},
      {stage1_62[170]}
   );
   gpc1_1 gpc2871 (
      {stage0_62[226]},
      {stage1_62[171]}
   );
   gpc1_1 gpc2872 (
      {stage0_62[227]},
      {stage1_62[172]}
   );
   gpc1_1 gpc2873 (
      {stage0_62[228]},
      {stage1_62[173]}
   );
   gpc1_1 gpc2874 (
      {stage0_62[229]},
      {stage1_62[174]}
   );
   gpc1_1 gpc2875 (
      {stage0_62[230]},
      {stage1_62[175]}
   );
   gpc1_1 gpc2876 (
      {stage0_62[231]},
      {stage1_62[176]}
   );
   gpc1_1 gpc2877 (
      {stage0_62[232]},
      {stage1_62[177]}
   );
   gpc1_1 gpc2878 (
      {stage0_62[233]},
      {stage1_62[178]}
   );
   gpc1_1 gpc2879 (
      {stage0_62[234]},
      {stage1_62[179]}
   );
   gpc1_1 gpc2880 (
      {stage0_62[235]},
      {stage1_62[180]}
   );
   gpc1_1 gpc2881 (
      {stage0_62[236]},
      {stage1_62[181]}
   );
   gpc1_1 gpc2882 (
      {stage0_62[237]},
      {stage1_62[182]}
   );
   gpc1_1 gpc2883 (
      {stage0_62[238]},
      {stage1_62[183]}
   );
   gpc1_1 gpc2884 (
      {stage0_62[239]},
      {stage1_62[184]}
   );
   gpc1_1 gpc2885 (
      {stage0_62[240]},
      {stage1_62[185]}
   );
   gpc1_1 gpc2886 (
      {stage0_62[241]},
      {stage1_62[186]}
   );
   gpc1_1 gpc2887 (
      {stage0_62[242]},
      {stage1_62[187]}
   );
   gpc1_1 gpc2888 (
      {stage0_62[243]},
      {stage1_62[188]}
   );
   gpc1_1 gpc2889 (
      {stage0_62[244]},
      {stage1_62[189]}
   );
   gpc1_1 gpc2890 (
      {stage0_62[245]},
      {stage1_62[190]}
   );
   gpc1_1 gpc2891 (
      {stage0_62[246]},
      {stage1_62[191]}
   );
   gpc1_1 gpc2892 (
      {stage0_62[247]},
      {stage1_62[192]}
   );
   gpc1_1 gpc2893 (
      {stage0_62[248]},
      {stage1_62[193]}
   );
   gpc1_1 gpc2894 (
      {stage0_62[249]},
      {stage1_62[194]}
   );
   gpc1_1 gpc2895 (
      {stage0_62[250]},
      {stage1_62[195]}
   );
   gpc1_1 gpc2896 (
      {stage0_62[251]},
      {stage1_62[196]}
   );
   gpc1_1 gpc2897 (
      {stage0_62[252]},
      {stage1_62[197]}
   );
   gpc1_1 gpc2898 (
      {stage0_62[253]},
      {stage1_62[198]}
   );
   gpc1_1 gpc2899 (
      {stage0_62[254]},
      {stage1_62[199]}
   );
   gpc1_1 gpc2900 (
      {stage0_62[255]},
      {stage1_62[200]}
   );
   gpc1_1 gpc2901 (
      {stage0_63[252]},
      {stage1_63[65]}
   );
   gpc1_1 gpc2902 (
      {stage0_63[253]},
      {stage1_63[66]}
   );
   gpc1_1 gpc2903 (
      {stage0_63[254]},
      {stage1_63[67]}
   );
   gpc1_1 gpc2904 (
      {stage0_63[255]},
      {stage1_63[68]}
   );
   gpc2135_5 gpc2905 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4]},
      {stage1_1[0], stage1_1[1], stage1_1[2]},
      {stage1_2[0]},
      {stage1_3[0], stage1_3[1]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc2135_5 gpc2906 (
      {stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9]},
      {stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[1]},
      {stage1_3[2], stage1_3[3]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc2135_5 gpc2907 (
      {stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_2[2]},
      {stage1_3[4], stage1_3[5]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc2908 (
      {stage1_0[15], stage1_0[16], stage1_0[17], stage1_0[18], stage1_0[19]},
      {stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[3]},
      {stage1_3[6], stage1_3[7]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc606_5 gpc2909 (
      {stage1_0[20], stage1_0[21], stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25]},
      {stage1_2[4], stage1_2[5], stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc2910 (
      {stage1_0[26], stage1_0[27], stage1_0[28], stage1_0[29], stage1_0[30], stage1_0[31]},
      {stage1_2[10], stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc606_5 gpc2911 (
      {stage1_0[32], stage1_0[33], stage1_0[34], stage1_0[35], stage1_0[36], stage1_0[37]},
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc606_5 gpc2912 (
      {stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41], stage1_0[42], stage1_0[43]},
      {stage1_2[22], stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc606_5 gpc2913 (
      {stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47], stage1_0[48], stage1_0[49]},
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc606_5 gpc2914 (
      {stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53], stage1_0[54], stage1_0[55]},
      {stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc606_5 gpc2915 (
      {stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59], stage1_0[60], stage1_0[61]},
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc606_5 gpc2916 (
      {stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65], stage1_0[66], stage1_0[67]},
      {stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc2917 (
      {stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71], stage1_0[72], stage1_0[73]},
      {stage1_2[52], stage1_2[53], stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc2918 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13]},
      {stage2_5[0],stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13]}
   );
   gpc606_5 gpc2919 (
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18], stage1_3[19]},
      {stage2_5[1],stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14]}
   );
   gpc606_5 gpc2920 (
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25]},
      {stage2_5[2],stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15]}
   );
   gpc606_5 gpc2921 (
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31]},
      {stage2_5[3],stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16]}
   );
   gpc606_5 gpc2922 (
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37]},
      {stage2_5[4],stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17]}
   );
   gpc606_5 gpc2923 (
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43]},
      {stage2_5[5],stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18]}
   );
   gpc606_5 gpc2924 (
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49]},
      {stage2_5[6],stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19]}
   );
   gpc615_5 gpc2925 (
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58]},
      {stage1_2[58]},
      {stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage2_5[7],stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20]}
   );
   gpc615_5 gpc2926 (
      {stage1_1[59], stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63]},
      {stage1_2[59]},
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60], stage1_3[61]},
      {stage2_5[8],stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21]}
   );
   gpc615_5 gpc2927 (
      {stage1_1[64], stage1_1[65], stage1_1[66], stage1_1[67], stage1_1[68]},
      {stage1_2[60]},
      {stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65], stage1_3[66], stage1_3[67]},
      {stage2_5[9],stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22]}
   );
   gpc615_5 gpc2928 (
      {stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage1_3[68]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[10],stage2_4[23],stage2_3[23],stage2_2[23]}
   );
   gpc615_5 gpc2929 (
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70]},
      {stage1_3[69]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[11],stage2_4[24],stage2_3[24],stage2_2[24]}
   );
   gpc615_5 gpc2930 (
      {stage1_2[71], stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75]},
      {stage1_3[70]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[12],stage2_4[25],stage2_3[25],stage2_2[25]}
   );
   gpc615_5 gpc2931 (
      {stage1_2[76], stage1_2[77], stage1_2[78], stage1_2[79], stage1_2[80]},
      {stage1_3[71]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[13],stage2_4[26],stage2_3[26],stage2_2[26]}
   );
   gpc615_5 gpc2932 (
      {stage1_2[81], stage1_2[82], stage1_2[83], stage1_2[84], stage1_2[85]},
      {stage1_3[72]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[14],stage2_4[27],stage2_3[27],stage2_2[27]}
   );
   gpc615_5 gpc2933 (
      {stage1_2[86], stage1_2[87], stage1_2[88], stage1_2[89], stage1_2[90]},
      {stage1_3[73]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[15],stage2_4[28],stage2_3[28],stage2_2[28]}
   );
   gpc615_5 gpc2934 (
      {stage1_2[91], stage1_2[92], stage1_2[93], stage1_2[94], stage1_2[95]},
      {stage1_3[74]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[16],stage2_4[29],stage2_3[29],stage2_2[29]}
   );
   gpc615_5 gpc2935 (
      {stage1_2[96], stage1_2[97], stage1_2[98], stage1_2[99], stage1_2[100]},
      {stage1_3[75]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[17],stage2_4[30],stage2_3[30],stage2_2[30]}
   );
   gpc615_5 gpc2936 (
      {stage1_2[101], stage1_2[102], stage1_2[103], stage1_2[104], stage1_2[105]},
      {stage1_3[76]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[18],stage2_4[31],stage2_3[31],stage2_2[31]}
   );
   gpc615_5 gpc2937 (
      {stage1_2[106], stage1_2[107], stage1_2[108], stage1_2[109], stage1_2[110]},
      {stage1_3[77]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[19],stage2_4[32],stage2_3[32],stage2_2[32]}
   );
   gpc615_5 gpc2938 (
      {stage1_2[111], stage1_2[112], stage1_2[113], stage1_2[114], stage1_2[115]},
      {stage1_3[78]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[20],stage2_4[33],stage2_3[33],stage2_2[33]}
   );
   gpc615_5 gpc2939 (
      {stage1_2[116], stage1_2[117], stage1_2[118], stage1_2[119], stage1_2[120]},
      {stage1_3[79]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[21],stage2_4[34],stage2_3[34],stage2_2[34]}
   );
   gpc615_5 gpc2940 (
      {stage1_2[121], stage1_2[122], stage1_2[123], stage1_2[124], stage1_2[125]},
      {stage1_3[80]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[22],stage2_4[35],stage2_3[35],stage2_2[35]}
   );
   gpc615_5 gpc2941 (
      {stage1_2[126], stage1_2[127], stage1_2[128], stage1_2[129], stage1_2[130]},
      {stage1_3[81]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[23],stage2_4[36],stage2_3[36],stage2_2[36]}
   );
   gpc615_5 gpc2942 (
      {stage1_3[82], stage1_3[83], stage1_3[84], stage1_3[85], stage1_3[86]},
      {stage1_4[84]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[14],stage2_5[24],stage2_4[37],stage2_3[37]}
   );
   gpc615_5 gpc2943 (
      {stage1_3[87], stage1_3[88], stage1_3[89], stage1_3[90], stage1_3[91]},
      {stage1_4[85]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[15],stage2_5[25],stage2_4[38],stage2_3[38]}
   );
   gpc606_5 gpc2944 (
      {stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89], stage1_4[90], stage1_4[91]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[2],stage2_6[16],stage2_5[26],stage2_4[39]}
   );
   gpc606_5 gpc2945 (
      {stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95], stage1_4[96], stage1_4[97]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[3],stage2_6[17],stage2_5[27],stage2_4[40]}
   );
   gpc606_5 gpc2946 (
      {stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101], stage1_4[102], stage1_4[103]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[4],stage2_6[18],stage2_5[28],stage2_4[41]}
   );
   gpc606_5 gpc2947 (
      {stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107], stage1_4[108], stage1_4[109]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[5],stage2_6[19],stage2_5[29],stage2_4[42]}
   );
   gpc606_5 gpc2948 (
      {stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113], stage1_4[114], stage1_4[115]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[6],stage2_6[20],stage2_5[30],stage2_4[43]}
   );
   gpc606_5 gpc2949 (
      {stage1_4[116], stage1_4[117], stage1_4[118], stage1_4[119], stage1_4[120], stage1_4[121]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[7],stage2_6[21],stage2_5[31],stage2_4[44]}
   );
   gpc606_5 gpc2950 (
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[6],stage2_7[8],stage2_6[22],stage2_5[32]}
   );
   gpc606_5 gpc2951 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[7],stage2_7[9],stage2_6[23],stage2_5[33]}
   );
   gpc606_5 gpc2952 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[8],stage2_7[10],stage2_6[24],stage2_5[34]}
   );
   gpc606_5 gpc2953 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[9],stage2_7[11],stage2_6[25],stage2_5[35]}
   );
   gpc606_5 gpc2954 (
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[10],stage2_7[12],stage2_6[26],stage2_5[36]}
   );
   gpc606_5 gpc2955 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[11],stage2_7[13],stage2_6[27],stage2_5[37]}
   );
   gpc606_5 gpc2956 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[12],stage2_7[14],stage2_6[28],stage2_5[38]}
   );
   gpc606_5 gpc2957 (
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[13],stage2_7[15],stage2_6[29],stage2_5[39]}
   );
   gpc606_5 gpc2958 (
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[14],stage2_7[16],stage2_6[30],stage2_5[40]}
   );
   gpc606_5 gpc2959 (
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[15],stage2_7[17],stage2_6[31],stage2_5[41]}
   );
   gpc606_5 gpc2960 (
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[16],stage2_7[18],stage2_6[32],stage2_5[42]}
   );
   gpc606_5 gpc2961 (
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[17],stage2_7[19],stage2_6[33],stage2_5[43]}
   );
   gpc606_5 gpc2962 (
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[18],stage2_7[20],stage2_6[34],stage2_5[44]}
   );
   gpc606_5 gpc2963 (
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[19],stage2_7[21],stage2_6[35],stage2_5[45]}
   );
   gpc615_5 gpc2964 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40]},
      {stage1_7[84]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[14],stage2_8[20],stage2_7[22],stage2_6[36]}
   );
   gpc615_5 gpc2965 (
      {stage1_6[41], stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45]},
      {stage1_7[85]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[15],stage2_8[21],stage2_7[23],stage2_6[37]}
   );
   gpc615_5 gpc2966 (
      {stage1_6[46], stage1_6[47], stage1_6[48], stage1_6[49], stage1_6[50]},
      {stage1_7[86]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[16],stage2_8[22],stage2_7[24],stage2_6[38]}
   );
   gpc615_5 gpc2967 (
      {stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54], stage1_6[55]},
      {stage1_7[87]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[17],stage2_8[23],stage2_7[25],stage2_6[39]}
   );
   gpc615_5 gpc2968 (
      {stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59], stage1_6[60]},
      {stage1_7[88]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[18],stage2_8[24],stage2_7[26],stage2_6[40]}
   );
   gpc615_5 gpc2969 (
      {stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage1_7[89]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[19],stage2_8[25],stage2_7[27],stage2_6[41]}
   );
   gpc615_5 gpc2970 (
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70]},
      {stage1_7[90]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[20],stage2_8[26],stage2_7[28],stage2_6[42]}
   );
   gpc615_5 gpc2971 (
      {stage1_6[71], stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75]},
      {stage1_7[91]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[21],stage2_8[27],stage2_7[29],stage2_6[43]}
   );
   gpc615_5 gpc2972 (
      {stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79], stage1_6[80]},
      {stage1_7[92]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[22],stage2_8[28],stage2_7[30],stage2_6[44]}
   );
   gpc615_5 gpc2973 (
      {stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84], stage1_6[85]},
      {stage1_7[93]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[23],stage2_8[29],stage2_7[31],stage2_6[45]}
   );
   gpc615_5 gpc2974 (
      {stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89], stage1_6[90]},
      {stage1_7[94]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[24],stage2_8[30],stage2_7[32],stage2_6[46]}
   );
   gpc615_5 gpc2975 (
      {stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_7[95]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[25],stage2_8[31],stage2_7[33],stage2_6[47]}
   );
   gpc615_5 gpc2976 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100]},
      {stage1_7[96]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[26],stage2_8[32],stage2_7[34],stage2_6[48]}
   );
   gpc615_5 gpc2977 (
      {stage1_6[101], stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105]},
      {stage1_7[97]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[27],stage2_8[33],stage2_7[35],stage2_6[49]}
   );
   gpc615_5 gpc2978 (
      {stage1_6[106], stage1_6[107], stage1_6[108], stage1_6[109], stage1_6[110]},
      {stage1_7[98]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[28],stage2_8[34],stage2_7[36],stage2_6[50]}
   );
   gpc615_5 gpc2979 (
      {stage1_6[111], stage1_6[112], stage1_6[113], stage1_6[114], stage1_6[115]},
      {stage1_7[99]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[29],stage2_8[35],stage2_7[37],stage2_6[51]}
   );
   gpc606_5 gpc2980 (
      {stage1_7[100], stage1_7[101], stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[16],stage2_9[30],stage2_8[36],stage2_7[38]}
   );
   gpc606_5 gpc2981 (
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[17],stage2_9[31],stage2_8[37]}
   );
   gpc606_5 gpc2982 (
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[2],stage2_10[18],stage2_9[32],stage2_8[38]}
   );
   gpc606_5 gpc2983 (
      {stage1_8[108], stage1_8[109], stage1_8[110], stage1_8[111], stage1_8[112], stage1_8[113]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[3],stage2_10[19],stage2_9[33],stage2_8[39]}
   );
   gpc606_5 gpc2984 (
      {stage1_8[114], stage1_8[115], stage1_8[116], stage1_8[117], stage1_8[118], stage1_8[119]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[4],stage2_10[20],stage2_9[34],stage2_8[40]}
   );
   gpc606_5 gpc2985 (
      {stage1_8[120], stage1_8[121], stage1_8[122], stage1_8[123], stage1_8[124], stage1_8[125]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[5],stage2_10[21],stage2_9[35],stage2_8[41]}
   );
   gpc606_5 gpc2986 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[6],stage2_10[22],stage2_9[36],stage2_8[42]}
   );
   gpc615_5 gpc2987 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10]},
      {stage1_10[36]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[6],stage2_11[7],stage2_10[23],stage2_9[37]}
   );
   gpc615_5 gpc2988 (
      {stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15]},
      {stage1_10[37]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[7],stage2_11[8],stage2_10[24],stage2_9[38]}
   );
   gpc615_5 gpc2989 (
      {stage1_9[16], stage1_9[17], stage1_9[18], stage1_9[19], stage1_9[20]},
      {stage1_10[38]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[8],stage2_11[9],stage2_10[25],stage2_9[39]}
   );
   gpc615_5 gpc2990 (
      {stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24], stage1_9[25]},
      {stage1_10[39]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[9],stage2_11[10],stage2_10[26],stage2_9[40]}
   );
   gpc615_5 gpc2991 (
      {stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30]},
      {stage1_10[40]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[10],stage2_11[11],stage2_10[27],stage2_9[41]}
   );
   gpc615_5 gpc2992 (
      {stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_10[41]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[11],stage2_11[12],stage2_10[28],stage2_9[42]}
   );
   gpc615_5 gpc2993 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40]},
      {stage1_10[42]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[12],stage2_11[13],stage2_10[29],stage2_9[43]}
   );
   gpc615_5 gpc2994 (
      {stage1_9[41], stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45]},
      {stage1_10[43]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[13],stage2_11[14],stage2_10[30],stage2_9[44]}
   );
   gpc615_5 gpc2995 (
      {stage1_9[46], stage1_9[47], stage1_9[48], stage1_9[49], stage1_9[50]},
      {stage1_10[44]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[14],stage2_11[15],stage2_10[31],stage2_9[45]}
   );
   gpc615_5 gpc2996 (
      {stage1_9[51], stage1_9[52], stage1_9[53], stage1_9[54], stage1_9[55]},
      {stage1_10[45]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[15],stage2_11[16],stage2_10[32],stage2_9[46]}
   );
   gpc615_5 gpc2997 (
      {stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59], stage1_9[60]},
      {stage1_10[46]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[16],stage2_11[17],stage2_10[33],stage2_9[47]}
   );
   gpc615_5 gpc2998 (
      {stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage1_10[47]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[17],stage2_11[18],stage2_10[34],stage2_9[48]}
   );
   gpc615_5 gpc2999 (
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70]},
      {stage1_10[48]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[18],stage2_11[19],stage2_10[35],stage2_9[49]}
   );
   gpc615_5 gpc3000 (
      {stage1_9[71], stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75]},
      {stage1_10[49]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[19],stage2_11[20],stage2_10[36],stage2_9[50]}
   );
   gpc615_5 gpc3001 (
      {stage1_9[76], stage1_9[77], stage1_9[78], stage1_9[79], stage1_9[80]},
      {stage1_10[50]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[20],stage2_11[21],stage2_10[37],stage2_9[51]}
   );
   gpc615_5 gpc3002 (
      {stage1_9[81], stage1_9[82], stage1_9[83], stage1_9[84], stage1_9[85]},
      {stage1_10[51]},
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94], stage1_11[95]},
      {stage2_13[15],stage2_12[21],stage2_11[22],stage2_10[38],stage2_9[52]}
   );
   gpc615_5 gpc3003 (
      {stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89], stage1_9[90]},
      {stage1_10[52]},
      {stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99], stage1_11[100], stage1_11[101]},
      {stage2_13[16],stage2_12[22],stage2_11[23],stage2_10[39],stage2_9[53]}
   );
   gpc615_5 gpc3004 (
      {stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage1_10[53]},
      {stage1_11[102], stage1_11[103], stage1_11[104], stage1_11[105], stage1_11[106], stage1_11[107]},
      {stage2_13[17],stage2_12[23],stage2_11[24],stage2_10[40],stage2_9[54]}
   );
   gpc615_5 gpc3005 (
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100]},
      {stage1_10[54]},
      {stage1_11[108], stage1_11[109], stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113]},
      {stage2_13[18],stage2_12[24],stage2_11[25],stage2_10[41],stage2_9[55]}
   );
   gpc615_5 gpc3006 (
      {stage1_9[101], stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105]},
      {stage1_10[55]},
      {stage1_11[114], stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage2_13[19],stage2_12[25],stage2_11[26],stage2_10[42],stage2_9[56]}
   );
   gpc615_5 gpc3007 (
      {stage1_9[106], stage1_9[107], stage1_9[108], stage1_9[109], stage1_9[110]},
      {stage1_10[56]},
      {stage1_11[120], stage1_11[121], stage1_11[122], stage1_11[123], stage1_11[124], stage1_11[125]},
      {stage2_13[20],stage2_12[26],stage2_11[27],stage2_10[43],stage2_9[57]}
   );
   gpc615_5 gpc3008 (
      {stage1_9[111], stage1_9[112], stage1_9[113], stage1_9[114], stage1_9[115]},
      {stage1_10[57]},
      {stage1_11[126], stage1_11[127], stage1_11[128], stage1_11[129], stage1_11[130], stage1_11[131]},
      {stage2_13[21],stage2_12[27],stage2_11[28],stage2_10[44],stage2_9[58]}
   );
   gpc615_5 gpc3009 (
      {stage1_9[116], stage1_9[117], stage1_9[118], stage1_9[119], 1'b0},
      {stage1_10[58]},
      {stage1_11[132], stage1_11[133], stage1_11[134], stage1_11[135], stage1_11[136], stage1_11[137]},
      {stage2_13[22],stage2_12[28],stage2_11[29],stage2_10[45],stage2_9[59]}
   );
   gpc606_5 gpc3010 (
      {stage1_10[59], stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[23],stage2_12[29],stage2_11[30],stage2_10[46]}
   );
   gpc606_5 gpc3011 (
      {stage1_10[65], stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[24],stage2_12[30],stage2_11[31],stage2_10[47]}
   );
   gpc606_5 gpc3012 (
      {stage1_10[71], stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[25],stage2_12[31],stage2_11[32],stage2_10[48]}
   );
   gpc606_5 gpc3013 (
      {stage1_10[77], stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[26],stage2_12[32],stage2_11[33],stage2_10[49]}
   );
   gpc606_5 gpc3014 (
      {stage1_10[83], stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[27],stage2_12[33],stage2_11[34],stage2_10[50]}
   );
   gpc606_5 gpc3015 (
      {stage1_10[89], stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[28],stage2_12[34],stage2_11[35],stage2_10[51]}
   );
   gpc606_5 gpc3016 (
      {stage1_10[95], stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[29],stage2_12[35],stage2_11[36],stage2_10[52]}
   );
   gpc606_5 gpc3017 (
      {stage1_10[101], stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[30],stage2_12[36],stage2_11[37],stage2_10[53]}
   );
   gpc606_5 gpc3018 (
      {stage1_10[107], stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[31],stage2_12[37],stage2_11[38],stage2_10[54]}
   );
   gpc606_5 gpc3019 (
      {stage1_10[113], stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[32],stage2_12[38],stage2_11[39],stage2_10[55]}
   );
   gpc606_5 gpc3020 (
      {stage1_10[119], stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[33],stage2_12[39],stage2_11[40],stage2_10[56]}
   );
   gpc606_5 gpc3021 (
      {stage1_10[125], stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[34],stage2_12[40],stage2_11[41],stage2_10[57]}
   );
   gpc606_5 gpc3022 (
      {stage1_10[131], stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[35],stage2_12[41],stage2_11[42],stage2_10[58]}
   );
   gpc615_5 gpc3023 (
      {stage1_10[137], stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141]},
      {stage1_11[138]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[36],stage2_12[42],stage2_11[43],stage2_10[59]}
   );
   gpc615_5 gpc3024 (
      {stage1_10[142], stage1_10[143], stage1_10[144], stage1_10[145], stage1_10[146]},
      {stage1_11[139]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[37],stage2_12[43],stage2_11[44],stage2_10[60]}
   );
   gpc1406_5 gpc3025 (
      {stage1_11[140], stage1_11[141], stage1_11[142], stage1_11[143], stage1_11[144], stage1_11[145]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[15],stage2_13[38],stage2_12[44],stage2_11[45]}
   );
   gpc606_5 gpc3026 (
      {stage1_11[146], stage1_11[147], stage1_11[148], stage1_11[149], stage1_11[150], stage1_11[151]},
      {stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9]},
      {stage2_15[1],stage2_14[16],stage2_13[39],stage2_12[45],stage2_11[46]}
   );
   gpc606_5 gpc3027 (
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[2],stage2_14[17],stage2_13[40],stage2_12[46]}
   );
   gpc606_5 gpc3028 (
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[3],stage2_14[18],stage2_13[41],stage2_12[47]}
   );
   gpc606_5 gpc3029 (
      {stage1_12[102], stage1_12[103], stage1_12[104], stage1_12[105], stage1_12[106], stage1_12[107]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage2_16[2],stage2_15[4],stage2_14[19],stage2_13[42],stage2_12[48]}
   );
   gpc606_5 gpc3030 (
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24]},
      {stage2_16[3],stage2_15[5],stage2_14[20],stage2_13[43],stage2_12[49]}
   );
   gpc606_5 gpc3031 (
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30]},
      {stage2_16[4],stage2_15[6],stage2_14[21],stage2_13[44],stage2_12[50]}
   );
   gpc606_5 gpc3032 (
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36]},
      {stage2_16[5],stage2_15[7],stage2_14[22],stage2_13[45],stage2_12[51]}
   );
   gpc606_5 gpc3033 (
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42]},
      {stage2_16[6],stage2_15[8],stage2_14[23],stage2_13[46],stage2_12[52]}
   );
   gpc606_5 gpc3034 (
      {stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[7],stage2_15[9],stage2_14[24],stage2_13[47]}
   );
   gpc606_5 gpc3035 (
      {stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[8],stage2_15[10],stage2_14[25],stage2_13[48]}
   );
   gpc606_5 gpc3036 (
      {stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[9],stage2_15[11],stage2_14[26],stage2_13[49]}
   );
   gpc606_5 gpc3037 (
      {stage1_13[28], stage1_13[29], stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[10],stage2_15[12],stage2_14[27],stage2_13[50]}
   );
   gpc606_5 gpc3038 (
      {stage1_13[34], stage1_13[35], stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[11],stage2_15[13],stage2_14[28],stage2_13[51]}
   );
   gpc606_5 gpc3039 (
      {stage1_13[40], stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[12],stage2_15[14],stage2_14[29],stage2_13[52]}
   );
   gpc606_5 gpc3040 (
      {stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[13],stage2_15[15],stage2_14[30],stage2_13[53]}
   );
   gpc606_5 gpc3041 (
      {stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[14],stage2_15[16],stage2_14[31],stage2_13[54]}
   );
   gpc606_5 gpc3042 (
      {stage1_13[58], stage1_13[59], stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[15],stage2_15[17],stage2_14[32],stage2_13[55]}
   );
   gpc606_5 gpc3043 (
      {stage1_13[64], stage1_13[65], stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[16],stage2_15[18],stage2_14[33],stage2_13[56]}
   );
   gpc606_5 gpc3044 (
      {stage1_13[70], stage1_13[71], stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[17],stage2_15[19],stage2_14[34],stage2_13[57]}
   );
   gpc606_5 gpc3045 (
      {stage1_13[76], stage1_13[77], stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[18],stage2_15[20],stage2_14[35],stage2_13[58]}
   );
   gpc606_5 gpc3046 (
      {stage1_13[82], stage1_13[83], stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[19],stage2_15[21],stage2_14[36],stage2_13[59]}
   );
   gpc606_5 gpc3047 (
      {stage1_13[88], stage1_13[89], stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[20],stage2_15[22],stage2_14[37],stage2_13[60]}
   );
   gpc606_5 gpc3048 (
      {stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[14],stage2_16[21],stage2_15[23],stage2_14[38]}
   );
   gpc606_5 gpc3049 (
      {stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[15],stage2_16[22],stage2_15[24],stage2_14[39]}
   );
   gpc606_5 gpc3050 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59], stage1_14[60]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[16],stage2_16[23],stage2_15[25],stage2_14[40]}
   );
   gpc606_5 gpc3051 (
      {stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65], stage1_14[66]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[17],stage2_16[24],stage2_15[26],stage2_14[41]}
   );
   gpc606_5 gpc3052 (
      {stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71], stage1_14[72]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[18],stage2_16[25],stage2_15[27],stage2_14[42]}
   );
   gpc606_5 gpc3053 (
      {stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77], stage1_14[78]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[19],stage2_16[26],stage2_15[28],stage2_14[43]}
   );
   gpc606_5 gpc3054 (
      {stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83], stage1_14[84]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[20],stage2_16[27],stage2_15[29],stage2_14[44]}
   );
   gpc615_5 gpc3055 (
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88]},
      {stage1_16[42]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[7],stage2_17[21],stage2_16[28],stage2_15[30]}
   );
   gpc207_4 gpc3056 (
      {stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49]},
      {stage1_18[0], stage1_18[1]},
      {stage2_19[1],stage2_18[8],stage2_17[22],stage2_16[29]}
   );
   gpc606_5 gpc3057 (
      {stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55]},
      {stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5], stage1_18[6], stage1_18[7]},
      {stage2_20[0],stage2_19[2],stage2_18[9],stage2_17[23],stage2_16[30]}
   );
   gpc606_5 gpc3058 (
      {stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61]},
      {stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11], stage1_18[12], stage1_18[13]},
      {stage2_20[1],stage2_19[3],stage2_18[10],stage2_17[24],stage2_16[31]}
   );
   gpc606_5 gpc3059 (
      {stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67]},
      {stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17], stage1_18[18], stage1_18[19]},
      {stage2_20[2],stage2_19[4],stage2_18[11],stage2_17[25],stage2_16[32]}
   );
   gpc606_5 gpc3060 (
      {stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73]},
      {stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23], stage1_18[24], stage1_18[25]},
      {stage2_20[3],stage2_19[5],stage2_18[12],stage2_17[26],stage2_16[33]}
   );
   gpc606_5 gpc3061 (
      {stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79]},
      {stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29], stage1_18[30], stage1_18[31]},
      {stage2_20[4],stage2_19[6],stage2_18[13],stage2_17[27],stage2_16[34]}
   );
   gpc606_5 gpc3062 (
      {stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85]},
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35], stage1_18[36], stage1_18[37]},
      {stage2_20[5],stage2_19[7],stage2_18[14],stage2_17[28],stage2_16[35]}
   );
   gpc606_5 gpc3063 (
      {stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89], stage1_16[90], stage1_16[91]},
      {stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41], stage1_18[42], stage1_18[43]},
      {stage2_20[6],stage2_19[8],stage2_18[15],stage2_17[29],stage2_16[36]}
   );
   gpc606_5 gpc3064 (
      {stage1_16[92], stage1_16[93], stage1_16[94], stage1_16[95], stage1_16[96], stage1_16[97]},
      {stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47], stage1_18[48], stage1_18[49]},
      {stage2_20[7],stage2_19[9],stage2_18[16],stage2_17[30],stage2_16[37]}
   );
   gpc606_5 gpc3065 (
      {stage1_16[98], stage1_16[99], stage1_16[100], stage1_16[101], stage1_16[102], stage1_16[103]},
      {stage1_18[50], stage1_18[51], stage1_18[52], stage1_18[53], stage1_18[54], stage1_18[55]},
      {stage2_20[8],stage2_19[10],stage2_18[17],stage2_17[31],stage2_16[38]}
   );
   gpc606_5 gpc3066 (
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[9],stage2_19[11],stage2_18[18],stage2_17[32]}
   );
   gpc606_5 gpc3067 (
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[10],stage2_19[12],stage2_18[19],stage2_17[33]}
   );
   gpc606_5 gpc3068 (
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[11],stage2_19[13],stage2_18[20],stage2_17[34]}
   );
   gpc606_5 gpc3069 (
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage2_21[3],stage2_20[12],stage2_19[14],stage2_18[21],stage2_17[35]}
   );
   gpc606_5 gpc3070 (
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28], stage1_19[29]},
      {stage2_21[4],stage2_20[13],stage2_19[15],stage2_18[22],stage2_17[36]}
   );
   gpc606_5 gpc3071 (
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35]},
      {stage2_21[5],stage2_20[14],stage2_19[16],stage2_18[23],stage2_17[37]}
   );
   gpc606_5 gpc3072 (
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage1_19[36], stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage2_21[6],stage2_20[15],stage2_19[17],stage2_18[24],stage2_17[38]}
   );
   gpc606_5 gpc3073 (
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage1_19[42], stage1_19[43], stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47]},
      {stage2_21[7],stage2_20[16],stage2_19[18],stage2_18[25],stage2_17[39]}
   );
   gpc606_5 gpc3074 (
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage1_19[48], stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage2_21[8],stage2_20[17],stage2_19[19],stage2_18[26],stage2_17[40]}
   );
   gpc606_5 gpc3075 (
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], stage1_17[64], stage1_17[65]},
      {stage1_19[54], stage1_19[55], stage1_19[56], stage1_19[57], stage1_19[58], stage1_19[59]},
      {stage2_21[9],stage2_20[18],stage2_19[20],stage2_18[27],stage2_17[41]}
   );
   gpc606_5 gpc3076 (
      {stage1_17[66], stage1_17[67], stage1_17[68], stage1_17[69], stage1_17[70], stage1_17[71]},
      {stage1_19[60], stage1_19[61], stage1_19[62], stage1_19[63], stage1_19[64], stage1_19[65]},
      {stage2_21[10],stage2_20[19],stage2_19[21],stage2_18[28],stage2_17[42]}
   );
   gpc606_5 gpc3077 (
      {stage1_17[72], stage1_17[73], stage1_17[74], stage1_17[75], stage1_17[76], stage1_17[77]},
      {stage1_19[66], stage1_19[67], stage1_19[68], stage1_19[69], stage1_19[70], stage1_19[71]},
      {stage2_21[11],stage2_20[20],stage2_19[22],stage2_18[29],stage2_17[43]}
   );
   gpc606_5 gpc3078 (
      {stage1_17[78], stage1_17[79], stage1_17[80], stage1_17[81], stage1_17[82], stage1_17[83]},
      {stage1_19[72], stage1_19[73], stage1_19[74], stage1_19[75], stage1_19[76], stage1_19[77]},
      {stage2_21[12],stage2_20[21],stage2_19[23],stage2_18[30],stage2_17[44]}
   );
   gpc606_5 gpc3079 (
      {stage1_17[84], stage1_17[85], stage1_17[86], stage1_17[87], stage1_17[88], stage1_17[89]},
      {stage1_19[78], stage1_19[79], stage1_19[80], stage1_19[81], stage1_19[82], stage1_19[83]},
      {stage2_21[13],stage2_20[22],stage2_19[24],stage2_18[31],stage2_17[45]}
   );
   gpc606_5 gpc3080 (
      {stage1_17[90], stage1_17[91], stage1_17[92], stage1_17[93], stage1_17[94], stage1_17[95]},
      {stage1_19[84], stage1_19[85], stage1_19[86], stage1_19[87], stage1_19[88], stage1_19[89]},
      {stage2_21[14],stage2_20[23],stage2_19[25],stage2_18[32],stage2_17[46]}
   );
   gpc606_5 gpc3081 (
      {stage1_17[96], stage1_17[97], stage1_17[98], stage1_17[99], stage1_17[100], stage1_17[101]},
      {stage1_19[90], stage1_19[91], stage1_19[92], stage1_19[93], stage1_19[94], stage1_19[95]},
      {stage2_21[15],stage2_20[24],stage2_19[26],stage2_18[33],stage2_17[47]}
   );
   gpc615_5 gpc3082 (
      {stage1_18[56], stage1_18[57], stage1_18[58], stage1_18[59], stage1_18[60]},
      {stage1_19[96]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[16],stage2_20[25],stage2_19[27],stage2_18[34]}
   );
   gpc615_5 gpc3083 (
      {stage1_18[61], stage1_18[62], stage1_18[63], stage1_18[64], stage1_18[65]},
      {stage1_19[97]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[17],stage2_20[26],stage2_19[28],stage2_18[35]}
   );
   gpc615_5 gpc3084 (
      {stage1_18[66], stage1_18[67], stage1_18[68], stage1_18[69], stage1_18[70]},
      {stage1_19[98]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[18],stage2_20[27],stage2_19[29],stage2_18[36]}
   );
   gpc615_5 gpc3085 (
      {stage1_19[99], stage1_19[100], stage1_19[101], stage1_19[102], stage1_19[103]},
      {stage1_20[18]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[19],stage2_20[28],stage2_19[30]}
   );
   gpc615_5 gpc3086 (
      {stage1_19[104], stage1_19[105], stage1_19[106], stage1_19[107], stage1_19[108]},
      {stage1_20[19]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[4],stage2_21[20],stage2_20[29],stage2_19[31]}
   );
   gpc615_5 gpc3087 (
      {stage1_19[109], stage1_19[110], stage1_19[111], stage1_19[112], stage1_19[113]},
      {stage1_20[20]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[5],stage2_21[21],stage2_20[30],stage2_19[32]}
   );
   gpc615_5 gpc3088 (
      {stage1_19[114], stage1_19[115], stage1_19[116], stage1_19[117], stage1_19[118]},
      {stage1_20[21]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[6],stage2_21[22],stage2_20[31],stage2_19[33]}
   );
   gpc615_5 gpc3089 (
      {stage1_19[119], stage1_19[120], stage1_19[121], stage1_19[122], stage1_19[123]},
      {stage1_20[22]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[7],stage2_21[23],stage2_20[32],stage2_19[34]}
   );
   gpc606_5 gpc3090 (
      {stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[5],stage2_22[8],stage2_21[24],stage2_20[33]}
   );
   gpc606_5 gpc3091 (
      {stage1_20[29], stage1_20[30], stage1_20[31], stage1_20[32], stage1_20[33], stage1_20[34]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[6],stage2_22[9],stage2_21[25],stage2_20[34]}
   );
   gpc606_5 gpc3092 (
      {stage1_20[35], stage1_20[36], stage1_20[37], stage1_20[38], stage1_20[39], stage1_20[40]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[7],stage2_22[10],stage2_21[26],stage2_20[35]}
   );
   gpc606_5 gpc3093 (
      {stage1_20[41], stage1_20[42], stage1_20[43], stage1_20[44], stage1_20[45], stage1_20[46]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[8],stage2_22[11],stage2_21[27],stage2_20[36]}
   );
   gpc606_5 gpc3094 (
      {stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50], stage1_20[51], stage1_20[52]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[9],stage2_22[12],stage2_21[28],stage2_20[37]}
   );
   gpc606_5 gpc3095 (
      {stage1_20[53], stage1_20[54], stage1_20[55], stage1_20[56], stage1_20[57], stage1_20[58]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[10],stage2_22[13],stage2_21[29],stage2_20[38]}
   );
   gpc606_5 gpc3096 (
      {stage1_20[59], stage1_20[60], stage1_20[61], stage1_20[62], stage1_20[63], stage1_20[64]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[11],stage2_22[14],stage2_21[30],stage2_20[39]}
   );
   gpc606_5 gpc3097 (
      {stage1_20[65], stage1_20[66], stage1_20[67], stage1_20[68], stage1_20[69], stage1_20[70]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[12],stage2_22[15],stage2_21[31],stage2_20[40]}
   );
   gpc606_5 gpc3098 (
      {stage1_20[71], stage1_20[72], stage1_20[73], stage1_20[74], stage1_20[75], stage1_20[76]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[13],stage2_22[16],stage2_21[32],stage2_20[41]}
   );
   gpc606_5 gpc3099 (
      {stage1_20[77], stage1_20[78], stage1_20[79], stage1_20[80], stage1_20[81], stage1_20[82]},
      {stage1_22[54], stage1_22[55], stage1_22[56], stage1_22[57], stage1_22[58], stage1_22[59]},
      {stage2_24[9],stage2_23[14],stage2_22[17],stage2_21[33],stage2_20[42]}
   );
   gpc606_5 gpc3100 (
      {stage1_20[83], stage1_20[84], stage1_20[85], stage1_20[86], stage1_20[87], stage1_20[88]},
      {stage1_22[60], stage1_22[61], stage1_22[62], stage1_22[63], stage1_22[64], stage1_22[65]},
      {stage2_24[10],stage2_23[15],stage2_22[18],stage2_21[34],stage2_20[43]}
   );
   gpc606_5 gpc3101 (
      {stage1_20[89], stage1_20[90], stage1_20[91], stage1_20[92], stage1_20[93], stage1_20[94]},
      {stage1_22[66], stage1_22[67], stage1_22[68], stage1_22[69], stage1_22[70], stage1_22[71]},
      {stage2_24[11],stage2_23[16],stage2_22[19],stage2_21[35],stage2_20[44]}
   );
   gpc606_5 gpc3102 (
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[12],stage2_23[17],stage2_22[20],stage2_21[36]}
   );
   gpc606_5 gpc3103 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[13],stage2_23[18],stage2_22[21],stage2_21[37]}
   );
   gpc606_5 gpc3104 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[14],stage2_23[19],stage2_22[22],stage2_21[38]}
   );
   gpc606_5 gpc3105 (
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[15],stage2_23[20],stage2_22[23],stage2_21[39]}
   );
   gpc606_5 gpc3106 (
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage1_23[24], stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage2_25[4],stage2_24[16],stage2_23[21],stage2_22[24],stage2_21[40]}
   );
   gpc606_5 gpc3107 (
      {stage1_21[60], stage1_21[61], stage1_21[62], stage1_21[63], stage1_21[64], stage1_21[65]},
      {stage1_23[30], stage1_23[31], stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35]},
      {stage2_25[5],stage2_24[17],stage2_23[22],stage2_22[25],stage2_21[41]}
   );
   gpc606_5 gpc3108 (
      {stage1_21[66], stage1_21[67], stage1_21[68], stage1_21[69], stage1_21[70], stage1_21[71]},
      {stage1_23[36], stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage2_25[6],stage2_24[18],stage2_23[23],stage2_22[26],stage2_21[42]}
   );
   gpc606_5 gpc3109 (
      {stage1_21[72], stage1_21[73], stage1_21[74], stage1_21[75], stage1_21[76], stage1_21[77]},
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46], stage1_23[47]},
      {stage2_25[7],stage2_24[19],stage2_23[24],stage2_22[27],stage2_21[43]}
   );
   gpc606_5 gpc3110 (
      {stage1_21[78], stage1_21[79], stage1_21[80], stage1_21[81], stage1_21[82], stage1_21[83]},
      {stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51], stage1_23[52], stage1_23[53]},
      {stage2_25[8],stage2_24[20],stage2_23[25],stage2_22[28],stage2_21[44]}
   );
   gpc606_5 gpc3111 (
      {stage1_21[84], stage1_21[85], stage1_21[86], stage1_21[87], stage1_21[88], stage1_21[89]},
      {stage1_23[54], stage1_23[55], stage1_23[56], stage1_23[57], stage1_23[58], stage1_23[59]},
      {stage2_25[9],stage2_24[21],stage2_23[26],stage2_22[29],stage2_21[45]}
   );
   gpc606_5 gpc3112 (
      {stage1_21[90], stage1_21[91], stage1_21[92], stage1_21[93], stage1_21[94], stage1_21[95]},
      {stage1_23[60], stage1_23[61], stage1_23[62], stage1_23[63], stage1_23[64], stage1_23[65]},
      {stage2_25[10],stage2_24[22],stage2_23[27],stage2_22[30],stage2_21[46]}
   );
   gpc606_5 gpc3113 (
      {stage1_21[96], stage1_21[97], stage1_21[98], stage1_21[99], stage1_21[100], stage1_21[101]},
      {stage1_23[66], stage1_23[67], stage1_23[68], stage1_23[69], stage1_23[70], stage1_23[71]},
      {stage2_25[11],stage2_24[23],stage2_23[28],stage2_22[31],stage2_21[47]}
   );
   gpc606_5 gpc3114 (
      {stage1_21[102], stage1_21[103], stage1_21[104], stage1_21[105], stage1_21[106], stage1_21[107]},
      {stage1_23[72], stage1_23[73], stage1_23[74], stage1_23[75], stage1_23[76], stage1_23[77]},
      {stage2_25[12],stage2_24[24],stage2_23[29],stage2_22[32],stage2_21[48]}
   );
   gpc615_5 gpc3115 (
      {stage1_22[72], stage1_22[73], stage1_22[74], stage1_22[75], stage1_22[76]},
      {stage1_23[78]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[13],stage2_24[25],stage2_23[30],stage2_22[33]}
   );
   gpc615_5 gpc3116 (
      {stage1_22[77], stage1_22[78], stage1_22[79], stage1_22[80], stage1_22[81]},
      {stage1_23[79]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[14],stage2_24[26],stage2_23[31],stage2_22[34]}
   );
   gpc615_5 gpc3117 (
      {stage1_22[82], stage1_22[83], stage1_22[84], stage1_22[85], stage1_22[86]},
      {stage1_23[80]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[15],stage2_24[27],stage2_23[32],stage2_22[35]}
   );
   gpc615_5 gpc3118 (
      {stage1_23[81], stage1_23[82], stage1_23[83], stage1_23[84], stage1_23[85]},
      {stage1_24[18]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[3],stage2_25[16],stage2_24[28],stage2_23[33]}
   );
   gpc615_5 gpc3119 (
      {stage1_23[86], stage1_23[87], stage1_23[88], stage1_23[89], stage1_23[90]},
      {stage1_24[19]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[4],stage2_25[17],stage2_24[29],stage2_23[34]}
   );
   gpc615_5 gpc3120 (
      {stage1_23[91], stage1_23[92], stage1_23[93], stage1_23[94], stage1_23[95]},
      {stage1_24[20]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[5],stage2_25[18],stage2_24[30],stage2_23[35]}
   );
   gpc615_5 gpc3121 (
      {stage1_23[96], stage1_23[97], stage1_23[98], stage1_23[99], stage1_23[100]},
      {stage1_24[21]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[6],stage2_25[19],stage2_24[31],stage2_23[36]}
   );
   gpc615_5 gpc3122 (
      {stage1_23[101], stage1_23[102], stage1_23[103], stage1_23[104], stage1_23[105]},
      {stage1_24[22]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[7],stage2_25[20],stage2_24[32],stage2_23[37]}
   );
   gpc1163_5 gpc3123 (
      {stage1_24[23], stage1_24[24], stage1_24[25]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage1_26[0]},
      {stage1_27[0]},
      {stage2_28[0],stage2_27[5],stage2_26[8],stage2_25[21],stage2_24[33]}
   );
   gpc1163_5 gpc3124 (
      {stage1_24[26], stage1_24[27], stage1_24[28]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage1_26[1]},
      {stage1_27[1]},
      {stage2_28[1],stage2_27[6],stage2_26[9],stage2_25[22],stage2_24[34]}
   );
   gpc1163_5 gpc3125 (
      {stage1_24[29], stage1_24[30], stage1_24[31]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage1_26[2]},
      {stage1_27[2]},
      {stage2_28[2],stage2_27[7],stage2_26[10],stage2_25[23],stage2_24[35]}
   );
   gpc1163_5 gpc3126 (
      {stage1_24[32], stage1_24[33], stage1_24[34]},
      {stage1_25[48], stage1_25[49], stage1_25[50], stage1_25[51], stage1_25[52], stage1_25[53]},
      {stage1_26[3]},
      {stage1_27[3]},
      {stage2_28[3],stage2_27[8],stage2_26[11],stage2_25[24],stage2_24[36]}
   );
   gpc615_5 gpc3127 (
      {stage1_24[35], stage1_24[36], stage1_24[37], stage1_24[38], stage1_24[39]},
      {stage1_25[54]},
      {stage1_26[4], stage1_26[5], stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9]},
      {stage2_28[4],stage2_27[9],stage2_26[12],stage2_25[25],stage2_24[37]}
   );
   gpc615_5 gpc3128 (
      {stage1_24[40], stage1_24[41], stage1_24[42], stage1_24[43], stage1_24[44]},
      {stage1_25[55]},
      {stage1_26[10], stage1_26[11], stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15]},
      {stage2_28[5],stage2_27[10],stage2_26[13],stage2_25[26],stage2_24[38]}
   );
   gpc615_5 gpc3129 (
      {stage1_24[45], stage1_24[46], stage1_24[47], stage1_24[48], stage1_24[49]},
      {stage1_25[56]},
      {stage1_26[16], stage1_26[17], stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21]},
      {stage2_28[6],stage2_27[11],stage2_26[14],stage2_25[27],stage2_24[39]}
   );
   gpc615_5 gpc3130 (
      {stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53], stage1_24[54]},
      {stage1_25[57]},
      {stage1_26[22], stage1_26[23], stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27]},
      {stage2_28[7],stage2_27[12],stage2_26[15],stage2_25[28],stage2_24[40]}
   );
   gpc615_5 gpc3131 (
      {stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59]},
      {stage1_25[58]},
      {stage1_26[28], stage1_26[29], stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33]},
      {stage2_28[8],stage2_27[13],stage2_26[16],stage2_25[29],stage2_24[41]}
   );
   gpc615_5 gpc3132 (
      {stage1_24[60], stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64]},
      {stage1_25[59]},
      {stage1_26[34], stage1_26[35], stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39]},
      {stage2_28[9],stage2_27[14],stage2_26[17],stage2_25[30],stage2_24[42]}
   );
   gpc615_5 gpc3133 (
      {stage1_24[65], stage1_24[66], stage1_24[67], stage1_24[68], stage1_24[69]},
      {stage1_25[60]},
      {stage1_26[40], stage1_26[41], stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45]},
      {stage2_28[10],stage2_27[15],stage2_26[18],stage2_25[31],stage2_24[43]}
   );
   gpc615_5 gpc3134 (
      {stage1_24[70], stage1_24[71], stage1_24[72], stage1_24[73], stage1_24[74]},
      {stage1_25[61]},
      {stage1_26[46], stage1_26[47], stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51]},
      {stage2_28[11],stage2_27[16],stage2_26[19],stage2_25[32],stage2_24[44]}
   );
   gpc615_5 gpc3135 (
      {stage1_24[75], stage1_24[76], stage1_24[77], stage1_24[78], stage1_24[79]},
      {stage1_25[62]},
      {stage1_26[52], stage1_26[53], stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57]},
      {stage2_28[12],stage2_27[17],stage2_26[20],stage2_25[33],stage2_24[45]}
   );
   gpc615_5 gpc3136 (
      {stage1_24[80], stage1_24[81], stage1_24[82], stage1_24[83], stage1_24[84]},
      {stage1_25[63]},
      {stage1_26[58], stage1_26[59], stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63]},
      {stage2_28[13],stage2_27[18],stage2_26[21],stage2_25[34],stage2_24[46]}
   );
   gpc615_5 gpc3137 (
      {stage1_24[85], stage1_24[86], stage1_24[87], stage1_24[88], stage1_24[89]},
      {stage1_25[64]},
      {stage1_26[64], stage1_26[65], stage1_26[66], stage1_26[67], stage1_26[68], stage1_26[69]},
      {stage2_28[14],stage2_27[19],stage2_26[22],stage2_25[35],stage2_24[47]}
   );
   gpc615_5 gpc3138 (
      {stage1_24[90], stage1_24[91], stage1_24[92], stage1_24[93], stage1_24[94]},
      {stage1_25[65]},
      {stage1_26[70], stage1_26[71], stage1_26[72], stage1_26[73], stage1_26[74], stage1_26[75]},
      {stage2_28[15],stage2_27[20],stage2_26[23],stage2_25[36],stage2_24[48]}
   );
   gpc615_5 gpc3139 (
      {stage1_24[95], stage1_24[96], stage1_24[97], stage1_24[98], stage1_24[99]},
      {stage1_25[66]},
      {stage1_26[76], stage1_26[77], stage1_26[78], stage1_26[79], stage1_26[80], stage1_26[81]},
      {stage2_28[16],stage2_27[21],stage2_26[24],stage2_25[37],stage2_24[49]}
   );
   gpc615_5 gpc3140 (
      {stage1_24[100], stage1_24[101], stage1_24[102], stage1_24[103], stage1_24[104]},
      {stage1_25[67]},
      {stage1_26[82], stage1_26[83], stage1_26[84], stage1_26[85], stage1_26[86], stage1_26[87]},
      {stage2_28[17],stage2_27[22],stage2_26[25],stage2_25[38],stage2_24[50]}
   );
   gpc615_5 gpc3141 (
      {stage1_24[105], stage1_24[106], stage1_24[107], stage1_24[108], stage1_24[109]},
      {stage1_25[68]},
      {stage1_26[88], stage1_26[89], stage1_26[90], stage1_26[91], stage1_26[92], stage1_26[93]},
      {stage2_28[18],stage2_27[23],stage2_26[26],stage2_25[39],stage2_24[51]}
   );
   gpc606_5 gpc3142 (
      {stage1_25[69], stage1_25[70], stage1_25[71], stage1_25[72], stage1_25[73], stage1_25[74]},
      {stage1_27[4], stage1_27[5], stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9]},
      {stage2_29[0],stage2_28[19],stage2_27[24],stage2_26[27],stage2_25[40]}
   );
   gpc606_5 gpc3143 (
      {stage1_25[75], stage1_25[76], stage1_25[77], stage1_25[78], stage1_25[79], stage1_25[80]},
      {stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15]},
      {stage2_29[1],stage2_28[20],stage2_27[25],stage2_26[28],stage2_25[41]}
   );
   gpc606_5 gpc3144 (
      {stage1_25[81], stage1_25[82], stage1_25[83], stage1_25[84], stage1_25[85], stage1_25[86]},
      {stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21]},
      {stage2_29[2],stage2_28[21],stage2_27[26],stage2_26[29],stage2_25[42]}
   );
   gpc606_5 gpc3145 (
      {stage1_25[87], stage1_25[88], stage1_25[89], stage1_25[90], stage1_25[91], stage1_25[92]},
      {stage1_27[22], stage1_27[23], stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27]},
      {stage2_29[3],stage2_28[22],stage2_27[27],stage2_26[30],stage2_25[43]}
   );
   gpc606_5 gpc3146 (
      {stage1_25[93], stage1_25[94], stage1_25[95], stage1_25[96], stage1_25[97], stage1_25[98]},
      {stage1_27[28], stage1_27[29], stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33]},
      {stage2_29[4],stage2_28[23],stage2_27[28],stage2_26[31],stage2_25[44]}
   );
   gpc606_5 gpc3147 (
      {stage1_25[99], stage1_25[100], stage1_25[101], stage1_25[102], stage1_25[103], stage1_25[104]},
      {stage1_27[34], stage1_27[35], stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39]},
      {stage2_29[5],stage2_28[24],stage2_27[29],stage2_26[32],stage2_25[45]}
   );
   gpc615_5 gpc3148 (
      {stage1_26[94], stage1_26[95], stage1_26[96], stage1_26[97], stage1_26[98]},
      {stage1_27[40]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[6],stage2_28[25],stage2_27[30],stage2_26[33]}
   );
   gpc615_5 gpc3149 (
      {stage1_26[99], stage1_26[100], stage1_26[101], stage1_26[102], stage1_26[103]},
      {stage1_27[41]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[7],stage2_28[26],stage2_27[31],stage2_26[34]}
   );
   gpc615_5 gpc3150 (
      {stage1_26[104], stage1_26[105], stage1_26[106], stage1_26[107], stage1_26[108]},
      {stage1_27[42]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[8],stage2_28[27],stage2_27[32],stage2_26[35]}
   );
   gpc615_5 gpc3151 (
      {stage1_26[109], stage1_26[110], stage1_26[111], stage1_26[112], stage1_26[113]},
      {stage1_27[43]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[9],stage2_28[28],stage2_27[33],stage2_26[36]}
   );
   gpc615_5 gpc3152 (
      {stage1_26[114], stage1_26[115], stage1_26[116], stage1_26[117], stage1_26[118]},
      {stage1_27[44]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[10],stage2_28[29],stage2_27[34],stage2_26[37]}
   );
   gpc615_5 gpc3153 (
      {stage1_26[119], stage1_26[120], stage1_26[121], stage1_26[122], stage1_26[123]},
      {stage1_27[45]},
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage2_30[5],stage2_29[11],stage2_28[30],stage2_27[35],stage2_26[38]}
   );
   gpc615_5 gpc3154 (
      {stage1_26[124], stage1_26[125], stage1_26[126], stage1_26[127], stage1_26[128]},
      {stage1_27[46]},
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage2_30[6],stage2_29[12],stage2_28[31],stage2_27[36],stage2_26[39]}
   );
   gpc606_5 gpc3155 (
      {stage1_27[47], stage1_27[48], stage1_27[49], stage1_27[50], stage1_27[51], stage1_27[52]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[7],stage2_29[13],stage2_28[32],stage2_27[37]}
   );
   gpc615_5 gpc3156 (
      {stage1_27[53], stage1_27[54], stage1_27[55], stage1_27[56], stage1_27[57]},
      {stage1_28[42]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[8],stage2_29[14],stage2_28[33],stage2_27[38]}
   );
   gpc615_5 gpc3157 (
      {stage1_27[58], stage1_27[59], stage1_27[60], stage1_27[61], stage1_27[62]},
      {stage1_28[43]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[9],stage2_29[15],stage2_28[34],stage2_27[39]}
   );
   gpc615_5 gpc3158 (
      {stage1_27[63], stage1_27[64], stage1_27[65], stage1_27[66], stage1_27[67]},
      {stage1_28[44]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[10],stage2_29[16],stage2_28[35],stage2_27[40]}
   );
   gpc615_5 gpc3159 (
      {stage1_27[68], stage1_27[69], stage1_27[70], stage1_27[71], stage1_27[72]},
      {stage1_28[45]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[11],stage2_29[17],stage2_28[36],stage2_27[41]}
   );
   gpc615_5 gpc3160 (
      {stage1_27[73], stage1_27[74], stage1_27[75], stage1_27[76], stage1_27[77]},
      {stage1_28[46]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[12],stage2_29[18],stage2_28[37],stage2_27[42]}
   );
   gpc615_5 gpc3161 (
      {stage1_27[78], stage1_27[79], stage1_27[80], stage1_27[81], stage1_27[82]},
      {stage1_28[47]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[13],stage2_29[19],stage2_28[38],stage2_27[43]}
   );
   gpc615_5 gpc3162 (
      {stage1_27[83], stage1_27[84], stage1_27[85], stage1_27[86], stage1_27[87]},
      {stage1_28[48]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[14],stage2_29[20],stage2_28[39],stage2_27[44]}
   );
   gpc615_5 gpc3163 (
      {stage1_27[88], stage1_27[89], stage1_27[90], stage1_27[91], stage1_27[92]},
      {stage1_28[49]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[15],stage2_29[21],stage2_28[40],stage2_27[45]}
   );
   gpc606_5 gpc3164 (
      {stage1_28[50], stage1_28[51], stage1_28[52], stage1_28[53], stage1_28[54], stage1_28[55]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[9],stage2_30[16],stage2_29[22],stage2_28[41]}
   );
   gpc606_5 gpc3165 (
      {stage1_28[56], stage1_28[57], stage1_28[58], stage1_28[59], stage1_28[60], stage1_28[61]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[10],stage2_30[17],stage2_29[23],stage2_28[42]}
   );
   gpc606_5 gpc3166 (
      {stage1_28[62], stage1_28[63], stage1_28[64], stage1_28[65], stage1_28[66], stage1_28[67]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[11],stage2_30[18],stage2_29[24],stage2_28[43]}
   );
   gpc606_5 gpc3167 (
      {stage1_28[68], stage1_28[69], stage1_28[70], stage1_28[71], stage1_28[72], stage1_28[73]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[12],stage2_30[19],stage2_29[25],stage2_28[44]}
   );
   gpc606_5 gpc3168 (
      {stage1_28[74], stage1_28[75], stage1_28[76], stage1_28[77], stage1_28[78], stage1_28[79]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[13],stage2_30[20],stage2_29[26],stage2_28[45]}
   );
   gpc606_5 gpc3169 (
      {stage1_28[80], stage1_28[81], stage1_28[82], stage1_28[83], stage1_28[84], stage1_28[85]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[14],stage2_30[21],stage2_29[27],stage2_28[46]}
   );
   gpc606_5 gpc3170 (
      {stage1_28[86], stage1_28[87], stage1_28[88], stage1_28[89], stage1_28[90], stage1_28[91]},
      {stage1_30[36], stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage2_32[6],stage2_31[15],stage2_30[22],stage2_29[28],stage2_28[47]}
   );
   gpc606_5 gpc3171 (
      {stage1_28[92], stage1_28[93], stage1_28[94], stage1_28[95], stage1_28[96], stage1_28[97]},
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47]},
      {stage2_32[7],stage2_31[16],stage2_30[23],stage2_29[29],stage2_28[48]}
   );
   gpc606_5 gpc3172 (
      {stage1_28[98], stage1_28[99], stage1_28[100], stage1_28[101], stage1_28[102], stage1_28[103]},
      {stage1_30[48], stage1_30[49], stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53]},
      {stage2_32[8],stage2_31[17],stage2_30[24],stage2_29[30],stage2_28[49]}
   );
   gpc1415_5 gpc3173 (
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58]},
      {stage1_30[54]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3]},
      {stage1_32[0]},
      {stage2_33[0],stage2_32[9],stage2_31[18],stage2_30[25],stage2_29[31]}
   );
   gpc606_5 gpc3174 (
      {stage1_29[59], stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64]},
      {stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9]},
      {stage2_33[1],stage2_32[10],stage2_31[19],stage2_30[26],stage2_29[32]}
   );
   gpc606_5 gpc3175 (
      {stage1_29[65], stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70]},
      {stage1_31[10], stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage2_33[2],stage2_32[11],stage2_31[20],stage2_30[27],stage2_29[33]}
   );
   gpc606_5 gpc3176 (
      {stage1_29[71], stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76]},
      {stage1_31[16], stage1_31[17], stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21]},
      {stage2_33[3],stage2_32[12],stage2_31[21],stage2_30[28],stage2_29[34]}
   );
   gpc606_5 gpc3177 (
      {stage1_29[77], stage1_29[78], stage1_29[79], stage1_29[80], stage1_29[81], stage1_29[82]},
      {stage1_31[22], stage1_31[23], stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27]},
      {stage2_33[4],stage2_32[13],stage2_31[22],stage2_30[29],stage2_29[35]}
   );
   gpc606_5 gpc3178 (
      {stage1_29[83], stage1_29[84], stage1_29[85], stage1_29[86], stage1_29[87], stage1_29[88]},
      {stage1_31[28], stage1_31[29], stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33]},
      {stage2_33[5],stage2_32[14],stage2_31[23],stage2_30[30],stage2_29[36]}
   );
   gpc615_5 gpc3179 (
      {stage1_29[89], stage1_29[90], stage1_29[91], stage1_29[92], stage1_29[93]},
      {stage1_30[55]},
      {stage1_31[34], stage1_31[35], stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39]},
      {stage2_33[6],stage2_32[15],stage2_31[24],stage2_30[31],stage2_29[37]}
   );
   gpc615_5 gpc3180 (
      {stage1_29[94], stage1_29[95], stage1_29[96], stage1_29[97], stage1_29[98]},
      {stage1_30[56]},
      {stage1_31[40], stage1_31[41], stage1_31[42], stage1_31[43], stage1_31[44], stage1_31[45]},
      {stage2_33[7],stage2_32[16],stage2_31[25],stage2_30[32],stage2_29[38]}
   );
   gpc615_5 gpc3181 (
      {stage1_29[99], stage1_29[100], stage1_29[101], stage1_29[102], stage1_29[103]},
      {stage1_30[57]},
      {stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49], stage1_31[50], stage1_31[51]},
      {stage2_33[8],stage2_32[17],stage2_31[26],stage2_30[33],stage2_29[39]}
   );
   gpc615_5 gpc3182 (
      {stage1_30[58], stage1_30[59], stage1_30[60], stage1_30[61], stage1_30[62]},
      {stage1_31[52]},
      {stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5], stage1_32[6]},
      {stage2_34[0],stage2_33[9],stage2_32[18],stage2_31[27],stage2_30[34]}
   );
   gpc615_5 gpc3183 (
      {stage1_30[63], stage1_30[64], stage1_30[65], stage1_30[66], stage1_30[67]},
      {stage1_31[53]},
      {stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11], stage1_32[12]},
      {stage2_34[1],stage2_33[10],stage2_32[19],stage2_31[28],stage2_30[35]}
   );
   gpc615_5 gpc3184 (
      {stage1_31[54], stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58]},
      {stage1_32[13]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[2],stage2_33[11],stage2_32[20],stage2_31[29]}
   );
   gpc615_5 gpc3185 (
      {stage1_31[59], stage1_31[60], stage1_31[61], stage1_31[62], stage1_31[63]},
      {stage1_32[14]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[3],stage2_33[12],stage2_32[21],stage2_31[30]}
   );
   gpc615_5 gpc3186 (
      {stage1_31[64], stage1_31[65], stage1_31[66], stage1_31[67], stage1_31[68]},
      {stage1_32[15]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[4],stage2_33[13],stage2_32[22],stage2_31[31]}
   );
   gpc615_5 gpc3187 (
      {stage1_31[69], stage1_31[70], stage1_31[71], stage1_31[72], stage1_31[73]},
      {stage1_32[16]},
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage2_35[3],stage2_34[5],stage2_33[14],stage2_32[23],stage2_31[32]}
   );
   gpc615_5 gpc3188 (
      {stage1_31[74], stage1_31[75], stage1_31[76], stage1_31[77], stage1_31[78]},
      {stage1_32[17]},
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage2_35[4],stage2_34[6],stage2_33[15],stage2_32[24],stage2_31[33]}
   );
   gpc615_5 gpc3189 (
      {stage1_31[79], stage1_31[80], stage1_31[81], stage1_31[82], stage1_31[83]},
      {stage1_32[18]},
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage2_35[5],stage2_34[7],stage2_33[16],stage2_32[25],stage2_31[34]}
   );
   gpc615_5 gpc3190 (
      {stage1_31[84], stage1_31[85], stage1_31[86], stage1_31[87], stage1_31[88]},
      {stage1_32[19]},
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41]},
      {stage2_35[6],stage2_34[8],stage2_33[17],stage2_32[26],stage2_31[35]}
   );
   gpc615_5 gpc3191 (
      {stage1_31[89], stage1_31[90], stage1_31[91], stage1_31[92], stage1_31[93]},
      {stage1_32[20]},
      {stage1_33[42], stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47]},
      {stage2_35[7],stage2_34[9],stage2_33[18],stage2_32[27],stage2_31[36]}
   );
   gpc615_5 gpc3192 (
      {stage1_31[94], stage1_31[95], stage1_31[96], stage1_31[97], stage1_31[98]},
      {stage1_32[21]},
      {stage1_33[48], stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53]},
      {stage2_35[8],stage2_34[10],stage2_33[19],stage2_32[28],stage2_31[37]}
   );
   gpc606_5 gpc3193 (
      {stage1_32[22], stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[9],stage2_34[11],stage2_33[20],stage2_32[29]}
   );
   gpc606_5 gpc3194 (
      {stage1_32[28], stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[10],stage2_34[12],stage2_33[21],stage2_32[30]}
   );
   gpc606_5 gpc3195 (
      {stage1_32[34], stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[11],stage2_34[13],stage2_33[22],stage2_32[31]}
   );
   gpc606_5 gpc3196 (
      {stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[12],stage2_34[14],stage2_33[23],stage2_32[32]}
   );
   gpc606_5 gpc3197 (
      {stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[13],stage2_34[15],stage2_33[24],stage2_32[33]}
   );
   gpc606_5 gpc3198 (
      {stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57]},
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage2_36[5],stage2_35[14],stage2_34[16],stage2_33[25],stage2_32[34]}
   );
   gpc606_5 gpc3199 (
      {stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63]},
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40], stage1_34[41]},
      {stage2_36[6],stage2_35[15],stage2_34[17],stage2_33[26],stage2_32[35]}
   );
   gpc606_5 gpc3200 (
      {stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69]},
      {stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45], stage1_34[46], stage1_34[47]},
      {stage2_36[7],stage2_35[16],stage2_34[18],stage2_33[27],stage2_32[36]}
   );
   gpc606_5 gpc3201 (
      {stage1_32[70], stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75]},
      {stage1_34[48], stage1_34[49], stage1_34[50], stage1_34[51], stage1_34[52], stage1_34[53]},
      {stage2_36[8],stage2_35[17],stage2_34[19],stage2_33[28],stage2_32[37]}
   );
   gpc606_5 gpc3202 (
      {stage1_32[76], stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81]},
      {stage1_34[54], stage1_34[55], stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59]},
      {stage2_36[9],stage2_35[18],stage2_34[20],stage2_33[29],stage2_32[38]}
   );
   gpc606_5 gpc3203 (
      {stage1_32[82], stage1_32[83], stage1_32[84], stage1_32[85], stage1_32[86], stage1_32[87]},
      {stage1_34[60], stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65]},
      {stage2_36[10],stage2_35[19],stage2_34[21],stage2_33[30],stage2_32[39]}
   );
   gpc606_5 gpc3204 (
      {stage1_32[88], stage1_32[89], stage1_32[90], stage1_32[91], stage1_32[92], stage1_32[93]},
      {stage1_34[66], stage1_34[67], stage1_34[68], stage1_34[69], stage1_34[70], stage1_34[71]},
      {stage2_36[11],stage2_35[20],stage2_34[22],stage2_33[31],stage2_32[40]}
   );
   gpc606_5 gpc3205 (
      {stage1_32[94], stage1_32[95], stage1_32[96], stage1_32[97], stage1_32[98], stage1_32[99]},
      {stage1_34[72], stage1_34[73], stage1_34[74], stage1_34[75], stage1_34[76], stage1_34[77]},
      {stage2_36[12],stage2_35[21],stage2_34[23],stage2_33[32],stage2_32[41]}
   );
   gpc606_5 gpc3206 (
      {stage1_32[100], stage1_32[101], stage1_32[102], stage1_32[103], stage1_32[104], stage1_32[105]},
      {stage1_34[78], stage1_34[79], stage1_34[80], stage1_34[81], stage1_34[82], stage1_34[83]},
      {stage2_36[13],stage2_35[22],stage2_34[24],stage2_33[33],stage2_32[42]}
   );
   gpc606_5 gpc3207 (
      {stage1_32[106], stage1_32[107], stage1_32[108], stage1_32[109], stage1_32[110], stage1_32[111]},
      {stage1_34[84], stage1_34[85], stage1_34[86], stage1_34[87], stage1_34[88], stage1_34[89]},
      {stage2_36[14],stage2_35[23],stage2_34[25],stage2_33[34],stage2_32[43]}
   );
   gpc606_5 gpc3208 (
      {stage1_33[54], stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[15],stage2_35[24],stage2_34[26],stage2_33[35]}
   );
   gpc606_5 gpc3209 (
      {stage1_33[60], stage1_33[61], stage1_33[62], stage1_33[63], stage1_33[64], stage1_33[65]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[16],stage2_35[25],stage2_34[27],stage2_33[36]}
   );
   gpc606_5 gpc3210 (
      {stage1_33[66], stage1_33[67], stage1_33[68], stage1_33[69], stage1_33[70], stage1_33[71]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[17],stage2_35[26],stage2_34[28],stage2_33[37]}
   );
   gpc606_5 gpc3211 (
      {stage1_33[72], stage1_33[73], stage1_33[74], stage1_33[75], stage1_33[76], stage1_33[77]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[18],stage2_35[27],stage2_34[29],stage2_33[38]}
   );
   gpc606_5 gpc3212 (
      {stage1_33[78], stage1_33[79], stage1_33[80], stage1_33[81], stage1_33[82], stage1_33[83]},
      {stage1_35[24], stage1_35[25], stage1_35[26], stage1_35[27], stage1_35[28], stage1_35[29]},
      {stage2_37[4],stage2_36[19],stage2_35[28],stage2_34[30],stage2_33[39]}
   );
   gpc606_5 gpc3213 (
      {stage1_33[84], stage1_33[85], stage1_33[86], stage1_33[87], stage1_33[88], stage1_33[89]},
      {stage1_35[30], stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage2_37[5],stage2_36[20],stage2_35[29],stage2_34[31],stage2_33[40]}
   );
   gpc606_5 gpc3214 (
      {stage1_33[90], stage1_33[91], stage1_33[92], stage1_33[93], stage1_33[94], stage1_33[95]},
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41]},
      {stage2_37[6],stage2_36[21],stage2_35[30],stage2_34[32],stage2_33[41]}
   );
   gpc606_5 gpc3215 (
      {stage1_33[96], stage1_33[97], stage1_33[98], stage1_33[99], stage1_33[100], stage1_33[101]},
      {stage1_35[42], stage1_35[43], stage1_35[44], stage1_35[45], stage1_35[46], stage1_35[47]},
      {stage2_37[7],stage2_36[22],stage2_35[31],stage2_34[33],stage2_33[42]}
   );
   gpc615_5 gpc3216 (
      {stage1_34[90], stage1_34[91], stage1_34[92], stage1_34[93], stage1_34[94]},
      {stage1_35[48]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[8],stage2_36[23],stage2_35[32],stage2_34[34]}
   );
   gpc615_5 gpc3217 (
      {stage1_34[95], stage1_34[96], stage1_34[97], stage1_34[98], stage1_34[99]},
      {stage1_35[49]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[9],stage2_36[24],stage2_35[33],stage2_34[35]}
   );
   gpc615_5 gpc3218 (
      {stage1_34[100], stage1_34[101], stage1_34[102], stage1_34[103], 1'b0},
      {stage1_35[50]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[10],stage2_36[25],stage2_35[34],stage2_34[36]}
   );
   gpc615_5 gpc3219 (
      {stage1_35[51], stage1_35[52], stage1_35[53], stage1_35[54], stage1_35[55]},
      {stage1_36[18]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[3],stage2_37[11],stage2_36[26],stage2_35[35]}
   );
   gpc615_5 gpc3220 (
      {stage1_35[56], stage1_35[57], stage1_35[58], stage1_35[59], stage1_35[60]},
      {stage1_36[19]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[4],stage2_37[12],stage2_36[27],stage2_35[36]}
   );
   gpc615_5 gpc3221 (
      {stage1_35[61], stage1_35[62], stage1_35[63], stage1_35[64], stage1_35[65]},
      {stage1_36[20]},
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage2_39[2],stage2_38[5],stage2_37[13],stage2_36[28],stage2_35[37]}
   );
   gpc615_5 gpc3222 (
      {stage1_35[66], stage1_35[67], stage1_35[68], stage1_35[69], stage1_35[70]},
      {stage1_36[21]},
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage2_39[3],stage2_38[6],stage2_37[14],stage2_36[29],stage2_35[38]}
   );
   gpc615_5 gpc3223 (
      {stage1_35[71], stage1_35[72], stage1_35[73], stage1_35[74], stage1_35[75]},
      {stage1_36[22]},
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28], stage1_37[29]},
      {stage2_39[4],stage2_38[7],stage2_37[15],stage2_36[30],stage2_35[39]}
   );
   gpc615_5 gpc3224 (
      {stage1_35[76], stage1_35[77], stage1_35[78], stage1_35[79], stage1_35[80]},
      {stage1_36[23]},
      {stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33], stage1_37[34], stage1_37[35]},
      {stage2_39[5],stage2_38[8],stage2_37[16],stage2_36[31],stage2_35[40]}
   );
   gpc615_5 gpc3225 (
      {stage1_35[81], stage1_35[82], stage1_35[83], stage1_35[84], stage1_35[85]},
      {stage1_36[24]},
      {stage1_37[36], stage1_37[37], stage1_37[38], stage1_37[39], stage1_37[40], stage1_37[41]},
      {stage2_39[6],stage2_38[9],stage2_37[17],stage2_36[32],stage2_35[41]}
   );
   gpc615_5 gpc3226 (
      {stage1_35[86], stage1_35[87], stage1_35[88], stage1_35[89], stage1_35[90]},
      {stage1_36[25]},
      {stage1_37[42], stage1_37[43], stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47]},
      {stage2_39[7],stage2_38[10],stage2_37[18],stage2_36[33],stage2_35[42]}
   );
   gpc615_5 gpc3227 (
      {stage1_35[91], stage1_35[92], stage1_35[93], stage1_35[94], stage1_35[95]},
      {stage1_36[26]},
      {stage1_37[48], stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage2_39[8],stage2_38[11],stage2_37[19],stage2_36[34],stage2_35[43]}
   );
   gpc615_5 gpc3228 (
      {stage1_35[96], stage1_35[97], stage1_35[98], stage1_35[99], stage1_35[100]},
      {stage1_36[27]},
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58], stage1_37[59]},
      {stage2_39[9],stage2_38[12],stage2_37[20],stage2_36[35],stage2_35[44]}
   );
   gpc615_5 gpc3229 (
      {stage1_35[101], stage1_35[102], stage1_35[103], stage1_35[104], stage1_35[105]},
      {stage1_36[28]},
      {stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63], stage1_37[64], stage1_37[65]},
      {stage2_39[10],stage2_38[13],stage2_37[21],stage2_36[36],stage2_35[45]}
   );
   gpc135_4 gpc3230 (
      {stage1_36[29], stage1_36[30], stage1_36[31], stage1_36[32], stage1_36[33]},
      {stage1_37[66], stage1_37[67], stage1_37[68]},
      {stage1_38[0]},
      {stage2_39[11],stage2_38[14],stage2_37[22],stage2_36[37]}
   );
   gpc135_4 gpc3231 (
      {stage1_36[34], stage1_36[35], stage1_36[36], stage1_36[37], stage1_36[38]},
      {stage1_37[69], stage1_37[70], stage1_37[71]},
      {stage1_38[1]},
      {stage2_39[12],stage2_38[15],stage2_37[23],stage2_36[38]}
   );
   gpc135_4 gpc3232 (
      {stage1_36[39], stage1_36[40], stage1_36[41], stage1_36[42], stage1_36[43]},
      {stage1_37[72], stage1_37[73], stage1_37[74]},
      {stage1_38[2]},
      {stage2_39[13],stage2_38[16],stage2_37[24],stage2_36[39]}
   );
   gpc135_4 gpc3233 (
      {stage1_36[44], stage1_36[45], stage1_36[46], stage1_36[47], stage1_36[48]},
      {stage1_37[75], stage1_37[76], stage1_37[77]},
      {stage1_38[3]},
      {stage2_39[14],stage2_38[17],stage2_37[25],stage2_36[40]}
   );
   gpc135_4 gpc3234 (
      {stage1_36[49], stage1_36[50], stage1_36[51], stage1_36[52], stage1_36[53]},
      {stage1_37[78], stage1_37[79], stage1_37[80]},
      {stage1_38[4]},
      {stage2_39[15],stage2_38[18],stage2_37[26],stage2_36[41]}
   );
   gpc606_5 gpc3235 (
      {stage1_36[54], stage1_36[55], stage1_36[56], stage1_36[57], stage1_36[58], stage1_36[59]},
      {stage1_38[5], stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10]},
      {stage2_40[0],stage2_39[16],stage2_38[19],stage2_37[27],stage2_36[42]}
   );
   gpc606_5 gpc3236 (
      {stage1_36[60], stage1_36[61], stage1_36[62], stage1_36[63], stage1_36[64], stage1_36[65]},
      {stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16]},
      {stage2_40[1],stage2_39[17],stage2_38[20],stage2_37[28],stage2_36[43]}
   );
   gpc606_5 gpc3237 (
      {stage1_36[66], stage1_36[67], stage1_36[68], stage1_36[69], stage1_36[70], stage1_36[71]},
      {stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20], stage1_38[21], stage1_38[22]},
      {stage2_40[2],stage2_39[18],stage2_38[21],stage2_37[29],stage2_36[44]}
   );
   gpc606_5 gpc3238 (
      {stage1_36[72], stage1_36[73], stage1_36[74], stage1_36[75], stage1_36[76], stage1_36[77]},
      {stage1_38[23], stage1_38[24], stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28]},
      {stage2_40[3],stage2_39[19],stage2_38[22],stage2_37[30],stage2_36[45]}
   );
   gpc606_5 gpc3239 (
      {stage1_36[78], stage1_36[79], stage1_36[80], stage1_36[81], stage1_36[82], stage1_36[83]},
      {stage1_38[29], stage1_38[30], stage1_38[31], stage1_38[32], stage1_38[33], stage1_38[34]},
      {stage2_40[4],stage2_39[20],stage2_38[23],stage2_37[31],stage2_36[46]}
   );
   gpc606_5 gpc3240 (
      {stage1_36[84], stage1_36[85], stage1_36[86], stage1_36[87], stage1_36[88], stage1_36[89]},
      {stage1_38[35], stage1_38[36], stage1_38[37], stage1_38[38], stage1_38[39], stage1_38[40]},
      {stage2_40[5],stage2_39[21],stage2_38[24],stage2_37[32],stage2_36[47]}
   );
   gpc606_5 gpc3241 (
      {stage1_36[90], stage1_36[91], stage1_36[92], stage1_36[93], stage1_36[94], stage1_36[95]},
      {stage1_38[41], stage1_38[42], stage1_38[43], stage1_38[44], stage1_38[45], stage1_38[46]},
      {stage2_40[6],stage2_39[22],stage2_38[25],stage2_37[33],stage2_36[48]}
   );
   gpc606_5 gpc3242 (
      {stage1_36[96], stage1_36[97], stage1_36[98], stage1_36[99], stage1_36[100], stage1_36[101]},
      {stage1_38[47], stage1_38[48], stage1_38[49], stage1_38[50], stage1_38[51], stage1_38[52]},
      {stage2_40[7],stage2_39[23],stage2_38[26],stage2_37[34],stage2_36[49]}
   );
   gpc606_5 gpc3243 (
      {stage1_36[102], stage1_36[103], stage1_36[104], stage1_36[105], stage1_36[106], stage1_36[107]},
      {stage1_38[53], stage1_38[54], stage1_38[55], stage1_38[56], stage1_38[57], stage1_38[58]},
      {stage2_40[8],stage2_39[24],stage2_38[27],stage2_37[35],stage2_36[50]}
   );
   gpc606_5 gpc3244 (
      {stage1_36[108], stage1_36[109], stage1_36[110], stage1_36[111], stage1_36[112], stage1_36[113]},
      {stage1_38[59], stage1_38[60], stage1_38[61], stage1_38[62], stage1_38[63], stage1_38[64]},
      {stage2_40[9],stage2_39[25],stage2_38[28],stage2_37[36],stage2_36[51]}
   );
   gpc606_5 gpc3245 (
      {stage1_36[114], stage1_36[115], stage1_36[116], stage1_36[117], stage1_36[118], stage1_36[119]},
      {stage1_38[65], stage1_38[66], stage1_38[67], stage1_38[68], stage1_38[69], stage1_38[70]},
      {stage2_40[10],stage2_39[26],stage2_38[29],stage2_37[37],stage2_36[52]}
   );
   gpc606_5 gpc3246 (
      {stage1_36[120], stage1_36[121], stage1_36[122], stage1_36[123], stage1_36[124], stage1_36[125]},
      {stage1_38[71], stage1_38[72], stage1_38[73], stage1_38[74], stage1_38[75], stage1_38[76]},
      {stage2_40[11],stage2_39[27],stage2_38[30],stage2_37[38],stage2_36[53]}
   );
   gpc606_5 gpc3247 (
      {stage1_36[126], stage1_36[127], stage1_36[128], stage1_36[129], stage1_36[130], stage1_36[131]},
      {stage1_38[77], stage1_38[78], stage1_38[79], stage1_38[80], stage1_38[81], stage1_38[82]},
      {stage2_40[12],stage2_39[28],stage2_38[31],stage2_37[39],stage2_36[54]}
   );
   gpc606_5 gpc3248 (
      {stage1_36[132], stage1_36[133], stage1_36[134], stage1_36[135], stage1_36[136], stage1_36[137]},
      {stage1_38[83], stage1_38[84], stage1_38[85], stage1_38[86], stage1_38[87], stage1_38[88]},
      {stage2_40[13],stage2_39[29],stage2_38[32],stage2_37[40],stage2_36[55]}
   );
   gpc606_5 gpc3249 (
      {stage1_37[81], stage1_37[82], stage1_37[83], stage1_37[84], stage1_37[85], stage1_37[86]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[14],stage2_39[30],stage2_38[33],stage2_37[41]}
   );
   gpc606_5 gpc3250 (
      {stage1_37[87], stage1_37[88], stage1_37[89], stage1_37[90], stage1_37[91], stage1_37[92]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[15],stage2_39[31],stage2_38[34],stage2_37[42]}
   );
   gpc615_5 gpc3251 (
      {stage1_38[89], stage1_38[90], stage1_38[91], stage1_38[92], stage1_38[93]},
      {stage1_39[12]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[2],stage2_40[16],stage2_39[32],stage2_38[35]}
   );
   gpc615_5 gpc3252 (
      {stage1_38[94], stage1_38[95], stage1_38[96], stage1_38[97], stage1_38[98]},
      {stage1_39[13]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[3],stage2_40[17],stage2_39[33],stage2_38[36]}
   );
   gpc615_5 gpc3253 (
      {stage1_38[99], stage1_38[100], stage1_38[101], stage1_38[102], stage1_38[103]},
      {stage1_39[14]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[4],stage2_40[18],stage2_39[34],stage2_38[37]}
   );
   gpc615_5 gpc3254 (
      {stage1_38[104], stage1_38[105], stage1_38[106], stage1_38[107], stage1_38[108]},
      {stage1_39[15]},
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage2_42[3],stage2_41[5],stage2_40[19],stage2_39[35],stage2_38[38]}
   );
   gpc615_5 gpc3255 (
      {stage1_38[109], stage1_38[110], stage1_38[111], stage1_38[112], stage1_38[113]},
      {stage1_39[16]},
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage2_42[4],stage2_41[6],stage2_40[20],stage2_39[36],stage2_38[39]}
   );
   gpc615_5 gpc3256 (
      {stage1_38[114], stage1_38[115], stage1_38[116], stage1_38[117], stage1_38[118]},
      {stage1_39[17]},
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage2_42[5],stage2_41[7],stage2_40[21],stage2_39[37],stage2_38[40]}
   );
   gpc615_5 gpc3257 (
      {stage1_38[119], stage1_38[120], stage1_38[121], stage1_38[122], stage1_38[123]},
      {stage1_39[18]},
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage2_42[6],stage2_41[8],stage2_40[22],stage2_39[38],stage2_38[41]}
   );
   gpc615_5 gpc3258 (
      {stage1_38[124], stage1_38[125], stage1_38[126], stage1_38[127], stage1_38[128]},
      {stage1_39[19]},
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage2_42[7],stage2_41[9],stage2_40[23],stage2_39[39],stage2_38[42]}
   );
   gpc615_5 gpc3259 (
      {stage1_38[129], stage1_38[130], stage1_38[131], stage1_38[132], stage1_38[133]},
      {stage1_39[20]},
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage2_42[8],stage2_41[10],stage2_40[24],stage2_39[40],stage2_38[43]}
   );
   gpc606_5 gpc3260 (
      {stage1_39[21], stage1_39[22], stage1_39[23], stage1_39[24], stage1_39[25], stage1_39[26]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage2_43[0],stage2_42[9],stage2_41[11],stage2_40[25],stage2_39[41]}
   );
   gpc606_5 gpc3261 (
      {stage1_39[27], stage1_39[28], stage1_39[29], stage1_39[30], stage1_39[31], stage1_39[32]},
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage2_43[1],stage2_42[10],stage2_41[12],stage2_40[26],stage2_39[42]}
   );
   gpc606_5 gpc3262 (
      {stage1_39[33], stage1_39[34], stage1_39[35], stage1_39[36], stage1_39[37], stage1_39[38]},
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage2_43[2],stage2_42[11],stage2_41[13],stage2_40[27],stage2_39[43]}
   );
   gpc606_5 gpc3263 (
      {stage1_39[39], stage1_39[40], stage1_39[41], stage1_39[42], stage1_39[43], stage1_39[44]},
      {stage1_41[18], stage1_41[19], stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23]},
      {stage2_43[3],stage2_42[12],stage2_41[14],stage2_40[28],stage2_39[44]}
   );
   gpc606_5 gpc3264 (
      {stage1_39[45], stage1_39[46], stage1_39[47], stage1_39[48], stage1_39[49], stage1_39[50]},
      {stage1_41[24], stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage2_43[4],stage2_42[13],stage2_41[15],stage2_40[29],stage2_39[45]}
   );
   gpc606_5 gpc3265 (
      {stage1_39[51], stage1_39[52], stage1_39[53], stage1_39[54], stage1_39[55], stage1_39[56]},
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34], stage1_41[35]},
      {stage2_43[5],stage2_42[14],stage2_41[16],stage2_40[30],stage2_39[46]}
   );
   gpc606_5 gpc3266 (
      {stage1_39[57], stage1_39[58], stage1_39[59], stage1_39[60], stage1_39[61], stage1_39[62]},
      {stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39], stage1_41[40], stage1_41[41]},
      {stage2_43[6],stage2_42[15],stage2_41[17],stage2_40[31],stage2_39[47]}
   );
   gpc606_5 gpc3267 (
      {stage1_39[63], stage1_39[64], stage1_39[65], stage1_39[66], stage1_39[67], stage1_39[68]},
      {stage1_41[42], stage1_41[43], stage1_41[44], stage1_41[45], stage1_41[46], stage1_41[47]},
      {stage2_43[7],stage2_42[16],stage2_41[18],stage2_40[32],stage2_39[48]}
   );
   gpc606_5 gpc3268 (
      {stage1_39[69], stage1_39[70], stage1_39[71], stage1_39[72], stage1_39[73], stage1_39[74]},
      {stage1_41[48], stage1_41[49], stage1_41[50], stage1_41[51], stage1_41[52], stage1_41[53]},
      {stage2_43[8],stage2_42[17],stage2_41[19],stage2_40[33],stage2_39[49]}
   );
   gpc606_5 gpc3269 (
      {stage1_39[75], stage1_39[76], stage1_39[77], stage1_39[78], stage1_39[79], stage1_39[80]},
      {stage1_41[54], stage1_41[55], stage1_41[56], stage1_41[57], stage1_41[58], stage1_41[59]},
      {stage2_43[9],stage2_42[18],stage2_41[20],stage2_40[34],stage2_39[50]}
   );
   gpc606_5 gpc3270 (
      {stage1_39[81], stage1_39[82], stage1_39[83], stage1_39[84], stage1_39[85], stage1_39[86]},
      {stage1_41[60], stage1_41[61], stage1_41[62], stage1_41[63], stage1_41[64], stage1_41[65]},
      {stage2_43[10],stage2_42[19],stage2_41[21],stage2_40[35],stage2_39[51]}
   );
   gpc606_5 gpc3271 (
      {stage1_39[87], stage1_39[88], stage1_39[89], stage1_39[90], stage1_39[91], stage1_39[92]},
      {stage1_41[66], stage1_41[67], stage1_41[68], stage1_41[69], stage1_41[70], stage1_41[71]},
      {stage2_43[11],stage2_42[20],stage2_41[22],stage2_40[36],stage2_39[52]}
   );
   gpc615_5 gpc3272 (
      {stage1_39[93], stage1_39[94], stage1_39[95], stage1_39[96], stage1_39[97]},
      {stage1_40[54]},
      {stage1_41[72], stage1_41[73], stage1_41[74], stage1_41[75], stage1_41[76], stage1_41[77]},
      {stage2_43[12],stage2_42[21],stage2_41[23],stage2_40[37],stage2_39[53]}
   );
   gpc606_5 gpc3273 (
      {stage1_40[55], stage1_40[56], stage1_40[57], stage1_40[58], stage1_40[59], stage1_40[60]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[13],stage2_42[22],stage2_41[24],stage2_40[38]}
   );
   gpc606_5 gpc3274 (
      {stage1_40[61], stage1_40[62], stage1_40[63], stage1_40[64], stage1_40[65], stage1_40[66]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[14],stage2_42[23],stage2_41[25],stage2_40[39]}
   );
   gpc606_5 gpc3275 (
      {stage1_40[67], stage1_40[68], stage1_40[69], stage1_40[70], stage1_40[71], stage1_40[72]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[15],stage2_42[24],stage2_41[26],stage2_40[40]}
   );
   gpc606_5 gpc3276 (
      {stage1_40[73], stage1_40[74], stage1_40[75], stage1_40[76], stage1_40[77], stage1_40[78]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[16],stage2_42[25],stage2_41[27],stage2_40[41]}
   );
   gpc606_5 gpc3277 (
      {stage1_40[79], stage1_40[80], stage1_40[81], stage1_40[82], stage1_40[83], stage1_40[84]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[17],stage2_42[26],stage2_41[28],stage2_40[42]}
   );
   gpc606_5 gpc3278 (
      {stage1_40[85], stage1_40[86], stage1_40[87], stage1_40[88], stage1_40[89], stage1_40[90]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[18],stage2_42[27],stage2_41[29],stage2_40[43]}
   );
   gpc606_5 gpc3279 (
      {stage1_41[78], stage1_41[79], stage1_41[80], stage1_41[81], stage1_41[82], stage1_41[83]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[6],stage2_43[19],stage2_42[28],stage2_41[30]}
   );
   gpc606_5 gpc3280 (
      {stage1_41[84], stage1_41[85], stage1_41[86], stage1_41[87], stage1_41[88], stage1_41[89]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[7],stage2_43[20],stage2_42[29],stage2_41[31]}
   );
   gpc606_5 gpc3281 (
      {stage1_41[90], stage1_41[91], stage1_41[92], stage1_41[93], stage1_41[94], stage1_41[95]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[8],stage2_43[21],stage2_42[30],stage2_41[32]}
   );
   gpc606_5 gpc3282 (
      {stage1_41[96], stage1_41[97], stage1_41[98], stage1_41[99], stage1_41[100], stage1_41[101]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[9],stage2_43[22],stage2_42[31],stage2_41[33]}
   );
   gpc606_5 gpc3283 (
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage2_46[0],stage2_45[4],stage2_44[10],stage2_43[23],stage2_42[32]}
   );
   gpc606_5 gpc3284 (
      {stage1_42[42], stage1_42[43], stage1_42[44], stage1_42[45], stage1_42[46], stage1_42[47]},
      {stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9], stage1_44[10], stage1_44[11]},
      {stage2_46[1],stage2_45[5],stage2_44[11],stage2_43[24],stage2_42[33]}
   );
   gpc606_5 gpc3285 (
      {stage1_42[48], stage1_42[49], stage1_42[50], stage1_42[51], stage1_42[52], stage1_42[53]},
      {stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16], stage1_44[17]},
      {stage2_46[2],stage2_45[6],stage2_44[12],stage2_43[25],stage2_42[34]}
   );
   gpc606_5 gpc3286 (
      {stage1_42[54], stage1_42[55], stage1_42[56], stage1_42[57], stage1_42[58], stage1_42[59]},
      {stage1_44[18], stage1_44[19], stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23]},
      {stage2_46[3],stage2_45[7],stage2_44[13],stage2_43[26],stage2_42[35]}
   );
   gpc606_5 gpc3287 (
      {stage1_42[60], stage1_42[61], stage1_42[62], stage1_42[63], stage1_42[64], stage1_42[65]},
      {stage1_44[24], stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage2_46[4],stage2_45[8],stage2_44[14],stage2_43[27],stage2_42[36]}
   );
   gpc606_5 gpc3288 (
      {stage1_42[66], stage1_42[67], stage1_42[68], stage1_42[69], stage1_42[70], stage1_42[71]},
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34], stage1_44[35]},
      {stage2_46[5],stage2_45[9],stage2_44[15],stage2_43[28],stage2_42[37]}
   );
   gpc606_5 gpc3289 (
      {stage1_42[72], stage1_42[73], stage1_42[74], stage1_42[75], stage1_42[76], stage1_42[77]},
      {stage1_44[36], stage1_44[37], stage1_44[38], stage1_44[39], stage1_44[40], stage1_44[41]},
      {stage2_46[6],stage2_45[10],stage2_44[16],stage2_43[29],stage2_42[38]}
   );
   gpc606_5 gpc3290 (
      {stage1_42[78], stage1_42[79], stage1_42[80], stage1_42[81], stage1_42[82], stage1_42[83]},
      {stage1_44[42], stage1_44[43], stage1_44[44], stage1_44[45], stage1_44[46], stage1_44[47]},
      {stage2_46[7],stage2_45[11],stage2_44[17],stage2_43[30],stage2_42[39]}
   );
   gpc606_5 gpc3291 (
      {stage1_42[84], stage1_42[85], stage1_42[86], stage1_42[87], stage1_42[88], stage1_42[89]},
      {stage1_44[48], stage1_44[49], stage1_44[50], stage1_44[51], stage1_44[52], stage1_44[53]},
      {stage2_46[8],stage2_45[12],stage2_44[18],stage2_43[31],stage2_42[40]}
   );
   gpc606_5 gpc3292 (
      {stage1_42[90], stage1_42[91], stage1_42[92], stage1_42[93], stage1_42[94], stage1_42[95]},
      {stage1_44[54], stage1_44[55], stage1_44[56], stage1_44[57], stage1_44[58], stage1_44[59]},
      {stage2_46[9],stage2_45[13],stage2_44[19],stage2_43[32],stage2_42[41]}
   );
   gpc606_5 gpc3293 (
      {stage1_42[96], stage1_42[97], stage1_42[98], stage1_42[99], stage1_42[100], stage1_42[101]},
      {stage1_44[60], stage1_44[61], stage1_44[62], stage1_44[63], stage1_44[64], stage1_44[65]},
      {stage2_46[10],stage2_45[14],stage2_44[20],stage2_43[33],stage2_42[42]}
   );
   gpc606_5 gpc3294 (
      {stage1_42[102], stage1_42[103], stage1_42[104], stage1_42[105], stage1_42[106], stage1_42[107]},
      {stage1_44[66], stage1_44[67], stage1_44[68], stage1_44[69], stage1_44[70], stage1_44[71]},
      {stage2_46[11],stage2_45[15],stage2_44[21],stage2_43[34],stage2_42[43]}
   );
   gpc606_5 gpc3295 (
      {stage1_42[108], stage1_42[109], stage1_42[110], stage1_42[111], stage1_42[112], stage1_42[113]},
      {stage1_44[72], stage1_44[73], stage1_44[74], stage1_44[75], stage1_44[76], stage1_44[77]},
      {stage2_46[12],stage2_45[16],stage2_44[22],stage2_43[35],stage2_42[44]}
   );
   gpc606_5 gpc3296 (
      {stage1_42[114], stage1_42[115], stage1_42[116], stage1_42[117], stage1_42[118], stage1_42[119]},
      {stage1_44[78], stage1_44[79], stage1_44[80], stage1_44[81], stage1_44[82], stage1_44[83]},
      {stage2_46[13],stage2_45[17],stage2_44[23],stage2_43[36],stage2_42[45]}
   );
   gpc606_5 gpc3297 (
      {stage1_42[120], stage1_42[121], stage1_42[122], stage1_42[123], stage1_42[124], stage1_42[125]},
      {stage1_44[84], stage1_44[85], stage1_44[86], stage1_44[87], stage1_44[88], stage1_44[89]},
      {stage2_46[14],stage2_45[18],stage2_44[24],stage2_43[37],stage2_42[46]}
   );
   gpc606_5 gpc3298 (
      {stage1_42[126], stage1_42[127], stage1_42[128], stage1_42[129], stage1_42[130], stage1_42[131]},
      {stage1_44[90], stage1_44[91], stage1_44[92], stage1_44[93], stage1_44[94], stage1_44[95]},
      {stage2_46[15],stage2_45[19],stage2_44[25],stage2_43[38],stage2_42[47]}
   );
   gpc606_5 gpc3299 (
      {stage1_42[132], stage1_42[133], stage1_42[134], stage1_42[135], stage1_42[136], stage1_42[137]},
      {stage1_44[96], stage1_44[97], stage1_44[98], stage1_44[99], stage1_44[100], stage1_44[101]},
      {stage2_46[16],stage2_45[20],stage2_44[26],stage2_43[39],stage2_42[48]}
   );
   gpc606_5 gpc3300 (
      {stage1_42[138], stage1_42[139], stage1_42[140], stage1_42[141], stage1_42[142], stage1_42[143]},
      {stage1_44[102], stage1_44[103], stage1_44[104], stage1_44[105], stage1_44[106], stage1_44[107]},
      {stage2_46[17],stage2_45[21],stage2_44[27],stage2_43[40],stage2_42[49]}
   );
   gpc606_5 gpc3301 (
      {stage1_42[144], stage1_42[145], stage1_42[146], stage1_42[147], stage1_42[148], stage1_42[149]},
      {stage1_44[108], stage1_44[109], stage1_44[110], stage1_44[111], stage1_44[112], stage1_44[113]},
      {stage2_46[18],stage2_45[22],stage2_44[28],stage2_43[41],stage2_42[50]}
   );
   gpc606_5 gpc3302 (
      {stage1_42[150], stage1_42[151], stage1_42[152], stage1_42[153], stage1_42[154], stage1_42[155]},
      {stage1_44[114], stage1_44[115], stage1_44[116], stage1_44[117], stage1_44[118], stage1_44[119]},
      {stage2_46[19],stage2_45[23],stage2_44[29],stage2_43[42],stage2_42[51]}
   );
   gpc606_5 gpc3303 (
      {stage1_42[156], stage1_42[157], stage1_42[158], stage1_42[159], stage1_42[160], stage1_42[161]},
      {stage1_44[120], stage1_44[121], stage1_44[122], stage1_44[123], stage1_44[124], stage1_44[125]},
      {stage2_46[20],stage2_45[24],stage2_44[30],stage2_43[43],stage2_42[52]}
   );
   gpc606_5 gpc3304 (
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[21],stage2_45[25],stage2_44[31],stage2_43[44]}
   );
   gpc615_5 gpc3305 (
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34]},
      {stage1_44[126]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[22],stage2_45[26],stage2_44[32],stage2_43[45]}
   );
   gpc615_5 gpc3306 (
      {stage1_43[35], stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39]},
      {stage1_44[127]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[23],stage2_45[27],stage2_44[33],stage2_43[46]}
   );
   gpc615_5 gpc3307 (
      {stage1_43[40], stage1_43[41], stage1_43[42], stage1_43[43], stage1_43[44]},
      {stage1_44[128]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[24],stage2_45[28],stage2_44[34],stage2_43[47]}
   );
   gpc615_5 gpc3308 (
      {stage1_43[45], stage1_43[46], stage1_43[47], stage1_43[48], stage1_43[49]},
      {stage1_44[129]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[25],stage2_45[29],stage2_44[35],stage2_43[48]}
   );
   gpc615_5 gpc3309 (
      {stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53], stage1_43[54]},
      {stage1_44[130]},
      {stage1_45[30], stage1_45[31], stage1_45[32], stage1_45[33], stage1_45[34], stage1_45[35]},
      {stage2_47[5],stage2_46[26],stage2_45[30],stage2_44[36],stage2_43[49]}
   );
   gpc615_5 gpc3310 (
      {stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage1_44[131]},
      {stage1_45[36], stage1_45[37], stage1_45[38], stage1_45[39], stage1_45[40], stage1_45[41]},
      {stage2_47[6],stage2_46[27],stage2_45[31],stage2_44[37],stage2_43[50]}
   );
   gpc615_5 gpc3311 (
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64]},
      {stage1_44[132]},
      {stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46], stage1_45[47]},
      {stage2_47[7],stage2_46[28],stage2_45[32],stage2_44[38],stage2_43[51]}
   );
   gpc615_5 gpc3312 (
      {stage1_43[65], stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69]},
      {stage1_44[133]},
      {stage1_45[48], stage1_45[49], stage1_45[50], stage1_45[51], stage1_45[52], stage1_45[53]},
      {stage2_47[8],stage2_46[29],stage2_45[33],stage2_44[39],stage2_43[52]}
   );
   gpc606_5 gpc3313 (
      {stage1_45[54], stage1_45[55], stage1_45[56], stage1_45[57], stage1_45[58], stage1_45[59]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[0],stage2_47[9],stage2_46[30],stage2_45[34]}
   );
   gpc606_5 gpc3314 (
      {stage1_45[60], stage1_45[61], stage1_45[62], stage1_45[63], stage1_45[64], stage1_45[65]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[1],stage2_47[10],stage2_46[31],stage2_45[35]}
   );
   gpc606_5 gpc3315 (
      {stage1_45[66], stage1_45[67], stage1_45[68], stage1_45[69], stage1_45[70], stage1_45[71]},
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17]},
      {stage2_49[2],stage2_48[2],stage2_47[11],stage2_46[32],stage2_45[36]}
   );
   gpc606_5 gpc3316 (
      {stage1_45[72], stage1_45[73], stage1_45[74], stage1_45[75], stage1_45[76], stage1_45[77]},
      {stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23]},
      {stage2_49[3],stage2_48[3],stage2_47[12],stage2_46[33],stage2_45[37]}
   );
   gpc606_5 gpc3317 (
      {stage1_45[78], stage1_45[79], stage1_45[80], stage1_45[81], stage1_45[82], stage1_45[83]},
      {stage1_47[24], stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29]},
      {stage2_49[4],stage2_48[4],stage2_47[13],stage2_46[34],stage2_45[38]}
   );
   gpc606_5 gpc3318 (
      {stage1_45[84], stage1_45[85], stage1_45[86], stage1_45[87], stage1_45[88], stage1_45[89]},
      {stage1_47[30], stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35]},
      {stage2_49[5],stage2_48[5],stage2_47[14],stage2_46[35],stage2_45[39]}
   );
   gpc606_5 gpc3319 (
      {stage1_45[90], stage1_45[91], stage1_45[92], stage1_45[93], stage1_45[94], stage1_45[95]},
      {stage1_47[36], stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41]},
      {stage2_49[6],stage2_48[6],stage2_47[15],stage2_46[36],stage2_45[40]}
   );
   gpc606_5 gpc3320 (
      {stage1_45[96], stage1_45[97], stage1_45[98], stage1_45[99], stage1_45[100], stage1_45[101]},
      {stage1_47[42], stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47]},
      {stage2_49[7],stage2_48[7],stage2_47[16],stage2_46[37],stage2_45[41]}
   );
   gpc606_5 gpc3321 (
      {stage1_45[102], stage1_45[103], stage1_45[104], stage1_45[105], stage1_45[106], stage1_45[107]},
      {stage1_47[48], stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage2_49[8],stage2_48[8],stage2_47[17],stage2_46[38],stage2_45[42]}
   );
   gpc606_5 gpc3322 (
      {stage1_45[108], stage1_45[109], stage1_45[110], stage1_45[111], stage1_45[112], stage1_45[113]},
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58], stage1_47[59]},
      {stage2_49[9],stage2_48[9],stage2_47[18],stage2_46[39],stage2_45[43]}
   );
   gpc606_5 gpc3323 (
      {stage1_45[114], stage1_45[115], stage1_45[116], stage1_45[117], stage1_45[118], stage1_45[119]},
      {stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63], stage1_47[64], stage1_47[65]},
      {stage2_49[10],stage2_48[10],stage2_47[19],stage2_46[40],stage2_45[44]}
   );
   gpc606_5 gpc3324 (
      {stage1_45[120], stage1_45[121], stage1_45[122], stage1_45[123], stage1_45[124], stage1_45[125]},
      {stage1_47[66], stage1_47[67], stage1_47[68], stage1_47[69], stage1_47[70], stage1_47[71]},
      {stage2_49[11],stage2_48[11],stage2_47[20],stage2_46[41],stage2_45[45]}
   );
   gpc606_5 gpc3325 (
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[12],stage2_48[12],stage2_47[21],stage2_46[42]}
   );
   gpc606_5 gpc3326 (
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[13],stage2_48[13],stage2_47[22],stage2_46[43]}
   );
   gpc606_5 gpc3327 (
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[14],stage2_48[14],stage2_47[23],stage2_46[44]}
   );
   gpc606_5 gpc3328 (
      {stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21], stage1_46[22], stage1_46[23]},
      {stage1_48[18], stage1_48[19], stage1_48[20], stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage2_50[3],stage2_49[15],stage2_48[15],stage2_47[24],stage2_46[45]}
   );
   gpc606_5 gpc3329 (
      {stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27], stage1_46[28], stage1_46[29]},
      {stage1_48[24], stage1_48[25], stage1_48[26], stage1_48[27], stage1_48[28], stage1_48[29]},
      {stage2_50[4],stage2_49[16],stage2_48[16],stage2_47[25],stage2_46[46]}
   );
   gpc606_5 gpc3330 (
      {stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35]},
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage2_50[5],stage2_49[17],stage2_48[17],stage2_47[26],stage2_46[47]}
   );
   gpc606_5 gpc3331 (
      {stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage2_50[6],stage2_49[18],stage2_48[18],stage2_47[27],stage2_46[48]}
   );
   gpc606_5 gpc3332 (
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46], stage1_46[47]},
      {stage1_48[42], stage1_48[43], stage1_48[44], stage1_48[45], stage1_48[46], stage1_48[47]},
      {stage2_50[7],stage2_49[19],stage2_48[19],stage2_47[28],stage2_46[49]}
   );
   gpc606_5 gpc3333 (
      {stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51], stage1_46[52], stage1_46[53]},
      {stage1_48[48], stage1_48[49], stage1_48[50], stage1_48[51], stage1_48[52], stage1_48[53]},
      {stage2_50[8],stage2_49[20],stage2_48[20],stage2_47[29],stage2_46[50]}
   );
   gpc606_5 gpc3334 (
      {stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57], stage1_46[58], stage1_46[59]},
      {stage1_48[54], stage1_48[55], stage1_48[56], stage1_48[57], stage1_48[58], stage1_48[59]},
      {stage2_50[9],stage2_49[21],stage2_48[21],stage2_47[30],stage2_46[51]}
   );
   gpc606_5 gpc3335 (
      {stage1_46[60], stage1_46[61], stage1_46[62], stage1_46[63], stage1_46[64], stage1_46[65]},
      {stage1_48[60], stage1_48[61], stage1_48[62], stage1_48[63], stage1_48[64], stage1_48[65]},
      {stage2_50[10],stage2_49[22],stage2_48[22],stage2_47[31],stage2_46[52]}
   );
   gpc606_5 gpc3336 (
      {stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69], stage1_46[70], stage1_46[71]},
      {stage1_48[66], stage1_48[67], stage1_48[68], stage1_48[69], stage1_48[70], stage1_48[71]},
      {stage2_50[11],stage2_49[23],stage2_48[23],stage2_47[32],stage2_46[53]}
   );
   gpc606_5 gpc3337 (
      {stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75], stage1_46[76], stage1_46[77]},
      {stage1_48[72], stage1_48[73], stage1_48[74], stage1_48[75], stage1_48[76], stage1_48[77]},
      {stage2_50[12],stage2_49[24],stage2_48[24],stage2_47[33],stage2_46[54]}
   );
   gpc606_5 gpc3338 (
      {stage1_46[78], stage1_46[79], stage1_46[80], stage1_46[81], stage1_46[82], stage1_46[83]},
      {stage1_48[78], stage1_48[79], stage1_48[80], stage1_48[81], stage1_48[82], stage1_48[83]},
      {stage2_50[13],stage2_49[25],stage2_48[25],stage2_47[34],stage2_46[55]}
   );
   gpc606_5 gpc3339 (
      {stage1_46[84], stage1_46[85], stage1_46[86], stage1_46[87], stage1_46[88], stage1_46[89]},
      {stage1_48[84], stage1_48[85], stage1_48[86], stage1_48[87], stage1_48[88], stage1_48[89]},
      {stage2_50[14],stage2_49[26],stage2_48[26],stage2_47[35],stage2_46[56]}
   );
   gpc606_5 gpc3340 (
      {stage1_46[90], stage1_46[91], stage1_46[92], stage1_46[93], stage1_46[94], stage1_46[95]},
      {stage1_48[90], stage1_48[91], stage1_48[92], stage1_48[93], stage1_48[94], stage1_48[95]},
      {stage2_50[15],stage2_49[27],stage2_48[27],stage2_47[36],stage2_46[57]}
   );
   gpc606_5 gpc3341 (
      {stage1_47[72], stage1_47[73], stage1_47[74], stage1_47[75], stage1_47[76], stage1_47[77]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[16],stage2_49[28],stage2_48[28],stage2_47[37]}
   );
   gpc606_5 gpc3342 (
      {stage1_47[78], stage1_47[79], stage1_47[80], stage1_47[81], stage1_47[82], stage1_47[83]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[17],stage2_49[29],stage2_48[29],stage2_47[38]}
   );
   gpc606_5 gpc3343 (
      {stage1_47[84], stage1_47[85], stage1_47[86], stage1_47[87], stage1_47[88], stage1_47[89]},
      {stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15], stage1_49[16], stage1_49[17]},
      {stage2_51[2],stage2_50[18],stage2_49[30],stage2_48[30],stage2_47[39]}
   );
   gpc606_5 gpc3344 (
      {stage1_47[90], stage1_47[91], stage1_47[92], stage1_47[93], stage1_47[94], stage1_47[95]},
      {stage1_49[18], stage1_49[19], stage1_49[20], stage1_49[21], stage1_49[22], stage1_49[23]},
      {stage2_51[3],stage2_50[19],stage2_49[31],stage2_48[31],stage2_47[40]}
   );
   gpc623_5 gpc3345 (
      {stage1_47[96], stage1_47[97], stage1_47[98]},
      {stage1_48[96], stage1_48[97]},
      {stage1_49[24], stage1_49[25], stage1_49[26], stage1_49[27], stage1_49[28], stage1_49[29]},
      {stage2_51[4],stage2_50[20],stage2_49[32],stage2_48[32],stage2_47[41]}
   );
   gpc623_5 gpc3346 (
      {stage1_47[99], stage1_47[100], stage1_47[101]},
      {stage1_48[98], stage1_48[99]},
      {stage1_49[30], stage1_49[31], stage1_49[32], stage1_49[33], stage1_49[34], stage1_49[35]},
      {stage2_51[5],stage2_50[21],stage2_49[33],stage2_48[33],stage2_47[42]}
   );
   gpc1406_5 gpc3347 (
      {stage1_49[36], stage1_49[37], stage1_49[38], stage1_49[39], stage1_49[40], stage1_49[41]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3]},
      {stage1_52[0]},
      {stage2_53[0],stage2_52[0],stage2_51[6],stage2_50[22],stage2_49[34]}
   );
   gpc606_5 gpc3348 (
      {stage1_49[42], stage1_49[43], stage1_49[44], stage1_49[45], stage1_49[46], stage1_49[47]},
      {stage1_51[4], stage1_51[5], stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9]},
      {stage2_53[1],stage2_52[1],stage2_51[7],stage2_50[23],stage2_49[35]}
   );
   gpc606_5 gpc3349 (
      {stage1_49[48], stage1_49[49], stage1_49[50], stage1_49[51], stage1_49[52], stage1_49[53]},
      {stage1_51[10], stage1_51[11], stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15]},
      {stage2_53[2],stage2_52[2],stage2_51[8],stage2_50[24],stage2_49[36]}
   );
   gpc606_5 gpc3350 (
      {stage1_49[54], stage1_49[55], stage1_49[56], stage1_49[57], stage1_49[58], stage1_49[59]},
      {stage1_51[16], stage1_51[17], stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21]},
      {stage2_53[3],stage2_52[3],stage2_51[9],stage2_50[25],stage2_49[37]}
   );
   gpc606_5 gpc3351 (
      {stage1_49[60], stage1_49[61], stage1_49[62], stage1_49[63], stage1_49[64], stage1_49[65]},
      {stage1_51[22], stage1_51[23], stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27]},
      {stage2_53[4],stage2_52[4],stage2_51[10],stage2_50[26],stage2_49[38]}
   );
   gpc606_5 gpc3352 (
      {stage1_49[66], stage1_49[67], stage1_49[68], stage1_49[69], stage1_49[70], stage1_49[71]},
      {stage1_51[28], stage1_51[29], stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33]},
      {stage2_53[5],stage2_52[5],stage2_51[11],stage2_50[27],stage2_49[39]}
   );
   gpc606_5 gpc3353 (
      {stage1_49[72], stage1_49[73], stage1_49[74], stage1_49[75], stage1_49[76], stage1_49[77]},
      {stage1_51[34], stage1_51[35], stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39]},
      {stage2_53[6],stage2_52[6],stage2_51[12],stage2_50[28],stage2_49[40]}
   );
   gpc615_5 gpc3354 (
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4]},
      {stage1_51[40]},
      {stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5], stage1_52[6]},
      {stage2_54[0],stage2_53[7],stage2_52[7],stage2_51[13],stage2_50[29]}
   );
   gpc615_5 gpc3355 (
      {stage1_50[5], stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9]},
      {stage1_51[41]},
      {stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11], stage1_52[12]},
      {stage2_54[1],stage2_53[8],stage2_52[8],stage2_51[14],stage2_50[30]}
   );
   gpc615_5 gpc3356 (
      {stage1_50[10], stage1_50[11], stage1_50[12], stage1_50[13], stage1_50[14]},
      {stage1_51[42]},
      {stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17], stage1_52[18]},
      {stage2_54[2],stage2_53[9],stage2_52[9],stage2_51[15],stage2_50[31]}
   );
   gpc615_5 gpc3357 (
      {stage1_50[15], stage1_50[16], stage1_50[17], stage1_50[18], stage1_50[19]},
      {stage1_51[43]},
      {stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23], stage1_52[24]},
      {stage2_54[3],stage2_53[10],stage2_52[10],stage2_51[16],stage2_50[32]}
   );
   gpc615_5 gpc3358 (
      {stage1_50[20], stage1_50[21], stage1_50[22], stage1_50[23], stage1_50[24]},
      {stage1_51[44]},
      {stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28], stage1_52[29], stage1_52[30]},
      {stage2_54[4],stage2_53[11],stage2_52[11],stage2_51[17],stage2_50[33]}
   );
   gpc615_5 gpc3359 (
      {stage1_50[25], stage1_50[26], stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage1_51[45]},
      {stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34], stage1_52[35], stage1_52[36]},
      {stage2_54[5],stage2_53[12],stage2_52[12],stage2_51[18],stage2_50[34]}
   );
   gpc615_5 gpc3360 (
      {stage1_50[30], stage1_50[31], stage1_50[32], stage1_50[33], stage1_50[34]},
      {stage1_51[46]},
      {stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41], stage1_52[42]},
      {stage2_54[6],stage2_53[13],stage2_52[13],stage2_51[19],stage2_50[35]}
   );
   gpc615_5 gpc3361 (
      {stage1_50[35], stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39]},
      {stage1_51[47]},
      {stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47], stage1_52[48]},
      {stage2_54[7],stage2_53[14],stage2_52[14],stage2_51[20],stage2_50[36]}
   );
   gpc615_5 gpc3362 (
      {stage1_50[40], stage1_50[41], stage1_50[42], stage1_50[43], stage1_50[44]},
      {stage1_51[48]},
      {stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53], stage1_52[54]},
      {stage2_54[8],stage2_53[15],stage2_52[15],stage2_51[21],stage2_50[37]}
   );
   gpc615_5 gpc3363 (
      {stage1_50[45], stage1_50[46], stage1_50[47], stage1_50[48], stage1_50[49]},
      {stage1_51[49]},
      {stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59], stage1_52[60]},
      {stage2_54[9],stage2_53[16],stage2_52[16],stage2_51[22],stage2_50[38]}
   );
   gpc615_5 gpc3364 (
      {stage1_50[50], stage1_50[51], stage1_50[52], stage1_50[53], stage1_50[54]},
      {stage1_51[50]},
      {stage1_52[61], stage1_52[62], stage1_52[63], stage1_52[64], stage1_52[65], stage1_52[66]},
      {stage2_54[10],stage2_53[17],stage2_52[17],stage2_51[23],stage2_50[39]}
   );
   gpc615_5 gpc3365 (
      {stage1_50[55], stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59]},
      {stage1_51[51]},
      {stage1_52[67], stage1_52[68], stage1_52[69], stage1_52[70], stage1_52[71], stage1_52[72]},
      {stage2_54[11],stage2_53[18],stage2_52[18],stage2_51[24],stage2_50[40]}
   );
   gpc615_5 gpc3366 (
      {stage1_50[60], stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64]},
      {stage1_51[52]},
      {stage1_52[73], stage1_52[74], stage1_52[75], stage1_52[76], stage1_52[77], stage1_52[78]},
      {stage2_54[12],stage2_53[19],stage2_52[19],stage2_51[25],stage2_50[41]}
   );
   gpc615_5 gpc3367 (
      {stage1_50[65], stage1_50[66], stage1_50[67], stage1_50[68], stage1_50[69]},
      {stage1_51[53]},
      {stage1_52[79], stage1_52[80], stage1_52[81], stage1_52[82], stage1_52[83], stage1_52[84]},
      {stage2_54[13],stage2_53[20],stage2_52[20],stage2_51[26],stage2_50[42]}
   );
   gpc615_5 gpc3368 (
      {stage1_50[70], stage1_50[71], stage1_50[72], stage1_50[73], stage1_50[74]},
      {stage1_51[54]},
      {stage1_52[85], stage1_52[86], stage1_52[87], stage1_52[88], stage1_52[89], stage1_52[90]},
      {stage2_54[14],stage2_53[21],stage2_52[21],stage2_51[27],stage2_50[43]}
   );
   gpc615_5 gpc3369 (
      {stage1_52[91], stage1_52[92], stage1_52[93], stage1_52[94], stage1_52[95]},
      {stage1_53[0]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[0],stage2_54[15],stage2_53[22],stage2_52[22]}
   );
   gpc615_5 gpc3370 (
      {stage1_52[96], stage1_52[97], stage1_52[98], stage1_52[99], stage1_52[100]},
      {stage1_53[1]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[1],stage2_54[16],stage2_53[23],stage2_52[23]}
   );
   gpc615_5 gpc3371 (
      {stage1_52[101], stage1_52[102], stage1_52[103], stage1_52[104], stage1_52[105]},
      {stage1_53[2]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[2],stage2_54[17],stage2_53[24],stage2_52[24]}
   );
   gpc615_5 gpc3372 (
      {stage1_52[106], stage1_52[107], stage1_52[108], stage1_52[109], stage1_52[110]},
      {stage1_53[3]},
      {stage1_54[18], stage1_54[19], stage1_54[20], stage1_54[21], stage1_54[22], stage1_54[23]},
      {stage2_56[3],stage2_55[3],stage2_54[18],stage2_53[25],stage2_52[25]}
   );
   gpc615_5 gpc3373 (
      {stage1_52[111], stage1_52[112], stage1_52[113], stage1_52[114], stage1_52[115]},
      {stage1_53[4]},
      {stage1_54[24], stage1_54[25], stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29]},
      {stage2_56[4],stage2_55[4],stage2_54[19],stage2_53[26],stage2_52[26]}
   );
   gpc615_5 gpc3374 (
      {stage1_53[5], stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9]},
      {stage1_54[30]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[5],stage2_55[5],stage2_54[20],stage2_53[27]}
   );
   gpc615_5 gpc3375 (
      {stage1_53[10], stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14]},
      {stage1_54[31]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[6],stage2_55[6],stage2_54[21],stage2_53[28]}
   );
   gpc615_5 gpc3376 (
      {stage1_53[15], stage1_53[16], stage1_53[17], stage1_53[18], stage1_53[19]},
      {stage1_54[32]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[7],stage2_55[7],stage2_54[22],stage2_53[29]}
   );
   gpc615_5 gpc3377 (
      {stage1_53[20], stage1_53[21], stage1_53[22], stage1_53[23], stage1_53[24]},
      {stage1_54[33]},
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23]},
      {stage2_57[3],stage2_56[8],stage2_55[8],stage2_54[23],stage2_53[30]}
   );
   gpc615_5 gpc3378 (
      {stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage1_54[34]},
      {stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29]},
      {stage2_57[4],stage2_56[9],stage2_55[9],stage2_54[24],stage2_53[31]}
   );
   gpc615_5 gpc3379 (
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34]},
      {stage1_54[35]},
      {stage1_55[30], stage1_55[31], stage1_55[32], stage1_55[33], stage1_55[34], stage1_55[35]},
      {stage2_57[5],stage2_56[10],stage2_55[10],stage2_54[25],stage2_53[32]}
   );
   gpc615_5 gpc3380 (
      {stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39]},
      {stage1_54[36]},
      {stage1_55[36], stage1_55[37], stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41]},
      {stage2_57[6],stage2_56[11],stage2_55[11],stage2_54[26],stage2_53[33]}
   );
   gpc615_5 gpc3381 (
      {stage1_53[40], stage1_53[41], stage1_53[42], stage1_53[43], stage1_53[44]},
      {stage1_54[37]},
      {stage1_55[42], stage1_55[43], stage1_55[44], stage1_55[45], stage1_55[46], stage1_55[47]},
      {stage2_57[7],stage2_56[12],stage2_55[12],stage2_54[27],stage2_53[34]}
   );
   gpc615_5 gpc3382 (
      {stage1_53[45], stage1_53[46], stage1_53[47], stage1_53[48], stage1_53[49]},
      {stage1_54[38]},
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52], stage1_55[53]},
      {stage2_57[8],stage2_56[13],stage2_55[13],stage2_54[28],stage2_53[35]}
   );
   gpc615_5 gpc3383 (
      {stage1_53[50], stage1_53[51], stage1_53[52], stage1_53[53], stage1_53[54]},
      {stage1_54[39]},
      {stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57], stage1_55[58], stage1_55[59]},
      {stage2_57[9],stage2_56[14],stage2_55[14],stage2_54[29],stage2_53[36]}
   );
   gpc615_5 gpc3384 (
      {stage1_53[55], stage1_53[56], stage1_53[57], stage1_53[58], stage1_53[59]},
      {stage1_54[40]},
      {stage1_55[60], stage1_55[61], stage1_55[62], stage1_55[63], stage1_55[64], stage1_55[65]},
      {stage2_57[10],stage2_56[15],stage2_55[15],stage2_54[30],stage2_53[37]}
   );
   gpc615_5 gpc3385 (
      {stage1_53[60], stage1_53[61], stage1_53[62], stage1_53[63], stage1_53[64]},
      {stage1_54[41]},
      {stage1_55[66], stage1_55[67], stage1_55[68], stage1_55[69], stage1_55[70], stage1_55[71]},
      {stage2_57[11],stage2_56[16],stage2_55[16],stage2_54[31],stage2_53[38]}
   );
   gpc615_5 gpc3386 (
      {stage1_53[65], stage1_53[66], stage1_53[67], stage1_53[68], stage1_53[69]},
      {stage1_54[42]},
      {stage1_55[72], stage1_55[73], stage1_55[74], stage1_55[75], stage1_55[76], stage1_55[77]},
      {stage2_57[12],stage2_56[17],stage2_55[17],stage2_54[32],stage2_53[39]}
   );
   gpc606_5 gpc3387 (
      {stage1_54[43], stage1_54[44], stage1_54[45], stage1_54[46], stage1_54[47], stage1_54[48]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[13],stage2_56[18],stage2_55[18],stage2_54[33]}
   );
   gpc606_5 gpc3388 (
      {stage1_54[49], stage1_54[50], stage1_54[51], stage1_54[52], stage1_54[53], stage1_54[54]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[14],stage2_56[19],stage2_55[19],stage2_54[34]}
   );
   gpc606_5 gpc3389 (
      {stage1_54[55], stage1_54[56], stage1_54[57], stage1_54[58], stage1_54[59], stage1_54[60]},
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage2_58[2],stage2_57[15],stage2_56[20],stage2_55[20],stage2_54[35]}
   );
   gpc606_5 gpc3390 (
      {stage1_54[61], stage1_54[62], stage1_54[63], stage1_54[64], stage1_54[65], stage1_54[66]},
      {stage1_56[18], stage1_56[19], stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage2_58[3],stage2_57[16],stage2_56[21],stage2_55[21],stage2_54[36]}
   );
   gpc606_5 gpc3391 (
      {stage1_54[67], stage1_54[68], stage1_54[69], stage1_54[70], stage1_54[71], stage1_54[72]},
      {stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage2_58[4],stage2_57[17],stage2_56[22],stage2_55[22],stage2_54[37]}
   );
   gpc606_5 gpc3392 (
      {stage1_54[73], stage1_54[74], stage1_54[75], stage1_54[76], stage1_54[77], stage1_54[78]},
      {stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage2_58[5],stage2_57[18],stage2_56[23],stage2_55[23],stage2_54[38]}
   );
   gpc606_5 gpc3393 (
      {stage1_54[79], stage1_54[80], stage1_54[81], stage1_54[82], stage1_54[83], stage1_54[84]},
      {stage1_56[36], stage1_56[37], stage1_56[38], stage1_56[39], stage1_56[40], stage1_56[41]},
      {stage2_58[6],stage2_57[19],stage2_56[24],stage2_55[24],stage2_54[39]}
   );
   gpc606_5 gpc3394 (
      {stage1_54[85], stage1_54[86], stage1_54[87], stage1_54[88], stage1_54[89], stage1_54[90]},
      {stage1_56[42], stage1_56[43], stage1_56[44], stage1_56[45], stage1_56[46], stage1_56[47]},
      {stage2_58[7],stage2_57[20],stage2_56[25],stage2_55[25],stage2_54[40]}
   );
   gpc606_5 gpc3395 (
      {stage1_54[91], stage1_54[92], stage1_54[93], stage1_54[94], stage1_54[95], stage1_54[96]},
      {stage1_56[48], stage1_56[49], stage1_56[50], stage1_56[51], stage1_56[52], stage1_56[53]},
      {stage2_58[8],stage2_57[21],stage2_56[26],stage2_55[26],stage2_54[41]}
   );
   gpc606_5 gpc3396 (
      {stage1_54[97], stage1_54[98], stage1_54[99], stage1_54[100], stage1_54[101], stage1_54[102]},
      {stage1_56[54], stage1_56[55], stage1_56[56], stage1_56[57], stage1_56[58], stage1_56[59]},
      {stage2_58[9],stage2_57[22],stage2_56[27],stage2_55[27],stage2_54[42]}
   );
   gpc606_5 gpc3397 (
      {stage1_54[103], stage1_54[104], stage1_54[105], stage1_54[106], stage1_54[107], stage1_54[108]},
      {stage1_56[60], stage1_56[61], stage1_56[62], stage1_56[63], stage1_56[64], stage1_56[65]},
      {stage2_58[10],stage2_57[23],stage2_56[28],stage2_55[28],stage2_54[43]}
   );
   gpc606_5 gpc3398 (
      {stage1_54[109], stage1_54[110], stage1_54[111], stage1_54[112], stage1_54[113], stage1_54[114]},
      {stage1_56[66], stage1_56[67], stage1_56[68], stage1_56[69], stage1_56[70], stage1_56[71]},
      {stage2_58[11],stage2_57[24],stage2_56[29],stage2_55[29],stage2_54[44]}
   );
   gpc606_5 gpc3399 (
      {stage1_54[115], stage1_54[116], stage1_54[117], stage1_54[118], stage1_54[119], stage1_54[120]},
      {stage1_56[72], stage1_56[73], stage1_56[74], stage1_56[75], stage1_56[76], stage1_56[77]},
      {stage2_58[12],stage2_57[25],stage2_56[30],stage2_55[30],stage2_54[45]}
   );
   gpc606_5 gpc3400 (
      {stage1_54[121], stage1_54[122], stage1_54[123], stage1_54[124], stage1_54[125], stage1_54[126]},
      {stage1_56[78], stage1_56[79], stage1_56[80], stage1_56[81], stage1_56[82], stage1_56[83]},
      {stage2_58[13],stage2_57[26],stage2_56[31],stage2_55[31],stage2_54[46]}
   );
   gpc606_5 gpc3401 (
      {stage1_54[127], stage1_54[128], stage1_54[129], stage1_54[130], stage1_54[131], stage1_54[132]},
      {stage1_56[84], stage1_56[85], stage1_56[86], stage1_56[87], stage1_56[88], stage1_56[89]},
      {stage2_58[14],stage2_57[27],stage2_56[32],stage2_55[32],stage2_54[47]}
   );
   gpc606_5 gpc3402 (
      {stage1_55[78], stage1_55[79], stage1_55[80], stage1_55[81], stage1_55[82], stage1_55[83]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[15],stage2_57[28],stage2_56[33],stage2_55[33]}
   );
   gpc606_5 gpc3403 (
      {stage1_55[84], stage1_55[85], stage1_55[86], stage1_55[87], stage1_55[88], stage1_55[89]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[16],stage2_57[29],stage2_56[34],stage2_55[34]}
   );
   gpc606_5 gpc3404 (
      {stage1_56[90], stage1_56[91], stage1_56[92], stage1_56[93], stage1_56[94], stage1_56[95]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[2],stage2_58[17],stage2_57[30],stage2_56[35]}
   );
   gpc606_5 gpc3405 (
      {stage1_56[96], stage1_56[97], stage1_56[98], stage1_56[99], stage1_56[100], stage1_56[101]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[3],stage2_58[18],stage2_57[31],stage2_56[36]}
   );
   gpc606_5 gpc3406 (
      {stage1_56[102], stage1_56[103], stage1_56[104], stage1_56[105], stage1_56[106], stage1_56[107]},
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage2_60[2],stage2_59[4],stage2_58[19],stage2_57[32],stage2_56[37]}
   );
   gpc606_5 gpc3407 (
      {stage1_56[108], stage1_56[109], stage1_56[110], stage1_56[111], stage1_56[112], stage1_56[113]},
      {stage1_58[18], stage1_58[19], stage1_58[20], stage1_58[21], stage1_58[22], stage1_58[23]},
      {stage2_60[3],stage2_59[5],stage2_58[20],stage2_57[33],stage2_56[38]}
   );
   gpc606_5 gpc3408 (
      {stage1_56[114], stage1_56[115], stage1_56[116], stage1_56[117], stage1_56[118], stage1_56[119]},
      {stage1_58[24], stage1_58[25], stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29]},
      {stage2_60[4],stage2_59[6],stage2_58[21],stage2_57[34],stage2_56[39]}
   );
   gpc606_5 gpc3409 (
      {stage1_56[120], stage1_56[121], stage1_56[122], stage1_56[123], stage1_56[124], stage1_56[125]},
      {stage1_58[30], stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage2_60[5],stage2_59[7],stage2_58[22],stage2_57[35],stage2_56[40]}
   );
   gpc606_5 gpc3410 (
      {stage1_56[126], stage1_56[127], stage1_56[128], stage1_56[129], stage1_56[130], stage1_56[131]},
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage2_60[6],stage2_59[8],stage2_58[23],stage2_57[36],stage2_56[41]}
   );
   gpc606_5 gpc3411 (
      {stage1_56[132], stage1_56[133], stage1_56[134], stage1_56[135], stage1_56[136], stage1_56[137]},
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage2_60[7],stage2_59[9],stage2_58[24],stage2_57[37],stage2_56[42]}
   );
   gpc606_5 gpc3412 (
      {stage1_56[138], stage1_56[139], stage1_56[140], stage1_56[141], stage1_56[142], stage1_56[143]},
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage2_60[8],stage2_59[10],stage2_58[25],stage2_57[38],stage2_56[43]}
   );
   gpc606_5 gpc3413 (
      {stage1_56[144], stage1_56[145], stage1_56[146], stage1_56[147], stage1_56[148], stage1_56[149]},
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage2_60[9],stage2_59[11],stage2_58[26],stage2_57[39],stage2_56[44]}
   );
   gpc606_5 gpc3414 (
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[10],stage2_59[12],stage2_58[27],stage2_57[40]}
   );
   gpc606_5 gpc3415 (
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[11],stage2_59[13],stage2_58[28],stage2_57[41]}
   );
   gpc606_5 gpc3416 (
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[12],stage2_59[14],stage2_58[29],stage2_57[42]}
   );
   gpc606_5 gpc3417 (
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[13],stage2_59[15],stage2_58[30],stage2_57[43]}
   );
   gpc606_5 gpc3418 (
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage1_59[24], stage1_59[25], stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29]},
      {stage2_61[4],stage2_60[14],stage2_59[16],stage2_58[31],stage2_57[44]}
   );
   gpc606_5 gpc3419 (
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage1_59[30], stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], stage1_59[35]},
      {stage2_61[5],stage2_60[15],stage2_59[17],stage2_58[32],stage2_57[45]}
   );
   gpc606_5 gpc3420 (
      {stage1_57[48], stage1_57[49], stage1_57[50], stage1_57[51], stage1_57[52], stage1_57[53]},
      {stage1_59[36], stage1_59[37], stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41]},
      {stage2_61[6],stage2_60[16],stage2_59[18],stage2_58[33],stage2_57[46]}
   );
   gpc606_5 gpc3421 (
      {stage1_57[54], stage1_57[55], stage1_57[56], stage1_57[57], stage1_57[58], stage1_57[59]},
      {stage1_59[42], stage1_59[43], stage1_59[44], stage1_59[45], stage1_59[46], stage1_59[47]},
      {stage2_61[7],stage2_60[17],stage2_59[19],stage2_58[34],stage2_57[47]}
   );
   gpc606_5 gpc3422 (
      {stage1_57[60], stage1_57[61], stage1_57[62], stage1_57[63], stage1_57[64], stage1_57[65]},
      {stage1_59[48], stage1_59[49], stage1_59[50], stage1_59[51], stage1_59[52], stage1_59[53]},
      {stage2_61[8],stage2_60[18],stage2_59[20],stage2_58[35],stage2_57[48]}
   );
   gpc606_5 gpc3423 (
      {stage1_57[66], stage1_57[67], stage1_57[68], stage1_57[69], stage1_57[70], stage1_57[71]},
      {stage1_59[54], stage1_59[55], stage1_59[56], stage1_59[57], stage1_59[58], stage1_59[59]},
      {stage2_61[9],stage2_60[19],stage2_59[21],stage2_58[36],stage2_57[49]}
   );
   gpc606_5 gpc3424 (
      {stage1_58[60], stage1_58[61], stage1_58[62], stage1_58[63], stage1_58[64], stage1_58[65]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[10],stage2_60[20],stage2_59[22],stage2_58[37]}
   );
   gpc606_5 gpc3425 (
      {stage1_58[66], stage1_58[67], stage1_58[68], stage1_58[69], stage1_58[70], stage1_58[71]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[11],stage2_60[21],stage2_59[23],stage2_58[38]}
   );
   gpc606_5 gpc3426 (
      {stage1_58[72], stage1_58[73], stage1_58[74], stage1_58[75], stage1_58[76], stage1_58[77]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[12],stage2_60[22],stage2_59[24],stage2_58[39]}
   );
   gpc606_5 gpc3427 (
      {stage1_59[60], stage1_59[61], stage1_59[62], stage1_59[63], stage1_59[64], stage1_59[65]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[3],stage2_61[13],stage2_60[23],stage2_59[25]}
   );
   gpc606_5 gpc3428 (
      {stage1_59[66], stage1_59[67], stage1_59[68], stage1_59[69], stage1_59[70], stage1_59[71]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[4],stage2_61[14],stage2_60[24],stage2_59[26]}
   );
   gpc606_5 gpc3429 (
      {stage1_59[72], stage1_59[73], stage1_59[74], stage1_59[75], stage1_59[76], stage1_59[77]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[5],stage2_61[15],stage2_60[25],stage2_59[27]}
   );
   gpc606_5 gpc3430 (
      {stage1_59[78], stage1_59[79], stage1_59[80], stage1_59[81], stage1_59[82], stage1_59[83]},
      {stage1_61[18], stage1_61[19], stage1_61[20], stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage2_63[3],stage2_62[6],stage2_61[16],stage2_60[26],stage2_59[28]}
   );
   gpc606_5 gpc3431 (
      {stage1_59[84], stage1_59[85], stage1_59[86], stage1_59[87], stage1_59[88], stage1_59[89]},
      {stage1_61[24], stage1_61[25], stage1_61[26], stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage2_63[4],stage2_62[7],stage2_61[17],stage2_60[27],stage2_59[29]}
   );
   gpc606_5 gpc3432 (
      {stage1_59[90], stage1_59[91], stage1_59[92], stage1_59[93], stage1_59[94], stage1_59[95]},
      {stage1_61[30], stage1_61[31], stage1_61[32], stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage2_63[5],stage2_62[8],stage2_61[18],stage2_60[28],stage2_59[30]}
   );
   gpc606_5 gpc3433 (
      {stage1_59[96], stage1_59[97], stage1_59[98], stage1_59[99], stage1_59[100], stage1_59[101]},
      {stage1_61[36], stage1_61[37], stage1_61[38], stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage2_63[6],stage2_62[9],stage2_61[19],stage2_60[29],stage2_59[31]}
   );
   gpc606_5 gpc3434 (
      {stage1_59[102], stage1_59[103], stage1_59[104], stage1_59[105], stage1_59[106], stage1_59[107]},
      {stage1_61[42], stage1_61[43], stage1_61[44], stage1_61[45], stage1_61[46], stage1_61[47]},
      {stage2_63[7],stage2_62[10],stage2_61[20],stage2_60[30],stage2_59[32]}
   );
   gpc606_5 gpc3435 (
      {stage1_59[108], stage1_59[109], stage1_59[110], stage1_59[111], stage1_59[112], stage1_59[113]},
      {stage1_61[48], stage1_61[49], stage1_61[50], stage1_61[51], stage1_61[52], stage1_61[53]},
      {stage2_63[8],stage2_62[11],stage2_61[21],stage2_60[31],stage2_59[33]}
   );
   gpc606_5 gpc3436 (
      {stage1_59[114], stage1_59[115], stage1_59[116], stage1_59[117], stage1_59[118], stage1_59[119]},
      {stage1_61[54], stage1_61[55], stage1_61[56], stage1_61[57], stage1_61[58], stage1_61[59]},
      {stage2_63[9],stage2_62[12],stage2_61[22],stage2_60[32],stage2_59[34]}
   );
   gpc606_5 gpc3437 (
      {stage1_59[120], stage1_59[121], stage1_59[122], stage1_59[123], stage1_59[124], stage1_59[125]},
      {stage1_61[60], stage1_61[61], stage1_61[62], stage1_61[63], stage1_61[64], stage1_61[65]},
      {stage2_63[10],stage2_62[13],stage2_61[23],stage2_60[33],stage2_59[35]}
   );
   gpc606_5 gpc3438 (
      {stage1_59[126], stage1_59[127], stage1_59[128], stage1_59[129], stage1_59[130], stage1_59[131]},
      {stage1_61[66], stage1_61[67], stage1_61[68], stage1_61[69], stage1_61[70], stage1_61[71]},
      {stage2_63[11],stage2_62[14],stage2_61[24],stage2_60[34],stage2_59[36]}
   );
   gpc606_5 gpc3439 (
      {stage1_59[132], stage1_59[133], stage1_59[134], stage1_59[135], stage1_59[136], stage1_59[137]},
      {stage1_61[72], stage1_61[73], stage1_61[74], stage1_61[75], stage1_61[76], stage1_61[77]},
      {stage2_63[12],stage2_62[15],stage2_61[25],stage2_60[35],stage2_59[37]}
   );
   gpc606_5 gpc3440 (
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[13],stage2_62[16],stage2_61[26],stage2_60[36]}
   );
   gpc606_5 gpc3441 (
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage2_64[1],stage2_63[14],stage2_62[17],stage2_61[27],stage2_60[37]}
   );
   gpc606_5 gpc3442 (
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage2_64[2],stage2_63[15],stage2_62[18],stage2_61[28],stage2_60[38]}
   );
   gpc606_5 gpc3443 (
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage2_64[3],stage2_63[16],stage2_62[19],stage2_61[29],stage2_60[39]}
   );
   gpc606_5 gpc3444 (
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage2_64[4],stage2_63[17],stage2_62[20],stage2_61[30],stage2_60[40]}
   );
   gpc615_5 gpc3445 (
      {stage1_60[48], stage1_60[49], stage1_60[50], stage1_60[51], stage1_60[52]},
      {stage1_61[78]},
      {stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35]},
      {stage2_64[5],stage2_63[18],stage2_62[21],stage2_61[31],stage2_60[41]}
   );
   gpc615_5 gpc3446 (
      {stage1_60[53], stage1_60[54], stage1_60[55], stage1_60[56], stage1_60[57]},
      {stage1_61[79]},
      {stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39], stage1_62[40], stage1_62[41]},
      {stage2_64[6],stage2_63[19],stage2_62[22],stage2_61[32],stage2_60[42]}
   );
   gpc615_5 gpc3447 (
      {stage1_60[58], stage1_60[59], stage1_60[60], stage1_60[61], stage1_60[62]},
      {stage1_61[80]},
      {stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45], stage1_62[46], stage1_62[47]},
      {stage2_64[7],stage2_63[20],stage2_62[23],stage2_61[33],stage2_60[43]}
   );
   gpc615_5 gpc3448 (
      {stage1_60[63], stage1_60[64], stage1_60[65], stage1_60[66], stage1_60[67]},
      {stage1_61[81]},
      {stage1_62[48], stage1_62[49], stage1_62[50], stage1_62[51], stage1_62[52], stage1_62[53]},
      {stage2_64[8],stage2_63[21],stage2_62[24],stage2_61[34],stage2_60[44]}
   );
   gpc615_5 gpc3449 (
      {stage1_60[68], stage1_60[69], stage1_60[70], stage1_60[71], stage1_60[72]},
      {stage1_61[82]},
      {stage1_62[54], stage1_62[55], stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59]},
      {stage2_64[9],stage2_63[22],stage2_62[25],stage2_61[35],stage2_60[45]}
   );
   gpc615_5 gpc3450 (
      {stage1_60[73], stage1_60[74], stage1_60[75], stage1_60[76], stage1_60[77]},
      {stage1_61[83]},
      {stage1_62[60], stage1_62[61], stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65]},
      {stage2_64[10],stage2_63[23],stage2_62[26],stage2_61[36],stage2_60[46]}
   );
   gpc615_5 gpc3451 (
      {stage1_60[78], stage1_60[79], stage1_60[80], stage1_60[81], stage1_60[82]},
      {stage1_61[84]},
      {stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69], stage1_62[70], stage1_62[71]},
      {stage2_64[11],stage2_63[24],stage2_62[27],stage2_61[37],stage2_60[47]}
   );
   gpc615_5 gpc3452 (
      {stage1_60[83], stage1_60[84], stage1_60[85], stage1_60[86], stage1_60[87]},
      {stage1_61[85]},
      {stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75], stage1_62[76], stage1_62[77]},
      {stage2_64[12],stage2_63[25],stage2_62[28],stage2_61[38],stage2_60[48]}
   );
   gpc615_5 gpc3453 (
      {stage1_60[88], stage1_60[89], stage1_60[90], stage1_60[91], stage1_60[92]},
      {stage1_61[86]},
      {stage1_62[78], stage1_62[79], stage1_62[80], stage1_62[81], stage1_62[82], stage1_62[83]},
      {stage2_64[13],stage2_63[26],stage2_62[29],stage2_61[39],stage2_60[49]}
   );
   gpc615_5 gpc3454 (
      {stage1_60[93], stage1_60[94], stage1_60[95], stage1_60[96], stage1_60[97]},
      {stage1_61[87]},
      {stage1_62[84], stage1_62[85], stage1_62[86], stage1_62[87], stage1_62[88], stage1_62[89]},
      {stage2_64[14],stage2_63[27],stage2_62[30],stage2_61[40],stage2_60[50]}
   );
   gpc615_5 gpc3455 (
      {stage1_60[98], stage1_60[99], stage1_60[100], stage1_60[101], stage1_60[102]},
      {stage1_61[88]},
      {stage1_62[90], stage1_62[91], stage1_62[92], stage1_62[93], stage1_62[94], stage1_62[95]},
      {stage2_64[15],stage2_63[28],stage2_62[31],stage2_61[41],stage2_60[51]}
   );
   gpc615_5 gpc3456 (
      {stage1_60[103], stage1_60[104], stage1_60[105], stage1_60[106], stage1_60[107]},
      {stage1_61[89]},
      {stage1_62[96], stage1_62[97], stage1_62[98], stage1_62[99], stage1_62[100], stage1_62[101]},
      {stage2_64[16],stage2_63[29],stage2_62[32],stage2_61[42],stage2_60[52]}
   );
   gpc615_5 gpc3457 (
      {stage1_60[108], stage1_60[109], stage1_60[110], stage1_60[111], stage1_60[112]},
      {stage1_61[90]},
      {stage1_62[102], stage1_62[103], stage1_62[104], stage1_62[105], stage1_62[106], stage1_62[107]},
      {stage2_64[17],stage2_63[30],stage2_62[33],stage2_61[43],stage2_60[53]}
   );
   gpc615_5 gpc3458 (
      {stage1_60[113], stage1_60[114], stage1_60[115], stage1_60[116], stage1_60[117]},
      {stage1_61[91]},
      {stage1_62[108], stage1_62[109], stage1_62[110], stage1_62[111], stage1_62[112], stage1_62[113]},
      {stage2_64[18],stage2_63[31],stage2_62[34],stage2_61[44],stage2_60[54]}
   );
   gpc615_5 gpc3459 (
      {stage1_60[118], stage1_60[119], stage1_60[120], stage1_60[121], stage1_60[122]},
      {stage1_61[92]},
      {stage1_62[114], stage1_62[115], stage1_62[116], stage1_62[117], stage1_62[118], stage1_62[119]},
      {stage2_64[19],stage2_63[32],stage2_62[35],stage2_61[45],stage2_60[55]}
   );
   gpc615_5 gpc3460 (
      {stage1_60[123], stage1_60[124], stage1_60[125], stage1_60[126], stage1_60[127]},
      {stage1_61[93]},
      {stage1_62[120], stage1_62[121], stage1_62[122], stage1_62[123], stage1_62[124], stage1_62[125]},
      {stage2_64[20],stage2_63[33],stage2_62[36],stage2_61[46],stage2_60[56]}
   );
   gpc615_5 gpc3461 (
      {stage1_60[128], stage1_60[129], stage1_60[130], stage1_60[131], stage1_60[132]},
      {stage1_61[94]},
      {stage1_62[126], stage1_62[127], stage1_62[128], stage1_62[129], stage1_62[130], stage1_62[131]},
      {stage2_64[21],stage2_63[34],stage2_62[37],stage2_61[47],stage2_60[57]}
   );
   gpc615_5 gpc3462 (
      {stage1_60[133], stage1_60[134], stage1_60[135], stage1_60[136], stage1_60[137]},
      {stage1_61[95]},
      {stage1_62[132], stage1_62[133], stage1_62[134], stage1_62[135], stage1_62[136], stage1_62[137]},
      {stage2_64[22],stage2_63[35],stage2_62[38],stage2_61[48],stage2_60[58]}
   );
   gpc606_5 gpc3463 (
      {stage1_61[96], stage1_61[97], stage1_61[98], stage1_61[99], stage1_61[100], stage1_61[101]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[23],stage2_63[36],stage2_62[39],stage2_61[49]}
   );
   gpc606_5 gpc3464 (
      {stage1_62[138], stage1_62[139], stage1_62[140], stage1_62[141], stage1_62[142], stage1_62[143]},
      {stage1_64[0], stage1_64[1], stage1_64[2], stage1_64[3], stage1_64[4], stage1_64[5]},
      {stage2_66[0],stage2_65[1],stage2_64[24],stage2_63[37],stage2_62[40]}
   );
   gpc606_5 gpc3465 (
      {stage1_62[144], stage1_62[145], stage1_62[146], stage1_62[147], stage1_62[148], stage1_62[149]},
      {stage1_64[6], stage1_64[7], stage1_64[8], stage1_64[9], stage1_64[10], stage1_64[11]},
      {stage2_66[1],stage2_65[2],stage2_64[25],stage2_63[38],stage2_62[41]}
   );
   gpc606_5 gpc3466 (
      {stage1_62[150], stage1_62[151], stage1_62[152], stage1_62[153], stage1_62[154], stage1_62[155]},
      {stage1_64[12], stage1_64[13], stage1_64[14], stage1_64[15], stage1_64[16], stage1_64[17]},
      {stage2_66[2],stage2_65[3],stage2_64[26],stage2_63[39],stage2_62[42]}
   );
   gpc606_5 gpc3467 (
      {stage1_62[156], stage1_62[157], stage1_62[158], stage1_62[159], stage1_62[160], stage1_62[161]},
      {stage1_64[18], stage1_64[19], stage1_64[20], stage1_64[21], stage1_64[22], stage1_64[23]},
      {stage2_66[3],stage2_65[4],stage2_64[27],stage2_63[40],stage2_62[43]}
   );
   gpc606_5 gpc3468 (
      {stage1_62[162], stage1_62[163], stage1_62[164], stage1_62[165], stage1_62[166], stage1_62[167]},
      {stage1_64[24], stage1_64[25], stage1_64[26], stage1_64[27], stage1_64[28], stage1_64[29]},
      {stage2_66[4],stage2_65[5],stage2_64[28],stage2_63[41],stage2_62[44]}
   );
   gpc606_5 gpc3469 (
      {stage1_62[168], stage1_62[169], stage1_62[170], stage1_62[171], stage1_62[172], stage1_62[173]},
      {stage1_64[30], stage1_64[31], stage1_64[32], stage1_64[33], stage1_64[34], stage1_64[35]},
      {stage2_66[5],stage2_65[6],stage2_64[29],stage2_63[42],stage2_62[45]}
   );
   gpc606_5 gpc3470 (
      {stage1_62[174], stage1_62[175], stage1_62[176], stage1_62[177], stage1_62[178], stage1_62[179]},
      {stage1_64[36], stage1_64[37], stage1_64[38], stage1_64[39], stage1_64[40], stage1_64[41]},
      {stage2_66[6],stage2_65[7],stage2_64[30],stage2_63[43],stage2_62[46]}
   );
   gpc606_5 gpc3471 (
      {stage1_62[180], stage1_62[181], stage1_62[182], stage1_62[183], stage1_62[184], stage1_62[185]},
      {stage1_64[42], stage1_64[43], stage1_64[44], stage1_64[45], stage1_64[46], stage1_64[47]},
      {stage2_66[7],stage2_65[8],stage2_64[31],stage2_63[44],stage2_62[47]}
   );
   gpc606_5 gpc3472 (
      {stage1_62[186], stage1_62[187], stage1_62[188], stage1_62[189], stage1_62[190], stage1_62[191]},
      {stage1_64[48], stage1_64[49], stage1_64[50], stage1_64[51], stage1_64[52], stage1_64[53]},
      {stage2_66[8],stage2_65[9],stage2_64[32],stage2_63[45],stage2_62[48]}
   );
   gpc606_5 gpc3473 (
      {stage1_62[192], stage1_62[193], stage1_62[194], stage1_62[195], stage1_62[196], stage1_62[197]},
      {stage1_64[54], stage1_64[55], stage1_64[56], stage1_64[57], stage1_64[58], stage1_64[59]},
      {stage2_66[9],stage2_65[10],stage2_64[33],stage2_63[46],stage2_62[49]}
   );
   gpc606_5 gpc3474 (
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage1_65[0], stage1_65[1], stage1_65[2], stage1_65[3], stage1_65[4], stage1_65[5]},
      {stage2_67[0],stage2_66[10],stage2_65[11],stage2_64[34],stage2_63[47]}
   );
   gpc606_5 gpc3475 (
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage1_65[6], stage1_65[7], stage1_65[8], stage1_65[9], stage1_65[10], stage1_65[11]},
      {stage2_67[1],stage2_66[11],stage2_65[12],stage2_64[35],stage2_63[48]}
   );
   gpc606_5 gpc3476 (
      {stage1_63[18], stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage1_65[12], stage1_65[13], stage1_65[14], stage1_65[15], stage1_65[16], stage1_65[17]},
      {stage2_67[2],stage2_66[12],stage2_65[13],stage2_64[36],stage2_63[49]}
   );
   gpc606_5 gpc3477 (
      {stage1_63[24], stage1_63[25], stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29]},
      {stage1_65[18], stage1_65[19], stage1_65[20], stage1_65[21], stage1_65[22], stage1_65[23]},
      {stage2_67[3],stage2_66[13],stage2_65[14],stage2_64[37],stage2_63[50]}
   );
   gpc606_5 gpc3478 (
      {stage1_63[30], stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage1_65[24], stage1_65[25], stage1_65[26], stage1_65[27], stage1_65[28], stage1_65[29]},
      {stage2_67[4],stage2_66[14],stage2_65[15],stage2_64[38],stage2_63[51]}
   );
   gpc606_5 gpc3479 (
      {stage1_63[36], stage1_63[37], stage1_63[38], stage1_63[39], stage1_63[40], stage1_63[41]},
      {stage1_65[30], stage1_65[31], stage1_65[32], stage1_65[33], stage1_65[34], stage1_65[35]},
      {stage2_67[5],stage2_66[15],stage2_65[16],stage2_64[39],stage2_63[52]}
   );
   gpc606_5 gpc3480 (
      {stage1_63[42], stage1_63[43], stage1_63[44], stage1_63[45], stage1_63[46], stage1_63[47]},
      {stage1_65[36], stage1_65[37], stage1_65[38], stage1_65[39], stage1_65[40], stage1_65[41]},
      {stage2_67[6],stage2_66[16],stage2_65[17],stage2_64[40],stage2_63[53]}
   );
   gpc1_1 gpc3481 (
      {stage1_0[74]},
      {stage2_0[13]}
   );
   gpc1_1 gpc3482 (
      {stage1_0[75]},
      {stage2_0[14]}
   );
   gpc1_1 gpc3483 (
      {stage1_0[76]},
      {stage2_0[15]}
   );
   gpc1_1 gpc3484 (
      {stage1_0[77]},
      {stage2_0[16]}
   );
   gpc1_1 gpc3485 (
      {stage1_0[78]},
      {stage2_0[17]}
   );
   gpc1_1 gpc3486 (
      {stage1_0[79]},
      {stage2_0[18]}
   );
   gpc1_1 gpc3487 (
      {stage1_0[80]},
      {stage2_0[19]}
   );
   gpc1_1 gpc3488 (
      {stage1_0[81]},
      {stage2_0[20]}
   );
   gpc1_1 gpc3489 (
      {stage1_0[82]},
      {stage2_0[21]}
   );
   gpc1_1 gpc3490 (
      {stage1_0[83]},
      {stage2_0[22]}
   );
   gpc1_1 gpc3491 (
      {stage1_0[84]},
      {stage2_0[23]}
   );
   gpc1_1 gpc3492 (
      {stage1_0[85]},
      {stage2_0[24]}
   );
   gpc1_1 gpc3493 (
      {stage1_0[86]},
      {stage2_0[25]}
   );
   gpc1_1 gpc3494 (
      {stage1_0[87]},
      {stage2_0[26]}
   );
   gpc1_1 gpc3495 (
      {stage1_0[88]},
      {stage2_0[27]}
   );
   gpc1_1 gpc3496 (
      {stage1_0[89]},
      {stage2_0[28]}
   );
   gpc1_1 gpc3497 (
      {stage1_0[90]},
      {stage2_0[29]}
   );
   gpc1_1 gpc3498 (
      {stage1_1[69]},
      {stage2_1[23]}
   );
   gpc1_1 gpc3499 (
      {stage1_1[70]},
      {stage2_1[24]}
   );
   gpc1_1 gpc3500 (
      {stage1_1[71]},
      {stage2_1[25]}
   );
   gpc1_1 gpc3501 (
      {stage1_1[72]},
      {stage2_1[26]}
   );
   gpc1_1 gpc3502 (
      {stage1_1[73]},
      {stage2_1[27]}
   );
   gpc1_1 gpc3503 (
      {stage1_1[74]},
      {stage2_1[28]}
   );
   gpc1_1 gpc3504 (
      {stage1_1[75]},
      {stage2_1[29]}
   );
   gpc1_1 gpc3505 (
      {stage1_1[76]},
      {stage2_1[30]}
   );
   gpc1_1 gpc3506 (
      {stage1_1[77]},
      {stage2_1[31]}
   );
   gpc1_1 gpc3507 (
      {stage1_1[78]},
      {stage2_1[32]}
   );
   gpc1_1 gpc3508 (
      {stage1_1[79]},
      {stage2_1[33]}
   );
   gpc1_1 gpc3509 (
      {stage1_1[80]},
      {stage2_1[34]}
   );
   gpc1_1 gpc3510 (
      {stage1_1[81]},
      {stage2_1[35]}
   );
   gpc1_1 gpc3511 (
      {stage1_1[82]},
      {stage2_1[36]}
   );
   gpc1_1 gpc3512 (
      {stage1_3[92]},
      {stage2_3[39]}
   );
   gpc1_1 gpc3513 (
      {stage1_3[93]},
      {stage2_3[40]}
   );
   gpc1_1 gpc3514 (
      {stage1_3[94]},
      {stage2_3[41]}
   );
   gpc1_1 gpc3515 (
      {stage1_3[95]},
      {stage2_3[42]}
   );
   gpc1_1 gpc3516 (
      {stage1_3[96]},
      {stage2_3[43]}
   );
   gpc1_1 gpc3517 (
      {stage1_3[97]},
      {stage2_3[44]}
   );
   gpc1_1 gpc3518 (
      {stage1_3[98]},
      {stage2_3[45]}
   );
   gpc1_1 gpc3519 (
      {stage1_3[99]},
      {stage2_3[46]}
   );
   gpc1_1 gpc3520 (
      {stage1_3[100]},
      {stage2_3[47]}
   );
   gpc1_1 gpc3521 (
      {stage1_3[101]},
      {stage2_3[48]}
   );
   gpc1_1 gpc3522 (
      {stage1_3[102]},
      {stage2_3[49]}
   );
   gpc1_1 gpc3523 (
      {stage1_3[103]},
      {stage2_3[50]}
   );
   gpc1_1 gpc3524 (
      {stage1_3[104]},
      {stage2_3[51]}
   );
   gpc1_1 gpc3525 (
      {stage1_3[105]},
      {stage2_3[52]}
   );
   gpc1_1 gpc3526 (
      {stage1_3[106]},
      {stage2_3[53]}
   );
   gpc1_1 gpc3527 (
      {stage1_7[106]},
      {stage2_7[39]}
   );
   gpc1_1 gpc3528 (
      {stage1_7[107]},
      {stage2_7[40]}
   );
   gpc1_1 gpc3529 (
      {stage1_7[108]},
      {stage2_7[41]}
   );
   gpc1_1 gpc3530 (
      {stage1_7[109]},
      {stage2_7[42]}
   );
   gpc1_1 gpc3531 (
      {stage1_10[147]},
      {stage2_10[61]}
   );
   gpc1_1 gpc3532 (
      {stage1_10[148]},
      {stage2_10[62]}
   );
   gpc1_1 gpc3533 (
      {stage1_10[149]},
      {stage2_10[63]}
   );
   gpc1_1 gpc3534 (
      {stage1_10[150]},
      {stage2_10[64]}
   );
   gpc1_1 gpc3535 (
      {stage1_10[151]},
      {stage2_10[65]}
   );
   gpc1_1 gpc3536 (
      {stage1_10[152]},
      {stage2_10[66]}
   );
   gpc1_1 gpc3537 (
      {stage1_10[153]},
      {stage2_10[67]}
   );
   gpc1_1 gpc3538 (
      {stage1_10[154]},
      {stage2_10[68]}
   );
   gpc1_1 gpc3539 (
      {stage1_10[155]},
      {stage2_10[69]}
   );
   gpc1_1 gpc3540 (
      {stage1_11[152]},
      {stage2_11[47]}
   );
   gpc1_1 gpc3541 (
      {stage1_11[153]},
      {stage2_11[48]}
   );
   gpc1_1 gpc3542 (
      {stage1_12[132]},
      {stage2_12[53]}
   );
   gpc1_1 gpc3543 (
      {stage1_13[94]},
      {stage2_13[61]}
   );
   gpc1_1 gpc3544 (
      {stage1_13[95]},
      {stage2_13[62]}
   );
   gpc1_1 gpc3545 (
      {stage1_13[96]},
      {stage2_13[63]}
   );
   gpc1_1 gpc3546 (
      {stage1_15[89]},
      {stage2_15[31]}
   );
   gpc1_1 gpc3547 (
      {stage1_15[90]},
      {stage2_15[32]}
   );
   gpc1_1 gpc3548 (
      {stage1_15[91]},
      {stage2_15[33]}
   );
   gpc1_1 gpc3549 (
      {stage1_15[92]},
      {stage2_15[34]}
   );
   gpc1_1 gpc3550 (
      {stage1_15[93]},
      {stage2_15[35]}
   );
   gpc1_1 gpc3551 (
      {stage1_15[94]},
      {stage2_15[36]}
   );
   gpc1_1 gpc3552 (
      {stage1_15[95]},
      {stage2_15[37]}
   );
   gpc1_1 gpc3553 (
      {stage1_15[96]},
      {stage2_15[38]}
   );
   gpc1_1 gpc3554 (
      {stage1_15[97]},
      {stage2_15[39]}
   );
   gpc1_1 gpc3555 (
      {stage1_15[98]},
      {stage2_15[40]}
   );
   gpc1_1 gpc3556 (
      {stage1_15[99]},
      {stage2_15[41]}
   );
   gpc1_1 gpc3557 (
      {stage1_15[100]},
      {stage2_15[42]}
   );
   gpc1_1 gpc3558 (
      {stage1_15[101]},
      {stage2_15[43]}
   );
   gpc1_1 gpc3559 (
      {stage1_15[102]},
      {stage2_15[44]}
   );
   gpc1_1 gpc3560 (
      {stage1_15[103]},
      {stage2_15[45]}
   );
   gpc1_1 gpc3561 (
      {stage1_15[104]},
      {stage2_15[46]}
   );
   gpc1_1 gpc3562 (
      {stage1_15[105]},
      {stage2_15[47]}
   );
   gpc1_1 gpc3563 (
      {stage1_15[106]},
      {stage2_15[48]}
   );
   gpc1_1 gpc3564 (
      {stage1_15[107]},
      {stage2_15[49]}
   );
   gpc1_1 gpc3565 (
      {stage1_15[108]},
      {stage2_15[50]}
   );
   gpc1_1 gpc3566 (
      {stage1_15[109]},
      {stage2_15[51]}
   );
   gpc1_1 gpc3567 (
      {stage1_15[110]},
      {stage2_15[52]}
   );
   gpc1_1 gpc3568 (
      {stage1_15[111]},
      {stage2_15[53]}
   );
   gpc1_1 gpc3569 (
      {stage1_15[112]},
      {stage2_15[54]}
   );
   gpc1_1 gpc3570 (
      {stage1_15[113]},
      {stage2_15[55]}
   );
   gpc1_1 gpc3571 (
      {stage1_15[114]},
      {stage2_15[56]}
   );
   gpc1_1 gpc3572 (
      {stage1_15[115]},
      {stage2_15[57]}
   );
   gpc1_1 gpc3573 (
      {stage1_15[116]},
      {stage2_15[58]}
   );
   gpc1_1 gpc3574 (
      {stage1_15[117]},
      {stage2_15[59]}
   );
   gpc1_1 gpc3575 (
      {stage1_15[118]},
      {stage2_15[60]}
   );
   gpc1_1 gpc3576 (
      {stage1_15[119]},
      {stage2_15[61]}
   );
   gpc1_1 gpc3577 (
      {stage1_15[120]},
      {stage2_15[62]}
   );
   gpc1_1 gpc3578 (
      {stage1_15[121]},
      {stage2_15[63]}
   );
   gpc1_1 gpc3579 (
      {stage1_15[122]},
      {stage2_15[64]}
   );
   gpc1_1 gpc3580 (
      {stage1_15[123]},
      {stage2_15[65]}
   );
   gpc1_1 gpc3581 (
      {stage1_15[124]},
      {stage2_15[66]}
   );
   gpc1_1 gpc3582 (
      {stage1_15[125]},
      {stage2_15[67]}
   );
   gpc1_1 gpc3583 (
      {stage1_15[126]},
      {stage2_15[68]}
   );
   gpc1_1 gpc3584 (
      {stage1_15[127]},
      {stage2_15[69]}
   );
   gpc1_1 gpc3585 (
      {stage1_15[128]},
      {stage2_15[70]}
   );
   gpc1_1 gpc3586 (
      {stage1_15[129]},
      {stage2_15[71]}
   );
   gpc1_1 gpc3587 (
      {stage1_15[130]},
      {stage2_15[72]}
   );
   gpc1_1 gpc3588 (
      {stage1_15[131]},
      {stage2_15[73]}
   );
   gpc1_1 gpc3589 (
      {stage1_16[104]},
      {stage2_16[39]}
   );
   gpc1_1 gpc3590 (
      {stage1_16[105]},
      {stage2_16[40]}
   );
   gpc1_1 gpc3591 (
      {stage1_16[106]},
      {stage2_16[41]}
   );
   gpc1_1 gpc3592 (
      {stage1_16[107]},
      {stage2_16[42]}
   );
   gpc1_1 gpc3593 (
      {stage1_16[108]},
      {stage2_16[43]}
   );
   gpc1_1 gpc3594 (
      {stage1_16[109]},
      {stage2_16[44]}
   );
   gpc1_1 gpc3595 (
      {stage1_16[110]},
      {stage2_16[45]}
   );
   gpc1_1 gpc3596 (
      {stage1_16[111]},
      {stage2_16[46]}
   );
   gpc1_1 gpc3597 (
      {stage1_16[112]},
      {stage2_16[47]}
   );
   gpc1_1 gpc3598 (
      {stage1_16[113]},
      {stage2_16[48]}
   );
   gpc1_1 gpc3599 (
      {stage1_16[114]},
      {stage2_16[49]}
   );
   gpc1_1 gpc3600 (
      {stage1_16[115]},
      {stage2_16[50]}
   );
   gpc1_1 gpc3601 (
      {stage1_16[116]},
      {stage2_16[51]}
   );
   gpc1_1 gpc3602 (
      {stage1_16[117]},
      {stage2_16[52]}
   );
   gpc1_1 gpc3603 (
      {stage1_16[118]},
      {stage2_16[53]}
   );
   gpc1_1 gpc3604 (
      {stage1_16[119]},
      {stage2_16[54]}
   );
   gpc1_1 gpc3605 (
      {stage1_17[102]},
      {stage2_17[48]}
   );
   gpc1_1 gpc3606 (
      {stage1_17[103]},
      {stage2_17[49]}
   );
   gpc1_1 gpc3607 (
      {stage1_17[104]},
      {stage2_17[50]}
   );
   gpc1_1 gpc3608 (
      {stage1_17[105]},
      {stage2_17[51]}
   );
   gpc1_1 gpc3609 (
      {stage1_17[106]},
      {stage2_17[52]}
   );
   gpc1_1 gpc3610 (
      {stage1_17[107]},
      {stage2_17[53]}
   );
   gpc1_1 gpc3611 (
      {stage1_17[108]},
      {stage2_17[54]}
   );
   gpc1_1 gpc3612 (
      {stage1_17[109]},
      {stage2_17[55]}
   );
   gpc1_1 gpc3613 (
      {stage1_17[110]},
      {stage2_17[56]}
   );
   gpc1_1 gpc3614 (
      {stage1_18[71]},
      {stage2_18[37]}
   );
   gpc1_1 gpc3615 (
      {stage1_18[72]},
      {stage2_18[38]}
   );
   gpc1_1 gpc3616 (
      {stage1_18[73]},
      {stage2_18[39]}
   );
   gpc1_1 gpc3617 (
      {stage1_18[74]},
      {stage2_18[40]}
   );
   gpc1_1 gpc3618 (
      {stage1_18[75]},
      {stage2_18[41]}
   );
   gpc1_1 gpc3619 (
      {stage1_18[76]},
      {stage2_18[42]}
   );
   gpc1_1 gpc3620 (
      {stage1_18[77]},
      {stage2_18[43]}
   );
   gpc1_1 gpc3621 (
      {stage1_18[78]},
      {stage2_18[44]}
   );
   gpc1_1 gpc3622 (
      {stage1_18[79]},
      {stage2_18[45]}
   );
   gpc1_1 gpc3623 (
      {stage1_18[80]},
      {stage2_18[46]}
   );
   gpc1_1 gpc3624 (
      {stage1_18[81]},
      {stage2_18[47]}
   );
   gpc1_1 gpc3625 (
      {stage1_18[82]},
      {stage2_18[48]}
   );
   gpc1_1 gpc3626 (
      {stage1_18[83]},
      {stage2_18[49]}
   );
   gpc1_1 gpc3627 (
      {stage1_18[84]},
      {stage2_18[50]}
   );
   gpc1_1 gpc3628 (
      {stage1_18[85]},
      {stage2_18[51]}
   );
   gpc1_1 gpc3629 (
      {stage1_18[86]},
      {stage2_18[52]}
   );
   gpc1_1 gpc3630 (
      {stage1_18[87]},
      {stage2_18[53]}
   );
   gpc1_1 gpc3631 (
      {stage1_18[88]},
      {stage2_18[54]}
   );
   gpc1_1 gpc3632 (
      {stage1_18[89]},
      {stage2_18[55]}
   );
   gpc1_1 gpc3633 (
      {stage1_18[90]},
      {stage2_18[56]}
   );
   gpc1_1 gpc3634 (
      {stage1_18[91]},
      {stage2_18[57]}
   );
   gpc1_1 gpc3635 (
      {stage1_18[92]},
      {stage2_18[58]}
   );
   gpc1_1 gpc3636 (
      {stage1_18[93]},
      {stage2_18[59]}
   );
   gpc1_1 gpc3637 (
      {stage1_18[94]},
      {stage2_18[60]}
   );
   gpc1_1 gpc3638 (
      {stage1_18[95]},
      {stage2_18[61]}
   );
   gpc1_1 gpc3639 (
      {stage1_18[96]},
      {stage2_18[62]}
   );
   gpc1_1 gpc3640 (
      {stage1_18[97]},
      {stage2_18[63]}
   );
   gpc1_1 gpc3641 (
      {stage1_18[98]},
      {stage2_18[64]}
   );
   gpc1_1 gpc3642 (
      {stage1_18[99]},
      {stage2_18[65]}
   );
   gpc1_1 gpc3643 (
      {stage1_19[124]},
      {stage2_19[35]}
   );
   gpc1_1 gpc3644 (
      {stage1_19[125]},
      {stage2_19[36]}
   );
   gpc1_1 gpc3645 (
      {stage1_20[95]},
      {stage2_20[45]}
   );
   gpc1_1 gpc3646 (
      {stage1_20[96]},
      {stage2_20[46]}
   );
   gpc1_1 gpc3647 (
      {stage1_20[97]},
      {stage2_20[47]}
   );
   gpc1_1 gpc3648 (
      {stage1_20[98]},
      {stage2_20[48]}
   );
   gpc1_1 gpc3649 (
      {stage1_20[99]},
      {stage2_20[49]}
   );
   gpc1_1 gpc3650 (
      {stage1_20[100]},
      {stage2_20[50]}
   );
   gpc1_1 gpc3651 (
      {stage1_20[101]},
      {stage2_20[51]}
   );
   gpc1_1 gpc3652 (
      {stage1_20[102]},
      {stage2_20[52]}
   );
   gpc1_1 gpc3653 (
      {stage1_20[103]},
      {stage2_20[53]}
   );
   gpc1_1 gpc3654 (
      {stage1_20[104]},
      {stage2_20[54]}
   );
   gpc1_1 gpc3655 (
      {stage1_20[105]},
      {stage2_20[55]}
   );
   gpc1_1 gpc3656 (
      {stage1_20[106]},
      {stage2_20[56]}
   );
   gpc1_1 gpc3657 (
      {stage1_20[107]},
      {stage2_20[57]}
   );
   gpc1_1 gpc3658 (
      {stage1_20[108]},
      {stage2_20[58]}
   );
   gpc1_1 gpc3659 (
      {stage1_20[109]},
      {stage2_20[59]}
   );
   gpc1_1 gpc3660 (
      {stage1_20[110]},
      {stage2_20[60]}
   );
   gpc1_1 gpc3661 (
      {stage1_20[111]},
      {stage2_20[61]}
   );
   gpc1_1 gpc3662 (
      {stage1_20[112]},
      {stage2_20[62]}
   );
   gpc1_1 gpc3663 (
      {stage1_20[113]},
      {stage2_20[63]}
   );
   gpc1_1 gpc3664 (
      {stage1_20[114]},
      {stage2_20[64]}
   );
   gpc1_1 gpc3665 (
      {stage1_20[115]},
      {stage2_20[65]}
   );
   gpc1_1 gpc3666 (
      {stage1_20[116]},
      {stage2_20[66]}
   );
   gpc1_1 gpc3667 (
      {stage1_20[117]},
      {stage2_20[67]}
   );
   gpc1_1 gpc3668 (
      {stage1_20[118]},
      {stage2_20[68]}
   );
   gpc1_1 gpc3669 (
      {stage1_20[119]},
      {stage2_20[69]}
   );
   gpc1_1 gpc3670 (
      {stage1_20[120]},
      {stage2_20[70]}
   );
   gpc1_1 gpc3671 (
      {stage1_20[121]},
      {stage2_20[71]}
   );
   gpc1_1 gpc3672 (
      {stage1_20[122]},
      {stage2_20[72]}
   );
   gpc1_1 gpc3673 (
      {stage1_20[123]},
      {stage2_20[73]}
   );
   gpc1_1 gpc3674 (
      {stage1_20[124]},
      {stage2_20[74]}
   );
   gpc1_1 gpc3675 (
      {stage1_20[125]},
      {stage2_20[75]}
   );
   gpc1_1 gpc3676 (
      {stage1_20[126]},
      {stage2_20[76]}
   );
   gpc1_1 gpc3677 (
      {stage1_20[127]},
      {stage2_20[77]}
   );
   gpc1_1 gpc3678 (
      {stage1_20[128]},
      {stage2_20[78]}
   );
   gpc1_1 gpc3679 (
      {stage1_20[129]},
      {stage2_20[79]}
   );
   gpc1_1 gpc3680 (
      {stage1_22[87]},
      {stage2_22[36]}
   );
   gpc1_1 gpc3681 (
      {stage1_22[88]},
      {stage2_22[37]}
   );
   gpc1_1 gpc3682 (
      {stage1_22[89]},
      {stage2_22[38]}
   );
   gpc1_1 gpc3683 (
      {stage1_22[90]},
      {stage2_22[39]}
   );
   gpc1_1 gpc3684 (
      {stage1_22[91]},
      {stage2_22[40]}
   );
   gpc1_1 gpc3685 (
      {stage1_23[106]},
      {stage2_23[38]}
   );
   gpc1_1 gpc3686 (
      {stage1_23[107]},
      {stage2_23[39]}
   );
   gpc1_1 gpc3687 (
      {stage1_23[108]},
      {stage2_23[40]}
   );
   gpc1_1 gpc3688 (
      {stage1_23[109]},
      {stage2_23[41]}
   );
   gpc1_1 gpc3689 (
      {stage1_23[110]},
      {stage2_23[42]}
   );
   gpc1_1 gpc3690 (
      {stage1_23[111]},
      {stage2_23[43]}
   );
   gpc1_1 gpc3691 (
      {stage1_23[112]},
      {stage2_23[44]}
   );
   gpc1_1 gpc3692 (
      {stage1_23[113]},
      {stage2_23[45]}
   );
   gpc1_1 gpc3693 (
      {stage1_23[114]},
      {stage2_23[46]}
   );
   gpc1_1 gpc3694 (
      {stage1_23[115]},
      {stage2_23[47]}
   );
   gpc1_1 gpc3695 (
      {stage1_23[116]},
      {stage2_23[48]}
   );
   gpc1_1 gpc3696 (
      {stage1_23[117]},
      {stage2_23[49]}
   );
   gpc1_1 gpc3697 (
      {stage1_23[118]},
      {stage2_23[50]}
   );
   gpc1_1 gpc3698 (
      {stage1_23[119]},
      {stage2_23[51]}
   );
   gpc1_1 gpc3699 (
      {stage1_23[120]},
      {stage2_23[52]}
   );
   gpc1_1 gpc3700 (
      {stage1_23[121]},
      {stage2_23[53]}
   );
   gpc1_1 gpc3701 (
      {stage1_23[122]},
      {stage2_23[54]}
   );
   gpc1_1 gpc3702 (
      {stage1_23[123]},
      {stage2_23[55]}
   );
   gpc1_1 gpc3703 (
      {stage1_23[124]},
      {stage2_23[56]}
   );
   gpc1_1 gpc3704 (
      {stage1_23[125]},
      {stage2_23[57]}
   );
   gpc1_1 gpc3705 (
      {stage1_23[126]},
      {stage2_23[58]}
   );
   gpc1_1 gpc3706 (
      {stage1_23[127]},
      {stage2_23[59]}
   );
   gpc1_1 gpc3707 (
      {stage1_23[128]},
      {stage2_23[60]}
   );
   gpc1_1 gpc3708 (
      {stage1_24[110]},
      {stage2_24[52]}
   );
   gpc1_1 gpc3709 (
      {stage1_24[111]},
      {stage2_24[53]}
   );
   gpc1_1 gpc3710 (
      {stage1_24[112]},
      {stage2_24[54]}
   );
   gpc1_1 gpc3711 (
      {stage1_24[113]},
      {stage2_24[55]}
   );
   gpc1_1 gpc3712 (
      {stage1_24[114]},
      {stage2_24[56]}
   );
   gpc1_1 gpc3713 (
      {stage1_24[115]},
      {stage2_24[57]}
   );
   gpc1_1 gpc3714 (
      {stage1_24[116]},
      {stage2_24[58]}
   );
   gpc1_1 gpc3715 (
      {stage1_24[117]},
      {stage2_24[59]}
   );
   gpc1_1 gpc3716 (
      {stage1_24[118]},
      {stage2_24[60]}
   );
   gpc1_1 gpc3717 (
      {stage1_24[119]},
      {stage2_24[61]}
   );
   gpc1_1 gpc3718 (
      {stage1_24[120]},
      {stage2_24[62]}
   );
   gpc1_1 gpc3719 (
      {stage1_24[121]},
      {stage2_24[63]}
   );
   gpc1_1 gpc3720 (
      {stage1_24[122]},
      {stage2_24[64]}
   );
   gpc1_1 gpc3721 (
      {stage1_24[123]},
      {stage2_24[65]}
   );
   gpc1_1 gpc3722 (
      {stage1_24[124]},
      {stage2_24[66]}
   );
   gpc1_1 gpc3723 (
      {stage1_24[125]},
      {stage2_24[67]}
   );
   gpc1_1 gpc3724 (
      {stage1_24[126]},
      {stage2_24[68]}
   );
   gpc1_1 gpc3725 (
      {stage1_24[127]},
      {stage2_24[69]}
   );
   gpc1_1 gpc3726 (
      {stage1_24[128]},
      {stage2_24[70]}
   );
   gpc1_1 gpc3727 (
      {stage1_24[129]},
      {stage2_24[71]}
   );
   gpc1_1 gpc3728 (
      {stage1_24[130]},
      {stage2_24[72]}
   );
   gpc1_1 gpc3729 (
      {stage1_24[131]},
      {stage2_24[73]}
   );
   gpc1_1 gpc3730 (
      {stage1_24[132]},
      {stage2_24[74]}
   );
   gpc1_1 gpc3731 (
      {stage1_24[133]},
      {stage2_24[75]}
   );
   gpc1_1 gpc3732 (
      {stage1_24[134]},
      {stage2_24[76]}
   );
   gpc1_1 gpc3733 (
      {stage1_24[135]},
      {stage2_24[77]}
   );
   gpc1_1 gpc3734 (
      {stage1_24[136]},
      {stage2_24[78]}
   );
   gpc1_1 gpc3735 (
      {stage1_24[137]},
      {stage2_24[79]}
   );
   gpc1_1 gpc3736 (
      {stage1_24[138]},
      {stage2_24[80]}
   );
   gpc1_1 gpc3737 (
      {stage1_24[139]},
      {stage2_24[81]}
   );
   gpc1_1 gpc3738 (
      {stage1_25[105]},
      {stage2_25[46]}
   );
   gpc1_1 gpc3739 (
      {stage1_25[106]},
      {stage2_25[47]}
   );
   gpc1_1 gpc3740 (
      {stage1_25[107]},
      {stage2_25[48]}
   );
   gpc1_1 gpc3741 (
      {stage1_25[108]},
      {stage2_25[49]}
   );
   gpc1_1 gpc3742 (
      {stage1_25[109]},
      {stage2_25[50]}
   );
   gpc1_1 gpc3743 (
      {stage1_26[129]},
      {stage2_26[40]}
   );
   gpc1_1 gpc3744 (
      {stage1_26[130]},
      {stage2_26[41]}
   );
   gpc1_1 gpc3745 (
      {stage1_26[131]},
      {stage2_26[42]}
   );
   gpc1_1 gpc3746 (
      {stage1_26[132]},
      {stage2_26[43]}
   );
   gpc1_1 gpc3747 (
      {stage1_26[133]},
      {stage2_26[44]}
   );
   gpc1_1 gpc3748 (
      {stage1_26[134]},
      {stage2_26[45]}
   );
   gpc1_1 gpc3749 (
      {stage1_26[135]},
      {stage2_26[46]}
   );
   gpc1_1 gpc3750 (
      {stage1_26[136]},
      {stage2_26[47]}
   );
   gpc1_1 gpc3751 (
      {stage1_26[137]},
      {stage2_26[48]}
   );
   gpc1_1 gpc3752 (
      {stage1_26[138]},
      {stage2_26[49]}
   );
   gpc1_1 gpc3753 (
      {stage1_26[139]},
      {stage2_26[50]}
   );
   gpc1_1 gpc3754 (
      {stage1_26[140]},
      {stage2_26[51]}
   );
   gpc1_1 gpc3755 (
      {stage1_27[93]},
      {stage2_27[46]}
   );
   gpc1_1 gpc3756 (
      {stage1_27[94]},
      {stage2_27[47]}
   );
   gpc1_1 gpc3757 (
      {stage1_27[95]},
      {stage2_27[48]}
   );
   gpc1_1 gpc3758 (
      {stage1_27[96]},
      {stage2_27[49]}
   );
   gpc1_1 gpc3759 (
      {stage1_27[97]},
      {stage2_27[50]}
   );
   gpc1_1 gpc3760 (
      {stage1_27[98]},
      {stage2_27[51]}
   );
   gpc1_1 gpc3761 (
      {stage1_27[99]},
      {stage2_27[52]}
   );
   gpc1_1 gpc3762 (
      {stage1_27[100]},
      {stage2_27[53]}
   );
   gpc1_1 gpc3763 (
      {stage1_27[101]},
      {stage2_27[54]}
   );
   gpc1_1 gpc3764 (
      {stage1_27[102]},
      {stage2_27[55]}
   );
   gpc1_1 gpc3765 (
      {stage1_27[103]},
      {stage2_27[56]}
   );
   gpc1_1 gpc3766 (
      {stage1_27[104]},
      {stage2_27[57]}
   );
   gpc1_1 gpc3767 (
      {stage1_27[105]},
      {stage2_27[58]}
   );
   gpc1_1 gpc3768 (
      {stage1_27[106]},
      {stage2_27[59]}
   );
   gpc1_1 gpc3769 (
      {stage1_27[107]},
      {stage2_27[60]}
   );
   gpc1_1 gpc3770 (
      {stage1_27[108]},
      {stage2_27[61]}
   );
   gpc1_1 gpc3771 (
      {stage1_27[109]},
      {stage2_27[62]}
   );
   gpc1_1 gpc3772 (
      {stage1_27[110]},
      {stage2_27[63]}
   );
   gpc1_1 gpc3773 (
      {stage1_27[111]},
      {stage2_27[64]}
   );
   gpc1_1 gpc3774 (
      {stage1_27[112]},
      {stage2_27[65]}
   );
   gpc1_1 gpc3775 (
      {stage1_27[113]},
      {stage2_27[66]}
   );
   gpc1_1 gpc3776 (
      {stage1_27[114]},
      {stage2_27[67]}
   );
   gpc1_1 gpc3777 (
      {stage1_27[115]},
      {stage2_27[68]}
   );
   gpc1_1 gpc3778 (
      {stage1_27[116]},
      {stage2_27[69]}
   );
   gpc1_1 gpc3779 (
      {stage1_27[117]},
      {stage2_27[70]}
   );
   gpc1_1 gpc3780 (
      {stage1_27[118]},
      {stage2_27[71]}
   );
   gpc1_1 gpc3781 (
      {stage1_28[104]},
      {stage2_28[50]}
   );
   gpc1_1 gpc3782 (
      {stage1_28[105]},
      {stage2_28[51]}
   );
   gpc1_1 gpc3783 (
      {stage1_28[106]},
      {stage2_28[52]}
   );
   gpc1_1 gpc3784 (
      {stage1_28[107]},
      {stage2_28[53]}
   );
   gpc1_1 gpc3785 (
      {stage1_28[108]},
      {stage2_28[54]}
   );
   gpc1_1 gpc3786 (
      {stage1_28[109]},
      {stage2_28[55]}
   );
   gpc1_1 gpc3787 (
      {stage1_28[110]},
      {stage2_28[56]}
   );
   gpc1_1 gpc3788 (
      {stage1_28[111]},
      {stage2_28[57]}
   );
   gpc1_1 gpc3789 (
      {stage1_28[112]},
      {stage2_28[58]}
   );
   gpc1_1 gpc3790 (
      {stage1_28[113]},
      {stage2_28[59]}
   );
   gpc1_1 gpc3791 (
      {stage1_28[114]},
      {stage2_28[60]}
   );
   gpc1_1 gpc3792 (
      {stage1_28[115]},
      {stage2_28[61]}
   );
   gpc1_1 gpc3793 (
      {stage1_28[116]},
      {stage2_28[62]}
   );
   gpc1_1 gpc3794 (
      {stage1_28[117]},
      {stage2_28[63]}
   );
   gpc1_1 gpc3795 (
      {stage1_28[118]},
      {stage2_28[64]}
   );
   gpc1_1 gpc3796 (
      {stage1_28[119]},
      {stage2_28[65]}
   );
   gpc1_1 gpc3797 (
      {stage1_28[120]},
      {stage2_28[66]}
   );
   gpc1_1 gpc3798 (
      {stage1_28[121]},
      {stage2_28[67]}
   );
   gpc1_1 gpc3799 (
      {stage1_28[122]},
      {stage2_28[68]}
   );
   gpc1_1 gpc3800 (
      {stage1_28[123]},
      {stage2_28[69]}
   );
   gpc1_1 gpc3801 (
      {stage1_28[124]},
      {stage2_28[70]}
   );
   gpc1_1 gpc3802 (
      {stage1_28[125]},
      {stage2_28[71]}
   );
   gpc1_1 gpc3803 (
      {stage1_28[126]},
      {stage2_28[72]}
   );
   gpc1_1 gpc3804 (
      {stage1_29[104]},
      {stage2_29[40]}
   );
   gpc1_1 gpc3805 (
      {stage1_29[105]},
      {stage2_29[41]}
   );
   gpc1_1 gpc3806 (
      {stage1_29[106]},
      {stage2_29[42]}
   );
   gpc1_1 gpc3807 (
      {stage1_29[107]},
      {stage2_29[43]}
   );
   gpc1_1 gpc3808 (
      {stage1_29[108]},
      {stage2_29[44]}
   );
   gpc1_1 gpc3809 (
      {stage1_29[109]},
      {stage2_29[45]}
   );
   gpc1_1 gpc3810 (
      {stage1_30[68]},
      {stage2_30[36]}
   );
   gpc1_1 gpc3811 (
      {stage1_30[69]},
      {stage2_30[37]}
   );
   gpc1_1 gpc3812 (
      {stage1_30[70]},
      {stage2_30[38]}
   );
   gpc1_1 gpc3813 (
      {stage1_30[71]},
      {stage2_30[39]}
   );
   gpc1_1 gpc3814 (
      {stage1_30[72]},
      {stage2_30[40]}
   );
   gpc1_1 gpc3815 (
      {stage1_30[73]},
      {stage2_30[41]}
   );
   gpc1_1 gpc3816 (
      {stage1_30[74]},
      {stage2_30[42]}
   );
   gpc1_1 gpc3817 (
      {stage1_30[75]},
      {stage2_30[43]}
   );
   gpc1_1 gpc3818 (
      {stage1_30[76]},
      {stage2_30[44]}
   );
   gpc1_1 gpc3819 (
      {stage1_30[77]},
      {stage2_30[45]}
   );
   gpc1_1 gpc3820 (
      {stage1_30[78]},
      {stage2_30[46]}
   );
   gpc1_1 gpc3821 (
      {stage1_30[79]},
      {stage2_30[47]}
   );
   gpc1_1 gpc3822 (
      {stage1_30[80]},
      {stage2_30[48]}
   );
   gpc1_1 gpc3823 (
      {stage1_30[81]},
      {stage2_30[49]}
   );
   gpc1_1 gpc3824 (
      {stage1_30[82]},
      {stage2_30[50]}
   );
   gpc1_1 gpc3825 (
      {stage1_30[83]},
      {stage2_30[51]}
   );
   gpc1_1 gpc3826 (
      {stage1_30[84]},
      {stage2_30[52]}
   );
   gpc1_1 gpc3827 (
      {stage1_30[85]},
      {stage2_30[53]}
   );
   gpc1_1 gpc3828 (
      {stage1_30[86]},
      {stage2_30[54]}
   );
   gpc1_1 gpc3829 (
      {stage1_30[87]},
      {stage2_30[55]}
   );
   gpc1_1 gpc3830 (
      {stage1_30[88]},
      {stage2_30[56]}
   );
   gpc1_1 gpc3831 (
      {stage1_30[89]},
      {stage2_30[57]}
   );
   gpc1_1 gpc3832 (
      {stage1_30[90]},
      {stage2_30[58]}
   );
   gpc1_1 gpc3833 (
      {stage1_31[99]},
      {stage2_31[38]}
   );
   gpc1_1 gpc3834 (
      {stage1_31[100]},
      {stage2_31[39]}
   );
   gpc1_1 gpc3835 (
      {stage1_31[101]},
      {stage2_31[40]}
   );
   gpc1_1 gpc3836 (
      {stage1_31[102]},
      {stage2_31[41]}
   );
   gpc1_1 gpc3837 (
      {stage1_31[103]},
      {stage2_31[42]}
   );
   gpc1_1 gpc3838 (
      {stage1_31[104]},
      {stage2_31[43]}
   );
   gpc1_1 gpc3839 (
      {stage1_31[105]},
      {stage2_31[44]}
   );
   gpc1_1 gpc3840 (
      {stage1_31[106]},
      {stage2_31[45]}
   );
   gpc1_1 gpc3841 (
      {stage1_31[107]},
      {stage2_31[46]}
   );
   gpc1_1 gpc3842 (
      {stage1_31[108]},
      {stage2_31[47]}
   );
   gpc1_1 gpc3843 (
      {stage1_31[109]},
      {stage2_31[48]}
   );
   gpc1_1 gpc3844 (
      {stage1_31[110]},
      {stage2_31[49]}
   );
   gpc1_1 gpc3845 (
      {stage1_31[111]},
      {stage2_31[50]}
   );
   gpc1_1 gpc3846 (
      {stage1_31[112]},
      {stage2_31[51]}
   );
   gpc1_1 gpc3847 (
      {stage1_31[113]},
      {stage2_31[52]}
   );
   gpc1_1 gpc3848 (
      {stage1_31[114]},
      {stage2_31[53]}
   );
   gpc1_1 gpc3849 (
      {stage1_32[112]},
      {stage2_32[44]}
   );
   gpc1_1 gpc3850 (
      {stage1_32[113]},
      {stage2_32[45]}
   );
   gpc1_1 gpc3851 (
      {stage1_32[114]},
      {stage2_32[46]}
   );
   gpc1_1 gpc3852 (
      {stage1_33[102]},
      {stage2_33[43]}
   );
   gpc1_1 gpc3853 (
      {stage1_33[103]},
      {stage2_33[44]}
   );
   gpc1_1 gpc3854 (
      {stage1_33[104]},
      {stage2_33[45]}
   );
   gpc1_1 gpc3855 (
      {stage1_33[105]},
      {stage2_33[46]}
   );
   gpc1_1 gpc3856 (
      {stage1_33[106]},
      {stage2_33[47]}
   );
   gpc1_1 gpc3857 (
      {stage1_33[107]},
      {stage2_33[48]}
   );
   gpc1_1 gpc3858 (
      {stage1_33[108]},
      {stage2_33[49]}
   );
   gpc1_1 gpc3859 (
      {stage1_33[109]},
      {stage2_33[50]}
   );
   gpc1_1 gpc3860 (
      {stage1_33[110]},
      {stage2_33[51]}
   );
   gpc1_1 gpc3861 (
      {stage1_35[106]},
      {stage2_35[46]}
   );
   gpc1_1 gpc3862 (
      {stage1_35[107]},
      {stage2_35[47]}
   );
   gpc1_1 gpc3863 (
      {stage1_35[108]},
      {stage2_35[48]}
   );
   gpc1_1 gpc3864 (
      {stage1_35[109]},
      {stage2_35[49]}
   );
   gpc1_1 gpc3865 (
      {stage1_35[110]},
      {stage2_35[50]}
   );
   gpc1_1 gpc3866 (
      {stage1_35[111]},
      {stage2_35[51]}
   );
   gpc1_1 gpc3867 (
      {stage1_35[112]},
      {stage2_35[52]}
   );
   gpc1_1 gpc3868 (
      {stage1_35[113]},
      {stage2_35[53]}
   );
   gpc1_1 gpc3869 (
      {stage1_35[114]},
      {stage2_35[54]}
   );
   gpc1_1 gpc3870 (
      {stage1_35[115]},
      {stage2_35[55]}
   );
   gpc1_1 gpc3871 (
      {stage1_35[116]},
      {stage2_35[56]}
   );
   gpc1_1 gpc3872 (
      {stage1_35[117]},
      {stage2_35[57]}
   );
   gpc1_1 gpc3873 (
      {stage1_35[118]},
      {stage2_35[58]}
   );
   gpc1_1 gpc3874 (
      {stage1_36[138]},
      {stage2_36[56]}
   );
   gpc1_1 gpc3875 (
      {stage1_36[139]},
      {stage2_36[57]}
   );
   gpc1_1 gpc3876 (
      {stage1_36[140]},
      {stage2_36[58]}
   );
   gpc1_1 gpc3877 (
      {stage1_36[141]},
      {stage2_36[59]}
   );
   gpc1_1 gpc3878 (
      {stage1_36[142]},
      {stage2_36[60]}
   );
   gpc1_1 gpc3879 (
      {stage1_36[143]},
      {stage2_36[61]}
   );
   gpc1_1 gpc3880 (
      {stage1_36[144]},
      {stage2_36[62]}
   );
   gpc1_1 gpc3881 (
      {stage1_37[93]},
      {stage2_37[43]}
   );
   gpc1_1 gpc3882 (
      {stage1_37[94]},
      {stage2_37[44]}
   );
   gpc1_1 gpc3883 (
      {stage1_37[95]},
      {stage2_37[45]}
   );
   gpc1_1 gpc3884 (
      {stage1_37[96]},
      {stage2_37[46]}
   );
   gpc1_1 gpc3885 (
      {stage1_37[97]},
      {stage2_37[47]}
   );
   gpc1_1 gpc3886 (
      {stage1_37[98]},
      {stage2_37[48]}
   );
   gpc1_1 gpc3887 (
      {stage1_37[99]},
      {stage2_37[49]}
   );
   gpc1_1 gpc3888 (
      {stage1_37[100]},
      {stage2_37[50]}
   );
   gpc1_1 gpc3889 (
      {stage1_37[101]},
      {stage2_37[51]}
   );
   gpc1_1 gpc3890 (
      {stage1_37[102]},
      {stage2_37[52]}
   );
   gpc1_1 gpc3891 (
      {stage1_37[103]},
      {stage2_37[53]}
   );
   gpc1_1 gpc3892 (
      {stage1_37[104]},
      {stage2_37[54]}
   );
   gpc1_1 gpc3893 (
      {stage1_38[134]},
      {stage2_38[44]}
   );
   gpc1_1 gpc3894 (
      {stage1_38[135]},
      {stage2_38[45]}
   );
   gpc1_1 gpc3895 (
      {stage1_38[136]},
      {stage2_38[46]}
   );
   gpc1_1 gpc3896 (
      {stage1_39[98]},
      {stage2_39[54]}
   );
   gpc1_1 gpc3897 (
      {stage1_39[99]},
      {stage2_39[55]}
   );
   gpc1_1 gpc3898 (
      {stage1_39[100]},
      {stage2_39[56]}
   );
   gpc1_1 gpc3899 (
      {stage1_39[101]},
      {stage2_39[57]}
   );
   gpc1_1 gpc3900 (
      {stage1_39[102]},
      {stage2_39[58]}
   );
   gpc1_1 gpc3901 (
      {stage1_39[103]},
      {stage2_39[59]}
   );
   gpc1_1 gpc3902 (
      {stage1_39[104]},
      {stage2_39[60]}
   );
   gpc1_1 gpc3903 (
      {stage1_39[105]},
      {stage2_39[61]}
   );
   gpc1_1 gpc3904 (
      {stage1_39[106]},
      {stage2_39[62]}
   );
   gpc1_1 gpc3905 (
      {stage1_39[107]},
      {stage2_39[63]}
   );
   gpc1_1 gpc3906 (
      {stage1_39[108]},
      {stage2_39[64]}
   );
   gpc1_1 gpc3907 (
      {stage1_39[109]},
      {stage2_39[65]}
   );
   gpc1_1 gpc3908 (
      {stage1_39[110]},
      {stage2_39[66]}
   );
   gpc1_1 gpc3909 (
      {stage1_39[111]},
      {stage2_39[67]}
   );
   gpc1_1 gpc3910 (
      {stage1_39[112]},
      {stage2_39[68]}
   );
   gpc1_1 gpc3911 (
      {stage1_39[113]},
      {stage2_39[69]}
   );
   gpc1_1 gpc3912 (
      {stage1_39[114]},
      {stage2_39[70]}
   );
   gpc1_1 gpc3913 (
      {stage1_39[115]},
      {stage2_39[71]}
   );
   gpc1_1 gpc3914 (
      {stage1_39[116]},
      {stage2_39[72]}
   );
   gpc1_1 gpc3915 (
      {stage1_39[117]},
      {stage2_39[73]}
   );
   gpc1_1 gpc3916 (
      {stage1_39[118]},
      {stage2_39[74]}
   );
   gpc1_1 gpc3917 (
      {stage1_39[119]},
      {stage2_39[75]}
   );
   gpc1_1 gpc3918 (
      {stage1_39[120]},
      {stage2_39[76]}
   );
   gpc1_1 gpc3919 (
      {stage1_39[121]},
      {stage2_39[77]}
   );
   gpc1_1 gpc3920 (
      {stage1_39[122]},
      {stage2_39[78]}
   );
   gpc1_1 gpc3921 (
      {stage1_39[123]},
      {stage2_39[79]}
   );
   gpc1_1 gpc3922 (
      {stage1_39[124]},
      {stage2_39[80]}
   );
   gpc1_1 gpc3923 (
      {stage1_40[91]},
      {stage2_40[44]}
   );
   gpc1_1 gpc3924 (
      {stage1_41[102]},
      {stage2_41[34]}
   );
   gpc1_1 gpc3925 (
      {stage1_41[103]},
      {stage2_41[35]}
   );
   gpc1_1 gpc3926 (
      {stage1_41[104]},
      {stage2_41[36]}
   );
   gpc1_1 gpc3927 (
      {stage1_41[105]},
      {stage2_41[37]}
   );
   gpc1_1 gpc3928 (
      {stage1_41[106]},
      {stage2_41[38]}
   );
   gpc1_1 gpc3929 (
      {stage1_41[107]},
      {stage2_41[39]}
   );
   gpc1_1 gpc3930 (
      {stage1_41[108]},
      {stage2_41[40]}
   );
   gpc1_1 gpc3931 (
      {stage1_41[109]},
      {stage2_41[41]}
   );
   gpc1_1 gpc3932 (
      {stage1_41[110]},
      {stage2_41[42]}
   );
   gpc1_1 gpc3933 (
      {stage1_41[111]},
      {stage2_41[43]}
   );
   gpc1_1 gpc3934 (
      {stage1_41[112]},
      {stage2_41[44]}
   );
   gpc1_1 gpc3935 (
      {stage1_41[113]},
      {stage2_41[45]}
   );
   gpc1_1 gpc3936 (
      {stage1_41[114]},
      {stage2_41[46]}
   );
   gpc1_1 gpc3937 (
      {stage1_41[115]},
      {stage2_41[47]}
   );
   gpc1_1 gpc3938 (
      {stage1_41[116]},
      {stage2_41[48]}
   );
   gpc1_1 gpc3939 (
      {stage1_41[117]},
      {stage2_41[49]}
   );
   gpc1_1 gpc3940 (
      {stage1_41[118]},
      {stage2_41[50]}
   );
   gpc1_1 gpc3941 (
      {stage1_41[119]},
      {stage2_41[51]}
   );
   gpc1_1 gpc3942 (
      {stage1_41[120]},
      {stage2_41[52]}
   );
   gpc1_1 gpc3943 (
      {stage1_41[121]},
      {stage2_41[53]}
   );
   gpc1_1 gpc3944 (
      {stage1_41[122]},
      {stage2_41[54]}
   );
   gpc1_1 gpc3945 (
      {stage1_41[123]},
      {stage2_41[55]}
   );
   gpc1_1 gpc3946 (
      {stage1_41[124]},
      {stage2_41[56]}
   );
   gpc1_1 gpc3947 (
      {stage1_41[125]},
      {stage2_41[57]}
   );
   gpc1_1 gpc3948 (
      {stage1_41[126]},
      {stage2_41[58]}
   );
   gpc1_1 gpc3949 (
      {stage1_41[127]},
      {stage2_41[59]}
   );
   gpc1_1 gpc3950 (
      {stage1_41[128]},
      {stage2_41[60]}
   );
   gpc1_1 gpc3951 (
      {stage1_41[129]},
      {stage2_41[61]}
   );
   gpc1_1 gpc3952 (
      {stage1_41[130]},
      {stage2_41[62]}
   );
   gpc1_1 gpc3953 (
      {stage1_41[131]},
      {stage2_41[63]}
   );
   gpc1_1 gpc3954 (
      {stage1_41[132]},
      {stage2_41[64]}
   );
   gpc1_1 gpc3955 (
      {stage1_41[133]},
      {stage2_41[65]}
   );
   gpc1_1 gpc3956 (
      {stage1_41[134]},
      {stage2_41[66]}
   );
   gpc1_1 gpc3957 (
      {stage1_41[135]},
      {stage2_41[67]}
   );
   gpc1_1 gpc3958 (
      {stage1_41[136]},
      {stage2_41[68]}
   );
   gpc1_1 gpc3959 (
      {stage1_41[137]},
      {stage2_41[69]}
   );
   gpc1_1 gpc3960 (
      {stage1_41[138]},
      {stage2_41[70]}
   );
   gpc1_1 gpc3961 (
      {stage1_41[139]},
      {stage2_41[71]}
   );
   gpc1_1 gpc3962 (
      {stage1_41[140]},
      {stage2_41[72]}
   );
   gpc1_1 gpc3963 (
      {stage1_41[141]},
      {stage2_41[73]}
   );
   gpc1_1 gpc3964 (
      {stage1_41[142]},
      {stage2_41[74]}
   );
   gpc1_1 gpc3965 (
      {stage1_42[162]},
      {stage2_42[53]}
   );
   gpc1_1 gpc3966 (
      {stage1_42[163]},
      {stage2_42[54]}
   );
   gpc1_1 gpc3967 (
      {stage1_42[164]},
      {stage2_42[55]}
   );
   gpc1_1 gpc3968 (
      {stage1_42[165]},
      {stage2_42[56]}
   );
   gpc1_1 gpc3969 (
      {stage1_42[166]},
      {stage2_42[57]}
   );
   gpc1_1 gpc3970 (
      {stage1_42[167]},
      {stage2_42[58]}
   );
   gpc1_1 gpc3971 (
      {stage1_42[168]},
      {stage2_42[59]}
   );
   gpc1_1 gpc3972 (
      {stage1_42[169]},
      {stage2_42[60]}
   );
   gpc1_1 gpc3973 (
      {stage1_42[170]},
      {stage2_42[61]}
   );
   gpc1_1 gpc3974 (
      {stage1_42[171]},
      {stage2_42[62]}
   );
   gpc1_1 gpc3975 (
      {stage1_43[70]},
      {stage2_43[53]}
   );
   gpc1_1 gpc3976 (
      {stage1_43[71]},
      {stage2_43[54]}
   );
   gpc1_1 gpc3977 (
      {stage1_43[72]},
      {stage2_43[55]}
   );
   gpc1_1 gpc3978 (
      {stage1_43[73]},
      {stage2_43[56]}
   );
   gpc1_1 gpc3979 (
      {stage1_43[74]},
      {stage2_43[57]}
   );
   gpc1_1 gpc3980 (
      {stage1_43[75]},
      {stage2_43[58]}
   );
   gpc1_1 gpc3981 (
      {stage1_43[76]},
      {stage2_43[59]}
   );
   gpc1_1 gpc3982 (
      {stage1_43[77]},
      {stage2_43[60]}
   );
   gpc1_1 gpc3983 (
      {stage1_43[78]},
      {stage2_43[61]}
   );
   gpc1_1 gpc3984 (
      {stage1_44[134]},
      {stage2_44[40]}
   );
   gpc1_1 gpc3985 (
      {stage1_44[135]},
      {stage2_44[41]}
   );
   gpc1_1 gpc3986 (
      {stage1_44[136]},
      {stage2_44[42]}
   );
   gpc1_1 gpc3987 (
      {stage1_44[137]},
      {stage2_44[43]}
   );
   gpc1_1 gpc3988 (
      {stage1_44[138]},
      {stage2_44[44]}
   );
   gpc1_1 gpc3989 (
      {stage1_44[139]},
      {stage2_44[45]}
   );
   gpc1_1 gpc3990 (
      {stage1_44[140]},
      {stage2_44[46]}
   );
   gpc1_1 gpc3991 (
      {stage1_44[141]},
      {stage2_44[47]}
   );
   gpc1_1 gpc3992 (
      {stage1_44[142]},
      {stage2_44[48]}
   );
   gpc1_1 gpc3993 (
      {stage1_44[143]},
      {stage2_44[49]}
   );
   gpc1_1 gpc3994 (
      {stage1_44[144]},
      {stage2_44[50]}
   );
   gpc1_1 gpc3995 (
      {stage1_44[145]},
      {stage2_44[51]}
   );
   gpc1_1 gpc3996 (
      {stage1_45[126]},
      {stage2_45[46]}
   );
   gpc1_1 gpc3997 (
      {stage1_45[127]},
      {stage2_45[47]}
   );
   gpc1_1 gpc3998 (
      {stage1_45[128]},
      {stage2_45[48]}
   );
   gpc1_1 gpc3999 (
      {stage1_45[129]},
      {stage2_45[49]}
   );
   gpc1_1 gpc4000 (
      {stage1_45[130]},
      {stage2_45[50]}
   );
   gpc1_1 gpc4001 (
      {stage1_45[131]},
      {stage2_45[51]}
   );
   gpc1_1 gpc4002 (
      {stage1_45[132]},
      {stage2_45[52]}
   );
   gpc1_1 gpc4003 (
      {stage1_45[133]},
      {stage2_45[53]}
   );
   gpc1_1 gpc4004 (
      {stage1_45[134]},
      {stage2_45[54]}
   );
   gpc1_1 gpc4005 (
      {stage1_45[135]},
      {stage2_45[55]}
   );
   gpc1_1 gpc4006 (
      {stage1_45[136]},
      {stage2_45[56]}
   );
   gpc1_1 gpc4007 (
      {stage1_45[137]},
      {stage2_45[57]}
   );
   gpc1_1 gpc4008 (
      {stage1_45[138]},
      {stage2_45[58]}
   );
   gpc1_1 gpc4009 (
      {stage1_45[139]},
      {stage2_45[59]}
   );
   gpc1_1 gpc4010 (
      {stage1_45[140]},
      {stage2_45[60]}
   );
   gpc1_1 gpc4011 (
      {stage1_45[141]},
      {stage2_45[61]}
   );
   gpc1_1 gpc4012 (
      {stage1_45[142]},
      {stage2_45[62]}
   );
   gpc1_1 gpc4013 (
      {stage1_45[143]},
      {stage2_45[63]}
   );
   gpc1_1 gpc4014 (
      {stage1_45[144]},
      {stage2_45[64]}
   );
   gpc1_1 gpc4015 (
      {stage1_45[145]},
      {stage2_45[65]}
   );
   gpc1_1 gpc4016 (
      {stage1_45[146]},
      {stage2_45[66]}
   );
   gpc1_1 gpc4017 (
      {stage1_45[147]},
      {stage2_45[67]}
   );
   gpc1_1 gpc4018 (
      {stage1_45[148]},
      {stage2_45[68]}
   );
   gpc1_1 gpc4019 (
      {stage1_45[149]},
      {stage2_45[69]}
   );
   gpc1_1 gpc4020 (
      {stage1_45[150]},
      {stage2_45[70]}
   );
   gpc1_1 gpc4021 (
      {stage1_45[151]},
      {stage2_45[71]}
   );
   gpc1_1 gpc4022 (
      {stage1_45[152]},
      {stage2_45[72]}
   );
   gpc1_1 gpc4023 (
      {stage1_45[153]},
      {stage2_45[73]}
   );
   gpc1_1 gpc4024 (
      {stage1_45[154]},
      {stage2_45[74]}
   );
   gpc1_1 gpc4025 (
      {stage1_45[155]},
      {stage2_45[75]}
   );
   gpc1_1 gpc4026 (
      {stage1_45[156]},
      {stage2_45[76]}
   );
   gpc1_1 gpc4027 (
      {stage1_45[157]},
      {stage2_45[77]}
   );
   gpc1_1 gpc4028 (
      {stage1_45[158]},
      {stage2_45[78]}
   );
   gpc1_1 gpc4029 (
      {stage1_46[96]},
      {stage2_46[58]}
   );
   gpc1_1 gpc4030 (
      {stage1_46[97]},
      {stage2_46[59]}
   );
   gpc1_1 gpc4031 (
      {stage1_46[98]},
      {stage2_46[60]}
   );
   gpc1_1 gpc4032 (
      {stage1_46[99]},
      {stage2_46[61]}
   );
   gpc1_1 gpc4033 (
      {stage1_46[100]},
      {stage2_46[62]}
   );
   gpc1_1 gpc4034 (
      {stage1_47[102]},
      {stage2_47[43]}
   );
   gpc1_1 gpc4035 (
      {stage1_47[103]},
      {stage2_47[44]}
   );
   gpc1_1 gpc4036 (
      {stage1_47[104]},
      {stage2_47[45]}
   );
   gpc1_1 gpc4037 (
      {stage1_47[105]},
      {stage2_47[46]}
   );
   gpc1_1 gpc4038 (
      {stage1_47[106]},
      {stage2_47[47]}
   );
   gpc1_1 gpc4039 (
      {stage1_47[107]},
      {stage2_47[48]}
   );
   gpc1_1 gpc4040 (
      {stage1_47[108]},
      {stage2_47[49]}
   );
   gpc1_1 gpc4041 (
      {stage1_47[109]},
      {stage2_47[50]}
   );
   gpc1_1 gpc4042 (
      {stage1_47[110]},
      {stage2_47[51]}
   );
   gpc1_1 gpc4043 (
      {stage1_47[111]},
      {stage2_47[52]}
   );
   gpc1_1 gpc4044 (
      {stage1_47[112]},
      {stage2_47[53]}
   );
   gpc1_1 gpc4045 (
      {stage1_47[113]},
      {stage2_47[54]}
   );
   gpc1_1 gpc4046 (
      {stage1_47[114]},
      {stage2_47[55]}
   );
   gpc1_1 gpc4047 (
      {stage1_47[115]},
      {stage2_47[56]}
   );
   gpc1_1 gpc4048 (
      {stage1_47[116]},
      {stage2_47[57]}
   );
   gpc1_1 gpc4049 (
      {stage1_47[117]},
      {stage2_47[58]}
   );
   gpc1_1 gpc4050 (
      {stage1_47[118]},
      {stage2_47[59]}
   );
   gpc1_1 gpc4051 (
      {stage1_47[119]},
      {stage2_47[60]}
   );
   gpc1_1 gpc4052 (
      {stage1_47[120]},
      {stage2_47[61]}
   );
   gpc1_1 gpc4053 (
      {stage1_47[121]},
      {stage2_47[62]}
   );
   gpc1_1 gpc4054 (
      {stage1_47[122]},
      {stage2_47[63]}
   );
   gpc1_1 gpc4055 (
      {stage1_47[123]},
      {stage2_47[64]}
   );
   gpc1_1 gpc4056 (
      {stage1_47[124]},
      {stage2_47[65]}
   );
   gpc1_1 gpc4057 (
      {stage1_47[125]},
      {stage2_47[66]}
   );
   gpc1_1 gpc4058 (
      {stage1_47[126]},
      {stage2_47[67]}
   );
   gpc1_1 gpc4059 (
      {stage1_47[127]},
      {stage2_47[68]}
   );
   gpc1_1 gpc4060 (
      {stage1_47[128]},
      {stage2_47[69]}
   );
   gpc1_1 gpc4061 (
      {stage1_47[129]},
      {stage2_47[70]}
   );
   gpc1_1 gpc4062 (
      {stage1_48[100]},
      {stage2_48[34]}
   );
   gpc1_1 gpc4063 (
      {stage1_48[101]},
      {stage2_48[35]}
   );
   gpc1_1 gpc4064 (
      {stage1_48[102]},
      {stage2_48[36]}
   );
   gpc1_1 gpc4065 (
      {stage1_48[103]},
      {stage2_48[37]}
   );
   gpc1_1 gpc4066 (
      {stage1_48[104]},
      {stage2_48[38]}
   );
   gpc1_1 gpc4067 (
      {stage1_48[105]},
      {stage2_48[39]}
   );
   gpc1_1 gpc4068 (
      {stage1_48[106]},
      {stage2_48[40]}
   );
   gpc1_1 gpc4069 (
      {stage1_48[107]},
      {stage2_48[41]}
   );
   gpc1_1 gpc4070 (
      {stage1_49[78]},
      {stage2_49[41]}
   );
   gpc1_1 gpc4071 (
      {stage1_49[79]},
      {stage2_49[42]}
   );
   gpc1_1 gpc4072 (
      {stage1_49[80]},
      {stage2_49[43]}
   );
   gpc1_1 gpc4073 (
      {stage1_49[81]},
      {stage2_49[44]}
   );
   gpc1_1 gpc4074 (
      {stage1_49[82]},
      {stage2_49[45]}
   );
   gpc1_1 gpc4075 (
      {stage1_49[83]},
      {stage2_49[46]}
   );
   gpc1_1 gpc4076 (
      {stage1_49[84]},
      {stage2_49[47]}
   );
   gpc1_1 gpc4077 (
      {stage1_49[85]},
      {stage2_49[48]}
   );
   gpc1_1 gpc4078 (
      {stage1_49[86]},
      {stage2_49[49]}
   );
   gpc1_1 gpc4079 (
      {stage1_49[87]},
      {stage2_49[50]}
   );
   gpc1_1 gpc4080 (
      {stage1_49[88]},
      {stage2_49[51]}
   );
   gpc1_1 gpc4081 (
      {stage1_49[89]},
      {stage2_49[52]}
   );
   gpc1_1 gpc4082 (
      {stage1_49[90]},
      {stage2_49[53]}
   );
   gpc1_1 gpc4083 (
      {stage1_49[91]},
      {stage2_49[54]}
   );
   gpc1_1 gpc4084 (
      {stage1_49[92]},
      {stage2_49[55]}
   );
   gpc1_1 gpc4085 (
      {stage1_49[93]},
      {stage2_49[56]}
   );
   gpc1_1 gpc4086 (
      {stage1_49[94]},
      {stage2_49[57]}
   );
   gpc1_1 gpc4087 (
      {stage1_49[95]},
      {stage2_49[58]}
   );
   gpc1_1 gpc4088 (
      {stage1_49[96]},
      {stage2_49[59]}
   );
   gpc1_1 gpc4089 (
      {stage1_49[97]},
      {stage2_49[60]}
   );
   gpc1_1 gpc4090 (
      {stage1_49[98]},
      {stage2_49[61]}
   );
   gpc1_1 gpc4091 (
      {stage1_49[99]},
      {stage2_49[62]}
   );
   gpc1_1 gpc4092 (
      {stage1_49[100]},
      {stage2_49[63]}
   );
   gpc1_1 gpc4093 (
      {stage1_49[101]},
      {stage2_49[64]}
   );
   gpc1_1 gpc4094 (
      {stage1_49[102]},
      {stage2_49[65]}
   );
   gpc1_1 gpc4095 (
      {stage1_49[103]},
      {stage2_49[66]}
   );
   gpc1_1 gpc4096 (
      {stage1_49[104]},
      {stage2_49[67]}
   );
   gpc1_1 gpc4097 (
      {stage1_49[105]},
      {stage2_49[68]}
   );
   gpc1_1 gpc4098 (
      {stage1_49[106]},
      {stage2_49[69]}
   );
   gpc1_1 gpc4099 (
      {stage1_49[107]},
      {stage2_49[70]}
   );
   gpc1_1 gpc4100 (
      {stage1_49[108]},
      {stage2_49[71]}
   );
   gpc1_1 gpc4101 (
      {stage1_49[109]},
      {stage2_49[72]}
   );
   gpc1_1 gpc4102 (
      {stage1_49[110]},
      {stage2_49[73]}
   );
   gpc1_1 gpc4103 (
      {stage1_49[111]},
      {stage2_49[74]}
   );
   gpc1_1 gpc4104 (
      {stage1_49[112]},
      {stage2_49[75]}
   );
   gpc1_1 gpc4105 (
      {stage1_49[113]},
      {stage2_49[76]}
   );
   gpc1_1 gpc4106 (
      {stage1_49[114]},
      {stage2_49[77]}
   );
   gpc1_1 gpc4107 (
      {stage1_49[115]},
      {stage2_49[78]}
   );
   gpc1_1 gpc4108 (
      {stage1_49[116]},
      {stage2_49[79]}
   );
   gpc1_1 gpc4109 (
      {stage1_49[117]},
      {stage2_49[80]}
   );
   gpc1_1 gpc4110 (
      {stage1_49[118]},
      {stage2_49[81]}
   );
   gpc1_1 gpc4111 (
      {stage1_49[119]},
      {stage2_49[82]}
   );
   gpc1_1 gpc4112 (
      {stage1_49[120]},
      {stage2_49[83]}
   );
   gpc1_1 gpc4113 (
      {stage1_49[121]},
      {stage2_49[84]}
   );
   gpc1_1 gpc4114 (
      {stage1_49[122]},
      {stage2_49[85]}
   );
   gpc1_1 gpc4115 (
      {stage1_49[123]},
      {stage2_49[86]}
   );
   gpc1_1 gpc4116 (
      {stage1_49[124]},
      {stage2_49[87]}
   );
   gpc1_1 gpc4117 (
      {stage1_49[125]},
      {stage2_49[88]}
   );
   gpc1_1 gpc4118 (
      {stage1_49[126]},
      {stage2_49[89]}
   );
   gpc1_1 gpc4119 (
      {stage1_49[127]},
      {stage2_49[90]}
   );
   gpc1_1 gpc4120 (
      {stage1_49[128]},
      {stage2_49[91]}
   );
   gpc1_1 gpc4121 (
      {stage1_49[129]},
      {stage2_49[92]}
   );
   gpc1_1 gpc4122 (
      {stage1_49[130]},
      {stage2_49[93]}
   );
   gpc1_1 gpc4123 (
      {stage1_49[131]},
      {stage2_49[94]}
   );
   gpc1_1 gpc4124 (
      {stage1_49[132]},
      {stage2_49[95]}
   );
   gpc1_1 gpc4125 (
      {stage1_49[133]},
      {stage2_49[96]}
   );
   gpc1_1 gpc4126 (
      {stage1_49[134]},
      {stage2_49[97]}
   );
   gpc1_1 gpc4127 (
      {stage1_49[135]},
      {stage2_49[98]}
   );
   gpc1_1 gpc4128 (
      {stage1_49[136]},
      {stage2_49[99]}
   );
   gpc1_1 gpc4129 (
      {stage1_49[137]},
      {stage2_49[100]}
   );
   gpc1_1 gpc4130 (
      {stage1_49[138]},
      {stage2_49[101]}
   );
   gpc1_1 gpc4131 (
      {stage1_49[139]},
      {stage2_49[102]}
   );
   gpc1_1 gpc4132 (
      {stage1_49[140]},
      {stage2_49[103]}
   );
   gpc1_1 gpc4133 (
      {stage1_49[141]},
      {stage2_49[104]}
   );
   gpc1_1 gpc4134 (
      {stage1_49[142]},
      {stage2_49[105]}
   );
   gpc1_1 gpc4135 (
      {stage1_49[143]},
      {stage2_49[106]}
   );
   gpc1_1 gpc4136 (
      {stage1_49[144]},
      {stage2_49[107]}
   );
   gpc1_1 gpc4137 (
      {stage1_49[145]},
      {stage2_49[108]}
   );
   gpc1_1 gpc4138 (
      {stage1_49[146]},
      {stage2_49[109]}
   );
   gpc1_1 gpc4139 (
      {stage1_49[147]},
      {stage2_49[110]}
   );
   gpc1_1 gpc4140 (
      {stage1_49[148]},
      {stage2_49[111]}
   );
   gpc1_1 gpc4141 (
      {stage1_49[149]},
      {stage2_49[112]}
   );
   gpc1_1 gpc4142 (
      {stage1_49[150]},
      {stage2_49[113]}
   );
   gpc1_1 gpc4143 (
      {stage1_49[151]},
      {stage2_49[114]}
   );
   gpc1_1 gpc4144 (
      {stage1_50[75]},
      {stage2_50[44]}
   );
   gpc1_1 gpc4145 (
      {stage1_50[76]},
      {stage2_50[45]}
   );
   gpc1_1 gpc4146 (
      {stage1_50[77]},
      {stage2_50[46]}
   );
   gpc1_1 gpc4147 (
      {stage1_50[78]},
      {stage2_50[47]}
   );
   gpc1_1 gpc4148 (
      {stage1_50[79]},
      {stage2_50[48]}
   );
   gpc1_1 gpc4149 (
      {stage1_50[80]},
      {stage2_50[49]}
   );
   gpc1_1 gpc4150 (
      {stage1_50[81]},
      {stage2_50[50]}
   );
   gpc1_1 gpc4151 (
      {stage1_50[82]},
      {stage2_50[51]}
   );
   gpc1_1 gpc4152 (
      {stage1_50[83]},
      {stage2_50[52]}
   );
   gpc1_1 gpc4153 (
      {stage1_50[84]},
      {stage2_50[53]}
   );
   gpc1_1 gpc4154 (
      {stage1_50[85]},
      {stage2_50[54]}
   );
   gpc1_1 gpc4155 (
      {stage1_50[86]},
      {stage2_50[55]}
   );
   gpc1_1 gpc4156 (
      {stage1_50[87]},
      {stage2_50[56]}
   );
   gpc1_1 gpc4157 (
      {stage1_50[88]},
      {stage2_50[57]}
   );
   gpc1_1 gpc4158 (
      {stage1_50[89]},
      {stage2_50[58]}
   );
   gpc1_1 gpc4159 (
      {stage1_50[90]},
      {stage2_50[59]}
   );
   gpc1_1 gpc4160 (
      {stage1_50[91]},
      {stage2_50[60]}
   );
   gpc1_1 gpc4161 (
      {stage1_50[92]},
      {stage2_50[61]}
   );
   gpc1_1 gpc4162 (
      {stage1_50[93]},
      {stage2_50[62]}
   );
   gpc1_1 gpc4163 (
      {stage1_50[94]},
      {stage2_50[63]}
   );
   gpc1_1 gpc4164 (
      {stage1_50[95]},
      {stage2_50[64]}
   );
   gpc1_1 gpc4165 (
      {stage1_50[96]},
      {stage2_50[65]}
   );
   gpc1_1 gpc4166 (
      {stage1_50[97]},
      {stage2_50[66]}
   );
   gpc1_1 gpc4167 (
      {stage1_50[98]},
      {stage2_50[67]}
   );
   gpc1_1 gpc4168 (
      {stage1_51[55]},
      {stage2_51[28]}
   );
   gpc1_1 gpc4169 (
      {stage1_51[56]},
      {stage2_51[29]}
   );
   gpc1_1 gpc4170 (
      {stage1_51[57]},
      {stage2_51[30]}
   );
   gpc1_1 gpc4171 (
      {stage1_51[58]},
      {stage2_51[31]}
   );
   gpc1_1 gpc4172 (
      {stage1_51[59]},
      {stage2_51[32]}
   );
   gpc1_1 gpc4173 (
      {stage1_51[60]},
      {stage2_51[33]}
   );
   gpc1_1 gpc4174 (
      {stage1_51[61]},
      {stage2_51[34]}
   );
   gpc1_1 gpc4175 (
      {stage1_51[62]},
      {stage2_51[35]}
   );
   gpc1_1 gpc4176 (
      {stage1_51[63]},
      {stage2_51[36]}
   );
   gpc1_1 gpc4177 (
      {stage1_51[64]},
      {stage2_51[37]}
   );
   gpc1_1 gpc4178 (
      {stage1_51[65]},
      {stage2_51[38]}
   );
   gpc1_1 gpc4179 (
      {stage1_51[66]},
      {stage2_51[39]}
   );
   gpc1_1 gpc4180 (
      {stage1_51[67]},
      {stage2_51[40]}
   );
   gpc1_1 gpc4181 (
      {stage1_51[68]},
      {stage2_51[41]}
   );
   gpc1_1 gpc4182 (
      {stage1_51[69]},
      {stage2_51[42]}
   );
   gpc1_1 gpc4183 (
      {stage1_51[70]},
      {stage2_51[43]}
   );
   gpc1_1 gpc4184 (
      {stage1_51[71]},
      {stage2_51[44]}
   );
   gpc1_1 gpc4185 (
      {stage1_51[72]},
      {stage2_51[45]}
   );
   gpc1_1 gpc4186 (
      {stage1_51[73]},
      {stage2_51[46]}
   );
   gpc1_1 gpc4187 (
      {stage1_51[74]},
      {stage2_51[47]}
   );
   gpc1_1 gpc4188 (
      {stage1_51[75]},
      {stage2_51[48]}
   );
   gpc1_1 gpc4189 (
      {stage1_51[76]},
      {stage2_51[49]}
   );
   gpc1_1 gpc4190 (
      {stage1_51[77]},
      {stage2_51[50]}
   );
   gpc1_1 gpc4191 (
      {stage1_51[78]},
      {stage2_51[51]}
   );
   gpc1_1 gpc4192 (
      {stage1_51[79]},
      {stage2_51[52]}
   );
   gpc1_1 gpc4193 (
      {stage1_51[80]},
      {stage2_51[53]}
   );
   gpc1_1 gpc4194 (
      {stage1_51[81]},
      {stage2_51[54]}
   );
   gpc1_1 gpc4195 (
      {stage1_51[82]},
      {stage2_51[55]}
   );
   gpc1_1 gpc4196 (
      {stage1_51[83]},
      {stage2_51[56]}
   );
   gpc1_1 gpc4197 (
      {stage1_51[84]},
      {stage2_51[57]}
   );
   gpc1_1 gpc4198 (
      {stage1_51[85]},
      {stage2_51[58]}
   );
   gpc1_1 gpc4199 (
      {stage1_51[86]},
      {stage2_51[59]}
   );
   gpc1_1 gpc4200 (
      {stage1_51[87]},
      {stage2_51[60]}
   );
   gpc1_1 gpc4201 (
      {stage1_51[88]},
      {stage2_51[61]}
   );
   gpc1_1 gpc4202 (
      {stage1_51[89]},
      {stage2_51[62]}
   );
   gpc1_1 gpc4203 (
      {stage1_51[90]},
      {stage2_51[63]}
   );
   gpc1_1 gpc4204 (
      {stage1_51[91]},
      {stage2_51[64]}
   );
   gpc1_1 gpc4205 (
      {stage1_51[92]},
      {stage2_51[65]}
   );
   gpc1_1 gpc4206 (
      {stage1_51[93]},
      {stage2_51[66]}
   );
   gpc1_1 gpc4207 (
      {stage1_51[94]},
      {stage2_51[67]}
   );
   gpc1_1 gpc4208 (
      {stage1_51[95]},
      {stage2_51[68]}
   );
   gpc1_1 gpc4209 (
      {stage1_51[96]},
      {stage2_51[69]}
   );
   gpc1_1 gpc4210 (
      {stage1_51[97]},
      {stage2_51[70]}
   );
   gpc1_1 gpc4211 (
      {stage1_51[98]},
      {stage2_51[71]}
   );
   gpc1_1 gpc4212 (
      {stage1_51[99]},
      {stage2_51[72]}
   );
   gpc1_1 gpc4213 (
      {stage1_51[100]},
      {stage2_51[73]}
   );
   gpc1_1 gpc4214 (
      {stage1_51[101]},
      {stage2_51[74]}
   );
   gpc1_1 gpc4215 (
      {stage1_51[102]},
      {stage2_51[75]}
   );
   gpc1_1 gpc4216 (
      {stage1_51[103]},
      {stage2_51[76]}
   );
   gpc1_1 gpc4217 (
      {stage1_51[104]},
      {stage2_51[77]}
   );
   gpc1_1 gpc4218 (
      {stage1_51[105]},
      {stage2_51[78]}
   );
   gpc1_1 gpc4219 (
      {stage1_52[116]},
      {stage2_52[27]}
   );
   gpc1_1 gpc4220 (
      {stage1_52[117]},
      {stage2_52[28]}
   );
   gpc1_1 gpc4221 (
      {stage1_52[118]},
      {stage2_52[29]}
   );
   gpc1_1 gpc4222 (
      {stage1_52[119]},
      {stage2_52[30]}
   );
   gpc1_1 gpc4223 (
      {stage1_52[120]},
      {stage2_52[31]}
   );
   gpc1_1 gpc4224 (
      {stage1_52[121]},
      {stage2_52[32]}
   );
   gpc1_1 gpc4225 (
      {stage1_52[122]},
      {stage2_52[33]}
   );
   gpc1_1 gpc4226 (
      {stage1_52[123]},
      {stage2_52[34]}
   );
   gpc1_1 gpc4227 (
      {stage1_52[124]},
      {stage2_52[35]}
   );
   gpc1_1 gpc4228 (
      {stage1_52[125]},
      {stage2_52[36]}
   );
   gpc1_1 gpc4229 (
      {stage1_52[126]},
      {stage2_52[37]}
   );
   gpc1_1 gpc4230 (
      {stage1_52[127]},
      {stage2_52[38]}
   );
   gpc1_1 gpc4231 (
      {stage1_52[128]},
      {stage2_52[39]}
   );
   gpc1_1 gpc4232 (
      {stage1_52[129]},
      {stage2_52[40]}
   );
   gpc1_1 gpc4233 (
      {stage1_52[130]},
      {stage2_52[41]}
   );
   gpc1_1 gpc4234 (
      {stage1_52[131]},
      {stage2_52[42]}
   );
   gpc1_1 gpc4235 (
      {stage1_52[132]},
      {stage2_52[43]}
   );
   gpc1_1 gpc4236 (
      {stage1_52[133]},
      {stage2_52[44]}
   );
   gpc1_1 gpc4237 (
      {stage1_52[134]},
      {stage2_52[45]}
   );
   gpc1_1 gpc4238 (
      {stage1_52[135]},
      {stage2_52[46]}
   );
   gpc1_1 gpc4239 (
      {stage1_52[136]},
      {stage2_52[47]}
   );
   gpc1_1 gpc4240 (
      {stage1_52[137]},
      {stage2_52[48]}
   );
   gpc1_1 gpc4241 (
      {stage1_52[138]},
      {stage2_52[49]}
   );
   gpc1_1 gpc4242 (
      {stage1_52[139]},
      {stage2_52[50]}
   );
   gpc1_1 gpc4243 (
      {stage1_53[70]},
      {stage2_53[40]}
   );
   gpc1_1 gpc4244 (
      {stage1_53[71]},
      {stage2_53[41]}
   );
   gpc1_1 gpc4245 (
      {stage1_53[72]},
      {stage2_53[42]}
   );
   gpc1_1 gpc4246 (
      {stage1_53[73]},
      {stage2_53[43]}
   );
   gpc1_1 gpc4247 (
      {stage1_53[74]},
      {stage2_53[44]}
   );
   gpc1_1 gpc4248 (
      {stage1_53[75]},
      {stage2_53[45]}
   );
   gpc1_1 gpc4249 (
      {stage1_53[76]},
      {stage2_53[46]}
   );
   gpc1_1 gpc4250 (
      {stage1_53[77]},
      {stage2_53[47]}
   );
   gpc1_1 gpc4251 (
      {stage1_53[78]},
      {stage2_53[48]}
   );
   gpc1_1 gpc4252 (
      {stage1_53[79]},
      {stage2_53[49]}
   );
   gpc1_1 gpc4253 (
      {stage1_53[80]},
      {stage2_53[50]}
   );
   gpc1_1 gpc4254 (
      {stage1_53[81]},
      {stage2_53[51]}
   );
   gpc1_1 gpc4255 (
      {stage1_53[82]},
      {stage2_53[52]}
   );
   gpc1_1 gpc4256 (
      {stage1_53[83]},
      {stage2_53[53]}
   );
   gpc1_1 gpc4257 (
      {stage1_53[84]},
      {stage2_53[54]}
   );
   gpc1_1 gpc4258 (
      {stage1_53[85]},
      {stage2_53[55]}
   );
   gpc1_1 gpc4259 (
      {stage1_53[86]},
      {stage2_53[56]}
   );
   gpc1_1 gpc4260 (
      {stage1_53[87]},
      {stage2_53[57]}
   );
   gpc1_1 gpc4261 (
      {stage1_53[88]},
      {stage2_53[58]}
   );
   gpc1_1 gpc4262 (
      {stage1_53[89]},
      {stage2_53[59]}
   );
   gpc1_1 gpc4263 (
      {stage1_53[90]},
      {stage2_53[60]}
   );
   gpc1_1 gpc4264 (
      {stage1_53[91]},
      {stage2_53[61]}
   );
   gpc1_1 gpc4265 (
      {stage1_53[92]},
      {stage2_53[62]}
   );
   gpc1_1 gpc4266 (
      {stage1_53[93]},
      {stage2_53[63]}
   );
   gpc1_1 gpc4267 (
      {stage1_53[94]},
      {stage2_53[64]}
   );
   gpc1_1 gpc4268 (
      {stage1_53[95]},
      {stage2_53[65]}
   );
   gpc1_1 gpc4269 (
      {stage1_53[96]},
      {stage2_53[66]}
   );
   gpc1_1 gpc4270 (
      {stage1_53[97]},
      {stage2_53[67]}
   );
   gpc1_1 gpc4271 (
      {stage1_53[98]},
      {stage2_53[68]}
   );
   gpc1_1 gpc4272 (
      {stage1_53[99]},
      {stage2_53[69]}
   );
   gpc1_1 gpc4273 (
      {stage1_53[100]},
      {stage2_53[70]}
   );
   gpc1_1 gpc4274 (
      {stage1_53[101]},
      {stage2_53[71]}
   );
   gpc1_1 gpc4275 (
      {stage1_53[102]},
      {stage2_53[72]}
   );
   gpc1_1 gpc4276 (
      {stage1_53[103]},
      {stage2_53[73]}
   );
   gpc1_1 gpc4277 (
      {stage1_53[104]},
      {stage2_53[74]}
   );
   gpc1_1 gpc4278 (
      {stage1_53[105]},
      {stage2_53[75]}
   );
   gpc1_1 gpc4279 (
      {stage1_53[106]},
      {stage2_53[76]}
   );
   gpc1_1 gpc4280 (
      {stage1_53[107]},
      {stage2_53[77]}
   );
   gpc1_1 gpc4281 (
      {stage1_54[133]},
      {stage2_54[48]}
   );
   gpc1_1 gpc4282 (
      {stage1_54[134]},
      {stage2_54[49]}
   );
   gpc1_1 gpc4283 (
      {stage1_54[135]},
      {stage2_54[50]}
   );
   gpc1_1 gpc4284 (
      {stage1_54[136]},
      {stage2_54[51]}
   );
   gpc1_1 gpc4285 (
      {stage1_54[137]},
      {stage2_54[52]}
   );
   gpc1_1 gpc4286 (
      {stage1_54[138]},
      {stage2_54[53]}
   );
   gpc1_1 gpc4287 (
      {stage1_54[139]},
      {stage2_54[54]}
   );
   gpc1_1 gpc4288 (
      {stage1_54[140]},
      {stage2_54[55]}
   );
   gpc1_1 gpc4289 (
      {stage1_54[141]},
      {stage2_54[56]}
   );
   gpc1_1 gpc4290 (
      {stage1_54[142]},
      {stage2_54[57]}
   );
   gpc1_1 gpc4291 (
      {stage1_54[143]},
      {stage2_54[58]}
   );
   gpc1_1 gpc4292 (
      {stage1_54[144]},
      {stage2_54[59]}
   );
   gpc1_1 gpc4293 (
      {stage1_54[145]},
      {stage2_54[60]}
   );
   gpc1_1 gpc4294 (
      {stage1_54[146]},
      {stage2_54[61]}
   );
   gpc1_1 gpc4295 (
      {stage1_54[147]},
      {stage2_54[62]}
   );
   gpc1_1 gpc4296 (
      {stage1_54[148]},
      {stage2_54[63]}
   );
   gpc1_1 gpc4297 (
      {stage1_54[149]},
      {stage2_54[64]}
   );
   gpc1_1 gpc4298 (
      {stage1_54[150]},
      {stage2_54[65]}
   );
   gpc1_1 gpc4299 (
      {stage1_54[151]},
      {stage2_54[66]}
   );
   gpc1_1 gpc4300 (
      {stage1_54[152]},
      {stage2_54[67]}
   );
   gpc1_1 gpc4301 (
      {stage1_54[153]},
      {stage2_54[68]}
   );
   gpc1_1 gpc4302 (
      {stage1_54[154]},
      {stage2_54[69]}
   );
   gpc1_1 gpc4303 (
      {stage1_54[155]},
      {stage2_54[70]}
   );
   gpc1_1 gpc4304 (
      {stage1_54[156]},
      {stage2_54[71]}
   );
   gpc1_1 gpc4305 (
      {stage1_54[157]},
      {stage2_54[72]}
   );
   gpc1_1 gpc4306 (
      {stage1_54[158]},
      {stage2_54[73]}
   );
   gpc1_1 gpc4307 (
      {stage1_54[159]},
      {stage2_54[74]}
   );
   gpc1_1 gpc4308 (
      {stage1_56[150]},
      {stage2_56[45]}
   );
   gpc1_1 gpc4309 (
      {stage1_56[151]},
      {stage2_56[46]}
   );
   gpc1_1 gpc4310 (
      {stage1_56[152]},
      {stage2_56[47]}
   );
   gpc1_1 gpc4311 (
      {stage1_56[153]},
      {stage2_56[48]}
   );
   gpc1_1 gpc4312 (
      {stage1_56[154]},
      {stage2_56[49]}
   );
   gpc1_1 gpc4313 (
      {stage1_56[155]},
      {stage2_56[50]}
   );
   gpc1_1 gpc4314 (
      {stage1_56[156]},
      {stage2_56[51]}
   );
   gpc1_1 gpc4315 (
      {stage1_56[157]},
      {stage2_56[52]}
   );
   gpc1_1 gpc4316 (
      {stage1_56[158]},
      {stage2_56[53]}
   );
   gpc1_1 gpc4317 (
      {stage1_56[159]},
      {stage2_56[54]}
   );
   gpc1_1 gpc4318 (
      {stage1_56[160]},
      {stage2_56[55]}
   );
   gpc1_1 gpc4319 (
      {stage1_56[161]},
      {stage2_56[56]}
   );
   gpc1_1 gpc4320 (
      {stage1_56[162]},
      {stage2_56[57]}
   );
   gpc1_1 gpc4321 (
      {stage1_56[163]},
      {stage2_56[58]}
   );
   gpc1_1 gpc4322 (
      {stage1_56[164]},
      {stage2_56[59]}
   );
   gpc1_1 gpc4323 (
      {stage1_56[165]},
      {stage2_56[60]}
   );
   gpc1_1 gpc4324 (
      {stage1_56[166]},
      {stage2_56[61]}
   );
   gpc1_1 gpc4325 (
      {stage1_56[167]},
      {stage2_56[62]}
   );
   gpc1_1 gpc4326 (
      {stage1_56[168]},
      {stage2_56[63]}
   );
   gpc1_1 gpc4327 (
      {stage1_56[169]},
      {stage2_56[64]}
   );
   gpc1_1 gpc4328 (
      {stage1_56[170]},
      {stage2_56[65]}
   );
   gpc1_1 gpc4329 (
      {stage1_56[171]},
      {stage2_56[66]}
   );
   gpc1_1 gpc4330 (
      {stage1_56[172]},
      {stage2_56[67]}
   );
   gpc1_1 gpc4331 (
      {stage1_56[173]},
      {stage2_56[68]}
   );
   gpc1_1 gpc4332 (
      {stage1_56[174]},
      {stage2_56[69]}
   );
   gpc1_1 gpc4333 (
      {stage1_56[175]},
      {stage2_56[70]}
   );
   gpc1_1 gpc4334 (
      {stage1_56[176]},
      {stage2_56[71]}
   );
   gpc1_1 gpc4335 (
      {stage1_56[177]},
      {stage2_56[72]}
   );
   gpc1_1 gpc4336 (
      {stage1_57[72]},
      {stage2_57[50]}
   );
   gpc1_1 gpc4337 (
      {stage1_57[73]},
      {stage2_57[51]}
   );
   gpc1_1 gpc4338 (
      {stage1_57[74]},
      {stage2_57[52]}
   );
   gpc1_1 gpc4339 (
      {stage1_57[75]},
      {stage2_57[53]}
   );
   gpc1_1 gpc4340 (
      {stage1_57[76]},
      {stage2_57[54]}
   );
   gpc1_1 gpc4341 (
      {stage1_57[77]},
      {stage2_57[55]}
   );
   gpc1_1 gpc4342 (
      {stage1_57[78]},
      {stage2_57[56]}
   );
   gpc1_1 gpc4343 (
      {stage1_57[79]},
      {stage2_57[57]}
   );
   gpc1_1 gpc4344 (
      {stage1_57[80]},
      {stage2_57[58]}
   );
   gpc1_1 gpc4345 (
      {stage1_57[81]},
      {stage2_57[59]}
   );
   gpc1_1 gpc4346 (
      {stage1_57[82]},
      {stage2_57[60]}
   );
   gpc1_1 gpc4347 (
      {stage1_57[83]},
      {stage2_57[61]}
   );
   gpc1_1 gpc4348 (
      {stage1_57[84]},
      {stage2_57[62]}
   );
   gpc1_1 gpc4349 (
      {stage1_57[85]},
      {stage2_57[63]}
   );
   gpc1_1 gpc4350 (
      {stage1_57[86]},
      {stage2_57[64]}
   );
   gpc1_1 gpc4351 (
      {stage1_57[87]},
      {stage2_57[65]}
   );
   gpc1_1 gpc4352 (
      {stage1_57[88]},
      {stage2_57[66]}
   );
   gpc1_1 gpc4353 (
      {stage1_57[89]},
      {stage2_57[67]}
   );
   gpc1_1 gpc4354 (
      {stage1_57[90]},
      {stage2_57[68]}
   );
   gpc1_1 gpc4355 (
      {stage1_57[91]},
      {stage2_57[69]}
   );
   gpc1_1 gpc4356 (
      {stage1_57[92]},
      {stage2_57[70]}
   );
   gpc1_1 gpc4357 (
      {stage1_57[93]},
      {stage2_57[71]}
   );
   gpc1_1 gpc4358 (
      {stage1_57[94]},
      {stage2_57[72]}
   );
   gpc1_1 gpc4359 (
      {stage1_57[95]},
      {stage2_57[73]}
   );
   gpc1_1 gpc4360 (
      {stage1_57[96]},
      {stage2_57[74]}
   );
   gpc1_1 gpc4361 (
      {stage1_57[97]},
      {stage2_57[75]}
   );
   gpc1_1 gpc4362 (
      {stage1_57[98]},
      {stage2_57[76]}
   );
   gpc1_1 gpc4363 (
      {stage1_57[99]},
      {stage2_57[77]}
   );
   gpc1_1 gpc4364 (
      {stage1_57[100]},
      {stage2_57[78]}
   );
   gpc1_1 gpc4365 (
      {stage1_57[101]},
      {stage2_57[79]}
   );
   gpc1_1 gpc4366 (
      {stage1_57[102]},
      {stage2_57[80]}
   );
   gpc1_1 gpc4367 (
      {stage1_57[103]},
      {stage2_57[81]}
   );
   gpc1_1 gpc4368 (
      {stage1_57[104]},
      {stage2_57[82]}
   );
   gpc1_1 gpc4369 (
      {stage1_58[78]},
      {stage2_58[40]}
   );
   gpc1_1 gpc4370 (
      {stage1_58[79]},
      {stage2_58[41]}
   );
   gpc1_1 gpc4371 (
      {stage1_58[80]},
      {stage2_58[42]}
   );
   gpc1_1 gpc4372 (
      {stage1_58[81]},
      {stage2_58[43]}
   );
   gpc1_1 gpc4373 (
      {stage1_58[82]},
      {stage2_58[44]}
   );
   gpc1_1 gpc4374 (
      {stage1_58[83]},
      {stage2_58[45]}
   );
   gpc1_1 gpc4375 (
      {stage1_58[84]},
      {stage2_58[46]}
   );
   gpc1_1 gpc4376 (
      {stage1_58[85]},
      {stage2_58[47]}
   );
   gpc1_1 gpc4377 (
      {stage1_59[138]},
      {stage2_59[38]}
   );
   gpc1_1 gpc4378 (
      {stage1_59[139]},
      {stage2_59[39]}
   );
   gpc1_1 gpc4379 (
      {stage1_59[140]},
      {stage2_59[40]}
   );
   gpc1_1 gpc4380 (
      {stage1_59[141]},
      {stage2_59[41]}
   );
   gpc1_1 gpc4381 (
      {stage1_59[142]},
      {stage2_59[42]}
   );
   gpc1_1 gpc4382 (
      {stage1_59[143]},
      {stage2_59[43]}
   );
   gpc1_1 gpc4383 (
      {stage1_59[144]},
      {stage2_59[44]}
   );
   gpc1_1 gpc4384 (
      {stage1_59[145]},
      {stage2_59[45]}
   );
   gpc1_1 gpc4385 (
      {stage1_59[146]},
      {stage2_59[46]}
   );
   gpc1_1 gpc4386 (
      {stage1_59[147]},
      {stage2_59[47]}
   );
   gpc1_1 gpc4387 (
      {stage1_60[138]},
      {stage2_60[59]}
   );
   gpc1_1 gpc4388 (
      {stage1_60[139]},
      {stage2_60[60]}
   );
   gpc1_1 gpc4389 (
      {stage1_60[140]},
      {stage2_60[61]}
   );
   gpc1_1 gpc4390 (
      {stage1_60[141]},
      {stage2_60[62]}
   );
   gpc1_1 gpc4391 (
      {stage1_61[102]},
      {stage2_61[50]}
   );
   gpc1_1 gpc4392 (
      {stage1_61[103]},
      {stage2_61[51]}
   );
   gpc1_1 gpc4393 (
      {stage1_61[104]},
      {stage2_61[52]}
   );
   gpc1_1 gpc4394 (
      {stage1_61[105]},
      {stage2_61[53]}
   );
   gpc1_1 gpc4395 (
      {stage1_61[106]},
      {stage2_61[54]}
   );
   gpc1_1 gpc4396 (
      {stage1_61[107]},
      {stage2_61[55]}
   );
   gpc1_1 gpc4397 (
      {stage1_61[108]},
      {stage2_61[56]}
   );
   gpc1_1 gpc4398 (
      {stage1_62[198]},
      {stage2_62[50]}
   );
   gpc1_1 gpc4399 (
      {stage1_62[199]},
      {stage2_62[51]}
   );
   gpc1_1 gpc4400 (
      {stage1_62[200]},
      {stage2_62[52]}
   );
   gpc1_1 gpc4401 (
      {stage1_63[48]},
      {stage2_63[54]}
   );
   gpc1_1 gpc4402 (
      {stage1_63[49]},
      {stage2_63[55]}
   );
   gpc1_1 gpc4403 (
      {stage1_63[50]},
      {stage2_63[56]}
   );
   gpc1_1 gpc4404 (
      {stage1_63[51]},
      {stage2_63[57]}
   );
   gpc1_1 gpc4405 (
      {stage1_63[52]},
      {stage2_63[58]}
   );
   gpc1_1 gpc4406 (
      {stage1_63[53]},
      {stage2_63[59]}
   );
   gpc1_1 gpc4407 (
      {stage1_63[54]},
      {stage2_63[60]}
   );
   gpc1_1 gpc4408 (
      {stage1_63[55]},
      {stage2_63[61]}
   );
   gpc1_1 gpc4409 (
      {stage1_63[56]},
      {stage2_63[62]}
   );
   gpc1_1 gpc4410 (
      {stage1_63[57]},
      {stage2_63[63]}
   );
   gpc1_1 gpc4411 (
      {stage1_63[58]},
      {stage2_63[64]}
   );
   gpc1_1 gpc4412 (
      {stage1_63[59]},
      {stage2_63[65]}
   );
   gpc1_1 gpc4413 (
      {stage1_63[60]},
      {stage2_63[66]}
   );
   gpc1_1 gpc4414 (
      {stage1_63[61]},
      {stage2_63[67]}
   );
   gpc1_1 gpc4415 (
      {stage1_63[62]},
      {stage2_63[68]}
   );
   gpc1_1 gpc4416 (
      {stage1_63[63]},
      {stage2_63[69]}
   );
   gpc1_1 gpc4417 (
      {stage1_63[64]},
      {stage2_63[70]}
   );
   gpc1_1 gpc4418 (
      {stage1_63[65]},
      {stage2_63[71]}
   );
   gpc1_1 gpc4419 (
      {stage1_63[66]},
      {stage2_63[72]}
   );
   gpc1_1 gpc4420 (
      {stage1_63[67]},
      {stage2_63[73]}
   );
   gpc1_1 gpc4421 (
      {stage1_63[68]},
      {stage2_63[74]}
   );
   gpc1_1 gpc4422 (
      {stage1_64[60]},
      {stage2_64[41]}
   );
   gpc1_1 gpc4423 (
      {stage1_64[61]},
      {stage2_64[42]}
   );
   gpc1_1 gpc4424 (
      {stage1_64[62]},
      {stage2_64[43]}
   );
   gpc1_1 gpc4425 (
      {stage1_64[63]},
      {stage2_64[44]}
   );
   gpc615_5 gpc4426 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc4427 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[1]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc4428 (
      {stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[2]},
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc4429 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19]},
      {stage2_1[3]},
      {stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc7_3 gpc4430 (
      {stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10]},
      {stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc4431 (
      {stage2_1[11], stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[4],stage3_3[5],stage3_2[5],stage3_1[5]}
   );
   gpc606_5 gpc4432 (
      {stage2_1[17], stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[5],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc4433 (
      {stage2_1[23], stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[2],stage3_4[6],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc4434 (
      {stage2_1[29], stage2_1[30], stage2_1[31], stage2_1[32], stage2_1[33], stage2_1[34]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[3],stage3_4[7],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc615_5 gpc4435 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28]},
      {stage2_3[24]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[4],stage3_4[8],stage3_3[9],stage3_2[9]}
   );
   gpc1163_5 gpc4436 (
      {stage2_3[25], stage2_3[26], stage2_3[27]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_5[0]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[1],stage3_5[5],stage3_4[9],stage3_3[10]}
   );
   gpc606_5 gpc4437 (
      {stage2_3[28], stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6]},
      {stage3_7[1],stage3_6[2],stage3_5[6],stage3_4[10],stage3_3[11]}
   );
   gpc606_5 gpc4438 (
      {stage2_3[34], stage2_3[35], stage2_3[36], stage2_3[37], stage2_3[38], stage2_3[39]},
      {stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12]},
      {stage3_7[2],stage3_6[3],stage3_5[7],stage3_4[11],stage3_3[12]}
   );
   gpc615_5 gpc4439 (
      {stage2_3[40], stage2_3[41], stage2_3[42], stage2_3[43], stage2_3[44]},
      {stage2_4[12]},
      {stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17], stage2_5[18]},
      {stage3_7[3],stage3_6[4],stage3_5[8],stage3_4[12],stage3_3[13]}
   );
   gpc615_5 gpc4440 (
      {stage2_3[45], stage2_3[46], stage2_3[47], stage2_3[48], stage2_3[49]},
      {stage2_4[13]},
      {stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23], stage2_5[24]},
      {stage3_7[4],stage3_6[5],stage3_5[9],stage3_4[13],stage3_3[14]}
   );
   gpc606_5 gpc4441 (
      {stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19]},
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5], stage2_6[6]},
      {stage3_8[0],stage3_7[5],stage3_6[6],stage3_5[10],stage3_4[14]}
   );
   gpc606_5 gpc4442 (
      {stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11], stage2_6[12]},
      {stage3_8[1],stage3_7[6],stage3_6[7],stage3_5[11],stage3_4[15]}
   );
   gpc606_5 gpc4443 (
      {stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29], stage2_4[30], stage2_4[31]},
      {stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17], stage2_6[18]},
      {stage3_8[2],stage3_7[7],stage3_6[8],stage3_5[12],stage3_4[16]}
   );
   gpc606_5 gpc4444 (
      {stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35], stage2_4[36], stage2_4[37]},
      {stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23], stage2_6[24]},
      {stage3_8[3],stage3_7[8],stage3_6[9],stage3_5[13],stage3_4[17]}
   );
   gpc615_5 gpc4445 (
      {stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41], stage2_4[42]},
      {stage2_5[25]},
      {stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29], stage2_6[30]},
      {stage3_8[4],stage3_7[9],stage3_6[10],stage3_5[14],stage3_4[18]}
   );
   gpc606_5 gpc4446 (
      {stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35], stage2_6[36]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[5],stage3_7[10],stage3_6[11]}
   );
   gpc606_5 gpc4447 (
      {stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41], stage2_6[42]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[6],stage3_7[11],stage3_6[12]}
   );
   gpc606_5 gpc4448 (
      {stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47], stage2_6[48]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[2],stage3_8[7],stage3_7[12],stage3_6[13]}
   );
   gpc615_5 gpc4449 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[18]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[3],stage3_9[3],stage3_8[8],stage3_7[13]}
   );
   gpc615_5 gpc4450 (
      {stage2_7[5], stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9]},
      {stage2_8[19]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[4],stage3_9[4],stage3_8[9],stage3_7[14]}
   );
   gpc615_5 gpc4451 (
      {stage2_7[10], stage2_7[11], stage2_7[12], stage2_7[13], stage2_7[14]},
      {stage2_8[20]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[5],stage3_9[5],stage3_8[10],stage3_7[15]}
   );
   gpc615_5 gpc4452 (
      {stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18], stage2_7[19]},
      {stage2_8[21]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[6],stage3_9[6],stage3_8[11],stage3_7[16]}
   );
   gpc615_5 gpc4453 (
      {stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24]},
      {stage2_8[22]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[7],stage3_9[7],stage3_8[12],stage3_7[17]}
   );
   gpc615_5 gpc4454 (
      {stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29]},
      {stage2_8[23]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[8],stage3_9[8],stage3_8[13],stage3_7[18]}
   );
   gpc615_5 gpc4455 (
      {stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34]},
      {stage2_8[24]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[9],stage3_9[9],stage3_8[14],stage3_7[19]}
   );
   gpc606_5 gpc4456 (
      {stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[7],stage3_10[10],stage3_9[10],stage3_8[15]}
   );
   gpc606_5 gpc4457 (
      {stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35], stage2_8[36]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[8],stage3_10[11],stage3_9[11],stage3_8[16]}
   );
   gpc606_5 gpc4458 (
      {stage2_8[37], stage2_8[38], stage2_8[39], stage2_8[40], stage2_8[41], stage2_8[42]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[9],stage3_10[12],stage3_9[12],stage3_8[17]}
   );
   gpc606_5 gpc4459 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[10],stage3_10[13],stage3_9[13]}
   );
   gpc606_5 gpc4460 (
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[4],stage3_11[11],stage3_10[14],stage3_9[14]}
   );
   gpc606_5 gpc4461 (
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[5],stage3_11[12],stage3_10[15],stage3_9[15]}
   );
   gpc606_5 gpc4462 (
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[3],stage3_12[6],stage3_11[13],stage3_10[16]}
   );
   gpc606_5 gpc4463 (
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[4],stage3_12[7],stage3_11[14],stage3_10[17]}
   );
   gpc606_5 gpc4464 (
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[5],stage3_12[8],stage3_11[15],stage3_10[18]}
   );
   gpc606_5 gpc4465 (
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage3_14[3],stage3_13[6],stage3_12[9],stage3_11[16],stage3_10[19]}
   );
   gpc606_5 gpc4466 (
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46], stage2_10[47]},
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage3_14[4],stage3_13[7],stage3_12[10],stage3_11[17],stage3_10[20]}
   );
   gpc606_5 gpc4467 (
      {stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51], stage2_10[52], stage2_10[53]},
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage3_14[5],stage3_13[8],stage3_12[11],stage3_11[18],stage3_10[21]}
   );
   gpc606_5 gpc4468 (
      {stage2_10[54], stage2_10[55], stage2_10[56], stage2_10[57], stage2_10[58], stage2_10[59]},
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage3_14[6],stage3_13[9],stage3_12[12],stage3_11[19],stage3_10[22]}
   );
   gpc615_5 gpc4469 (
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22]},
      {stage2_12[42]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[7],stage3_13[10],stage3_12[13],stage3_11[20]}
   );
   gpc615_5 gpc4470 (
      {stage2_11[23], stage2_11[24], stage2_11[25], stage2_11[26], stage2_11[27]},
      {stage2_12[43]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[8],stage3_13[11],stage3_12[14],stage3_11[21]}
   );
   gpc615_5 gpc4471 (
      {stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_12[44]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[9],stage3_13[12],stage3_12[15],stage3_11[22]}
   );
   gpc615_5 gpc4472 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37]},
      {stage2_12[45]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[10],stage3_13[13],stage3_12[16],stage3_11[23]}
   );
   gpc615_5 gpc4473 (
      {stage2_11[38], stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42]},
      {stage2_12[46]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[11],stage3_13[14],stage3_12[17],stage3_11[24]}
   );
   gpc606_5 gpc4474 (
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[0],stage3_15[5],stage3_14[12],stage3_13[15]}
   );
   gpc606_5 gpc4475 (
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[1],stage3_15[6],stage3_14[13],stage3_13[16]}
   );
   gpc606_5 gpc4476 (
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[2],stage3_15[7],stage3_14[14],stage3_13[17]}
   );
   gpc606_5 gpc4477 (
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[3],stage3_15[8],stage3_14[15],stage3_13[18]}
   );
   gpc606_5 gpc4478 (
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[4],stage3_15[9],stage3_14[16],stage3_13[19]}
   );
   gpc606_5 gpc4479 (
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[5],stage3_16[5],stage3_15[10],stage3_14[17]}
   );
   gpc606_5 gpc4480 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[6],stage3_16[6],stage3_15[11],stage3_14[18]}
   );
   gpc606_5 gpc4481 (
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[7],stage3_16[7],stage3_15[12],stage3_14[19]}
   );
   gpc606_5 gpc4482 (
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[8],stage3_16[8],stage3_15[13],stage3_14[20]}
   );
   gpc606_5 gpc4483 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[9],stage3_16[9],stage3_15[14],stage3_14[21]}
   );
   gpc606_5 gpc4484 (
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[10],stage3_16[10],stage3_15[15],stage3_14[22]}
   );
   gpc606_5 gpc4485 (
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[11],stage3_16[11],stage3_15[16],stage3_14[23]}
   );
   gpc615_5 gpc4486 (
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34]},
      {stage2_16[42]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[7],stage3_17[12],stage3_16[12],stage3_15[17]}
   );
   gpc615_5 gpc4487 (
      {stage2_15[35], stage2_15[36], stage2_15[37], stage2_15[38], stage2_15[39]},
      {stage2_16[43]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[8],stage3_17[13],stage3_16[13],stage3_15[18]}
   );
   gpc615_5 gpc4488 (
      {stage2_15[40], stage2_15[41], stage2_15[42], stage2_15[43], stage2_15[44]},
      {stage2_16[44]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[9],stage3_17[14],stage3_16[14],stage3_15[19]}
   );
   gpc615_5 gpc4489 (
      {stage2_15[45], stage2_15[46], stage2_15[47], stage2_15[48], stage2_15[49]},
      {stage2_16[45]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[10],stage3_17[15],stage3_16[15],stage3_15[20]}
   );
   gpc615_5 gpc4490 (
      {stage2_15[50], stage2_15[51], stage2_15[52], stage2_15[53], stage2_15[54]},
      {stage2_16[46]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[11],stage3_17[16],stage3_16[16],stage3_15[21]}
   );
   gpc606_5 gpc4491 (
      {stage2_16[47], stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[5],stage3_18[12],stage3_17[17],stage3_16[17]}
   );
   gpc606_5 gpc4492 (
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[6],stage3_18[13],stage3_17[18]}
   );
   gpc606_5 gpc4493 (
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], stage2_19[11]},
      {stage3_21[1],stage3_20[2],stage3_19[7],stage3_18[14],stage3_17[19]}
   );
   gpc606_5 gpc4494 (
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage2_19[12], stage2_19[13], stage2_19[14], stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage3_21[2],stage3_20[3],stage3_19[8],stage3_18[15],stage3_17[20]}
   );
   gpc615_5 gpc4495 (
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10]},
      {stage2_19[18]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[3],stage3_20[4],stage3_19[9],stage3_18[16]}
   );
   gpc615_5 gpc4496 (
      {stage2_18[11], stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15]},
      {stage2_19[19]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[4],stage3_20[5],stage3_19[10],stage3_18[17]}
   );
   gpc615_5 gpc4497 (
      {stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19], stage2_18[20]},
      {stage2_19[20]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[5],stage3_20[6],stage3_19[11],stage3_18[18]}
   );
   gpc615_5 gpc4498 (
      {stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24], stage2_18[25]},
      {stage2_19[21]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[6],stage3_20[7],stage3_19[12],stage3_18[19]}
   );
   gpc615_5 gpc4499 (
      {stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_19[22]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[7],stage3_20[8],stage3_19[13],stage3_18[20]}
   );
   gpc615_5 gpc4500 (
      {stage2_18[31], stage2_18[32], stage2_18[33], stage2_18[34], stage2_18[35]},
      {stage2_19[23]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[8],stage3_20[9],stage3_19[14],stage3_18[21]}
   );
   gpc615_5 gpc4501 (
      {stage2_18[36], stage2_18[37], stage2_18[38], stage2_18[39], stage2_18[40]},
      {stage2_19[24]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[9],stage3_20[10],stage3_19[15],stage3_18[22]}
   );
   gpc615_5 gpc4502 (
      {stage2_18[41], stage2_18[42], stage2_18[43], stage2_18[44], stage2_18[45]},
      {stage2_19[25]},
      {stage2_20[42], stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47]},
      {stage3_22[7],stage3_21[10],stage3_20[11],stage3_19[16],stage3_18[23]}
   );
   gpc615_5 gpc4503 (
      {stage2_18[46], stage2_18[47], stage2_18[48], stage2_18[49], stage2_18[50]},
      {stage2_19[26]},
      {stage2_20[48], stage2_20[49], stage2_20[50], stage2_20[51], stage2_20[52], stage2_20[53]},
      {stage3_22[8],stage3_21[11],stage3_20[12],stage3_19[17],stage3_18[24]}
   );
   gpc615_5 gpc4504 (
      {stage2_18[51], stage2_18[52], stage2_18[53], stage2_18[54], stage2_18[55]},
      {stage2_19[27]},
      {stage2_20[54], stage2_20[55], stage2_20[56], stage2_20[57], stage2_20[58], stage2_20[59]},
      {stage3_22[9],stage3_21[12],stage3_20[13],stage3_19[18],stage3_18[25]}
   );
   gpc615_5 gpc4505 (
      {stage2_18[56], stage2_18[57], stage2_18[58], stage2_18[59], stage2_18[60]},
      {stage2_19[28]},
      {stage2_20[60], stage2_20[61], stage2_20[62], stage2_20[63], stage2_20[64], stage2_20[65]},
      {stage3_22[10],stage3_21[13],stage3_20[14],stage3_19[19],stage3_18[26]}
   );
   gpc615_5 gpc4506 (
      {stage2_18[61], stage2_18[62], stage2_18[63], stage2_18[64], stage2_18[65]},
      {stage2_19[29]},
      {stage2_20[66], stage2_20[67], stage2_20[68], stage2_20[69], stage2_20[70], stage2_20[71]},
      {stage3_22[11],stage3_21[14],stage3_20[15],stage3_19[20],stage3_18[27]}
   );
   gpc606_5 gpc4507 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[12],stage3_21[15]}
   );
   gpc606_5 gpc4508 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[13],stage3_21[16]}
   );
   gpc606_5 gpc4509 (
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[14],stage3_21[17]}
   );
   gpc606_5 gpc4510 (
      {stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21], stage2_21[22], stage2_21[23]},
      {stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21], stage2_23[22], stage2_23[23]},
      {stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[15],stage3_21[18]}
   );
   gpc615_5 gpc4511 (
      {stage2_21[24], stage2_21[25], stage2_21[26], stage2_21[27], stage2_21[28]},
      {stage2_22[0]},
      {stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27], stage2_23[28], stage2_23[29]},
      {stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[16],stage3_21[19]}
   );
   gpc615_5 gpc4512 (
      {stage2_21[29], stage2_21[30], stage2_21[31], stage2_21[32], stage2_21[33]},
      {stage2_22[1]},
      {stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33], stage2_23[34], stage2_23[35]},
      {stage3_25[5],stage3_24[5],stage3_23[5],stage3_22[17],stage3_21[20]}
   );
   gpc615_5 gpc4513 (
      {stage2_21[34], stage2_21[35], stage2_21[36], stage2_21[37], stage2_21[38]},
      {stage2_22[2]},
      {stage2_23[36], stage2_23[37], stage2_23[38], stage2_23[39], stage2_23[40], stage2_23[41]},
      {stage3_25[6],stage3_24[6],stage3_23[6],stage3_22[18],stage3_21[21]}
   );
   gpc615_5 gpc4514 (
      {stage2_21[39], stage2_21[40], stage2_21[41], stage2_21[42], stage2_21[43]},
      {stage2_22[3]},
      {stage2_23[42], stage2_23[43], stage2_23[44], stage2_23[45], stage2_23[46], stage2_23[47]},
      {stage3_25[7],stage3_24[7],stage3_23[7],stage3_22[19],stage3_21[22]}
   );
   gpc615_5 gpc4515 (
      {stage2_21[44], stage2_21[45], stage2_21[46], stage2_21[47], stage2_21[48]},
      {stage2_22[4]},
      {stage2_23[48], stage2_23[49], stage2_23[50], stage2_23[51], stage2_23[52], stage2_23[53]},
      {stage3_25[8],stage3_24[8],stage3_23[8],stage3_22[20],stage3_21[23]}
   );
   gpc615_5 gpc4516 (
      {stage2_22[5], stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9]},
      {stage2_23[54]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[9],stage3_24[9],stage3_23[9],stage3_22[21]}
   );
   gpc615_5 gpc4517 (
      {stage2_22[10], stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14]},
      {stage2_23[55]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[10],stage3_24[10],stage3_23[10],stage3_22[22]}
   );
   gpc615_5 gpc4518 (
      {stage2_22[15], stage2_22[16], stage2_22[17], stage2_22[18], stage2_22[19]},
      {stage2_23[56]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[11],stage3_24[11],stage3_23[11],stage3_22[23]}
   );
   gpc615_5 gpc4519 (
      {stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23], stage2_22[24]},
      {stage2_23[57]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[12],stage3_24[12],stage3_23[12],stage3_22[24]}
   );
   gpc615_5 gpc4520 (
      {stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage2_23[58]},
      {stage2_24[24], stage2_24[25], stage2_24[26], stage2_24[27], stage2_24[28], stage2_24[29]},
      {stage3_26[4],stage3_25[13],stage3_24[13],stage3_23[13],stage3_22[25]}
   );
   gpc615_5 gpc4521 (
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34]},
      {stage2_23[59]},
      {stage2_24[30], stage2_24[31], stage2_24[32], stage2_24[33], stage2_24[34], stage2_24[35]},
      {stage3_26[5],stage3_25[14],stage3_24[14],stage3_23[14],stage3_22[26]}
   );
   gpc615_5 gpc4522 (
      {stage2_22[35], stage2_22[36], stage2_22[37], stage2_22[38], stage2_22[39]},
      {stage2_23[60]},
      {stage2_24[36], stage2_24[37], stage2_24[38], stage2_24[39], stage2_24[40], stage2_24[41]},
      {stage3_26[6],stage3_25[15],stage3_24[15],stage3_23[15],stage3_22[27]}
   );
   gpc606_5 gpc4523 (
      {stage2_24[42], stage2_24[43], stage2_24[44], stage2_24[45], stage2_24[46], stage2_24[47]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[0],stage3_26[7],stage3_25[16],stage3_24[16]}
   );
   gpc606_5 gpc4524 (
      {stage2_24[48], stage2_24[49], stage2_24[50], stage2_24[51], stage2_24[52], stage2_24[53]},
      {stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11]},
      {stage3_28[1],stage3_27[1],stage3_26[8],stage3_25[17],stage3_24[17]}
   );
   gpc606_5 gpc4525 (
      {stage2_24[54], stage2_24[55], stage2_24[56], stage2_24[57], stage2_24[58], stage2_24[59]},
      {stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17]},
      {stage3_28[2],stage3_27[2],stage3_26[9],stage3_25[18],stage3_24[18]}
   );
   gpc606_5 gpc4526 (
      {stage2_24[60], stage2_24[61], stage2_24[62], stage2_24[63], stage2_24[64], stage2_24[65]},
      {stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23]},
      {stage3_28[3],stage3_27[3],stage3_26[10],stage3_25[19],stage3_24[19]}
   );
   gpc606_5 gpc4527 (
      {stage2_24[66], stage2_24[67], stage2_24[68], stage2_24[69], stage2_24[70], stage2_24[71]},
      {stage2_26[24], stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29]},
      {stage3_28[4],stage3_27[4],stage3_26[11],stage3_25[20],stage3_24[20]}
   );
   gpc2135_5 gpc4528 (
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4]},
      {stage2_26[30], stage2_26[31], stage2_26[32]},
      {stage2_27[0]},
      {stage2_28[0], stage2_28[1]},
      {stage3_29[0],stage3_28[5],stage3_27[5],stage3_26[12],stage3_25[21]}
   );
   gpc606_5 gpc4529 (
      {stage2_25[5], stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10]},
      {stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5], stage2_27[6]},
      {stage3_29[1],stage3_28[6],stage3_27[6],stage3_26[13],stage3_25[22]}
   );
   gpc606_5 gpc4530 (
      {stage2_25[11], stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16]},
      {stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11], stage2_27[12]},
      {stage3_29[2],stage3_28[7],stage3_27[7],stage3_26[14],stage3_25[23]}
   );
   gpc606_5 gpc4531 (
      {stage2_25[17], stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22]},
      {stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17], stage2_27[18]},
      {stage3_29[3],stage3_28[8],stage3_27[8],stage3_26[15],stage3_25[24]}
   );
   gpc606_5 gpc4532 (
      {stage2_25[23], stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28]},
      {stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23], stage2_27[24]},
      {stage3_29[4],stage3_28[9],stage3_27[9],stage3_26[16],stage3_25[25]}
   );
   gpc606_5 gpc4533 (
      {stage2_25[29], stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34]},
      {stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30]},
      {stage3_29[5],stage3_28[10],stage3_27[10],stage3_26[17],stage3_25[26]}
   );
   gpc606_5 gpc4534 (
      {stage2_25[35], stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40]},
      {stage2_27[31], stage2_27[32], stage2_27[33], stage2_27[34], stage2_27[35], stage2_27[36]},
      {stage3_29[6],stage3_28[11],stage3_27[11],stage3_26[18],stage3_25[27]}
   );
   gpc615_5 gpc4535 (
      {stage2_25[41], stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45]},
      {stage2_26[33]},
      {stage2_27[37], stage2_27[38], stage2_27[39], stage2_27[40], stage2_27[41], stage2_27[42]},
      {stage3_29[7],stage3_28[12],stage3_27[12],stage3_26[19],stage3_25[28]}
   );
   gpc615_5 gpc4536 (
      {stage2_26[34], stage2_26[35], stage2_26[36], stage2_26[37], stage2_26[38]},
      {stage2_27[43]},
      {stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7]},
      {stage3_30[0],stage3_29[8],stage3_28[13],stage3_27[13],stage3_26[20]}
   );
   gpc615_5 gpc4537 (
      {stage2_26[39], stage2_26[40], stage2_26[41], stage2_26[42], stage2_26[43]},
      {stage2_27[44]},
      {stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage3_30[1],stage3_29[9],stage3_28[14],stage3_27[14],stage3_26[21]}
   );
   gpc615_5 gpc4538 (
      {stage2_26[44], stage2_26[45], stage2_26[46], stage2_26[47], stage2_26[48]},
      {stage2_27[45]},
      {stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18], stage2_28[19]},
      {stage3_30[2],stage3_29[10],stage3_28[15],stage3_27[15],stage3_26[22]}
   );
   gpc615_5 gpc4539 (
      {stage2_26[49], stage2_26[50], stage2_26[51], 1'b0, 1'b0},
      {stage2_27[46]},
      {stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23], stage2_28[24], stage2_28[25]},
      {stage3_30[3],stage3_29[11],stage3_28[16],stage3_27[16],stage3_26[23]}
   );
   gpc615_5 gpc4540 (
      {stage2_27[47], stage2_27[48], stage2_27[49], stage2_27[50], stage2_27[51]},
      {stage2_28[26]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[4],stage3_29[12],stage3_28[17],stage3_27[17]}
   );
   gpc615_5 gpc4541 (
      {stage2_27[52], stage2_27[53], stage2_27[54], stage2_27[55], stage2_27[56]},
      {stage2_28[27]},
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage3_31[1],stage3_30[5],stage3_29[13],stage3_28[18],stage3_27[18]}
   );
   gpc615_5 gpc4542 (
      {stage2_27[57], stage2_27[58], stage2_27[59], stage2_27[60], stage2_27[61]},
      {stage2_28[28]},
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage3_31[2],stage3_30[6],stage3_29[14],stage3_28[19],stage3_27[19]}
   );
   gpc615_5 gpc4543 (
      {stage2_27[62], stage2_27[63], stage2_27[64], stage2_27[65], stage2_27[66]},
      {stage2_28[29]},
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage3_31[3],stage3_30[7],stage3_29[15],stage3_28[20],stage3_27[20]}
   );
   gpc615_5 gpc4544 (
      {stage2_27[67], stage2_27[68], stage2_27[69], stage2_27[70], stage2_27[71]},
      {stage2_28[30]},
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage3_31[4],stage3_30[8],stage3_29[16],stage3_28[21],stage3_27[21]}
   );
   gpc606_5 gpc4545 (
      {stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34], stage2_28[35], stage2_28[36]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[5],stage3_30[9],stage3_29[17],stage3_28[22]}
   );
   gpc606_5 gpc4546 (
      {stage2_28[37], stage2_28[38], stage2_28[39], stage2_28[40], stage2_28[41], stage2_28[42]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[1],stage3_31[6],stage3_30[10],stage3_29[18],stage3_28[23]}
   );
   gpc606_5 gpc4547 (
      {stage2_28[43], stage2_28[44], stage2_28[45], stage2_28[46], stage2_28[47], stage2_28[48]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[2],stage3_31[7],stage3_30[11],stage3_29[19],stage3_28[24]}
   );
   gpc606_5 gpc4548 (
      {stage2_28[49], stage2_28[50], stage2_28[51], stage2_28[52], stage2_28[53], stage2_28[54]},
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22], stage2_30[23]},
      {stage3_32[3],stage3_31[8],stage3_30[12],stage3_29[20],stage3_28[25]}
   );
   gpc606_5 gpc4549 (
      {stage2_28[55], stage2_28[56], stage2_28[57], stage2_28[58], stage2_28[59], stage2_28[60]},
      {stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27], stage2_30[28], stage2_30[29]},
      {stage3_32[4],stage3_31[9],stage3_30[13],stage3_29[21],stage3_28[26]}
   );
   gpc606_5 gpc4550 (
      {stage2_28[61], stage2_28[62], stage2_28[63], stage2_28[64], stage2_28[65], stage2_28[66]},
      {stage2_30[30], stage2_30[31], stage2_30[32], stage2_30[33], stage2_30[34], stage2_30[35]},
      {stage3_32[5],stage3_31[10],stage3_30[14],stage3_29[22],stage3_28[27]}
   );
   gpc606_5 gpc4551 (
      {stage2_28[67], stage2_28[68], stage2_28[69], stage2_28[70], stage2_28[71], stage2_28[72]},
      {stage2_30[36], stage2_30[37], stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41]},
      {stage3_32[6],stage3_31[11],stage3_30[15],stage3_29[23],stage3_28[28]}
   );
   gpc606_5 gpc4552 (
      {stage2_29[30], stage2_29[31], stage2_29[32], stage2_29[33], stage2_29[34], stage2_29[35]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[7],stage3_31[12],stage3_30[16],stage3_29[24]}
   );
   gpc615_5 gpc4553 (
      {stage2_30[42], stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46]},
      {stage2_31[6]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[1],stage3_32[8],stage3_31[13],stage3_30[17]}
   );
   gpc615_5 gpc4554 (
      {stage2_30[47], stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51]},
      {stage2_31[7]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[2],stage3_32[9],stage3_31[14],stage3_30[18]}
   );
   gpc606_5 gpc4555 (
      {stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11], stage2_31[12], stage2_31[13]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[2],stage3_33[3],stage3_32[10],stage3_31[15]}
   );
   gpc606_5 gpc4556 (
      {stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17], stage2_31[18], stage2_31[19]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[3],stage3_33[4],stage3_32[11],stage3_31[16]}
   );
   gpc606_5 gpc4557 (
      {stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23], stage2_31[24], stage2_31[25]},
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16], stage2_33[17]},
      {stage3_35[2],stage3_34[4],stage3_33[5],stage3_32[12],stage3_31[17]}
   );
   gpc606_5 gpc4558 (
      {stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29], stage2_31[30], stage2_31[31]},
      {stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22], stage2_33[23]},
      {stage3_35[3],stage3_34[5],stage3_33[6],stage3_32[13],stage3_31[18]}
   );
   gpc606_5 gpc4559 (
      {stage2_31[32], stage2_31[33], stage2_31[34], stage2_31[35], stage2_31[36], stage2_31[37]},
      {stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28], stage2_33[29]},
      {stage3_35[4],stage3_34[6],stage3_33[7],stage3_32[14],stage3_31[19]}
   );
   gpc615_5 gpc4560 (
      {stage2_31[38], stage2_31[39], stage2_31[40], stage2_31[41], stage2_31[42]},
      {stage2_32[12]},
      {stage2_33[30], stage2_33[31], stage2_33[32], stage2_33[33], stage2_33[34], stage2_33[35]},
      {stage3_35[5],stage3_34[7],stage3_33[8],stage3_32[15],stage3_31[20]}
   );
   gpc117_4 gpc4561 (
      {stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17], stage2_32[18], stage2_32[19]},
      {stage2_33[36]},
      {stage2_34[0]},
      {stage3_35[6],stage3_34[8],stage3_33[9],stage3_32[16]}
   );
   gpc117_4 gpc4562 (
      {stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23], stage2_32[24], stage2_32[25], stage2_32[26]},
      {stage2_33[37]},
      {stage2_34[1]},
      {stage3_35[7],stage3_34[9],stage3_33[10],stage3_32[17]}
   );
   gpc606_5 gpc4563 (
      {stage2_32[27], stage2_32[28], stage2_32[29], stage2_32[30], stage2_32[31], stage2_32[32]},
      {stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5], stage2_34[6], stage2_34[7]},
      {stage3_36[0],stage3_35[8],stage3_34[10],stage3_33[11],stage3_32[18]}
   );
   gpc606_5 gpc4564 (
      {stage2_32[33], stage2_32[34], stage2_32[35], stage2_32[36], stage2_32[37], stage2_32[38]},
      {stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11], stage2_34[12], stage2_34[13]},
      {stage3_36[1],stage3_35[9],stage3_34[11],stage3_33[12],stage3_32[19]}
   );
   gpc615_5 gpc4565 (
      {stage2_34[14], stage2_34[15], stage2_34[16], stage2_34[17], stage2_34[18]},
      {stage2_35[0]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[0],stage3_36[2],stage3_35[10],stage3_34[12]}
   );
   gpc615_5 gpc4566 (
      {stage2_34[19], stage2_34[20], stage2_34[21], stage2_34[22], stage2_34[23]},
      {stage2_35[1]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[1],stage3_36[3],stage3_35[11],stage3_34[13]}
   );
   gpc615_5 gpc4567 (
      {stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5], stage2_35[6]},
      {stage2_36[12]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[2],stage3_37[2],stage3_36[4],stage3_35[12]}
   );
   gpc615_5 gpc4568 (
      {stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage2_36[13]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage3_39[1],stage3_38[3],stage3_37[3],stage3_36[5],stage3_35[13]}
   );
   gpc615_5 gpc4569 (
      {stage2_35[12], stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16]},
      {stage2_36[14]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage3_39[2],stage3_38[4],stage3_37[4],stage3_36[6],stage3_35[14]}
   );
   gpc615_5 gpc4570 (
      {stage2_35[17], stage2_35[18], stage2_35[19], stage2_35[20], stage2_35[21]},
      {stage2_36[15]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage3_39[3],stage3_38[5],stage3_37[5],stage3_36[7],stage3_35[15]}
   );
   gpc615_5 gpc4571 (
      {stage2_35[22], stage2_35[23], stage2_35[24], stage2_35[25], stage2_35[26]},
      {stage2_36[16]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage3_39[4],stage3_38[6],stage3_37[6],stage3_36[8],stage3_35[16]}
   );
   gpc615_5 gpc4572 (
      {stage2_35[27], stage2_35[28], stage2_35[29], stage2_35[30], stage2_35[31]},
      {stage2_36[17]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage3_39[5],stage3_38[7],stage3_37[7],stage3_36[9],stage3_35[17]}
   );
   gpc615_5 gpc4573 (
      {stage2_35[32], stage2_35[33], stage2_35[34], stage2_35[35], stage2_35[36]},
      {stage2_36[18]},
      {stage2_37[36], stage2_37[37], stage2_37[38], stage2_37[39], stage2_37[40], stage2_37[41]},
      {stage3_39[6],stage3_38[8],stage3_37[8],stage3_36[10],stage3_35[18]}
   );
   gpc615_5 gpc4574 (
      {stage2_35[37], stage2_35[38], stage2_35[39], stage2_35[40], stage2_35[41]},
      {stage2_36[19]},
      {stage2_37[42], stage2_37[43], stage2_37[44], stage2_37[45], stage2_37[46], stage2_37[47]},
      {stage3_39[7],stage3_38[9],stage3_37[9],stage3_36[11],stage3_35[19]}
   );
   gpc615_5 gpc4575 (
      {stage2_35[42], stage2_35[43], stage2_35[44], stage2_35[45], stage2_35[46]},
      {stage2_36[20]},
      {stage2_37[48], stage2_37[49], stage2_37[50], stage2_37[51], stage2_37[52], stage2_37[53]},
      {stage3_39[8],stage3_38[10],stage3_37[10],stage3_36[12],stage3_35[20]}
   );
   gpc606_5 gpc4576 (
      {stage2_36[21], stage2_36[22], stage2_36[23], stage2_36[24], stage2_36[25], stage2_36[26]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[9],stage3_38[11],stage3_37[11],stage3_36[13]}
   );
   gpc606_5 gpc4577 (
      {stage2_36[27], stage2_36[28], stage2_36[29], stage2_36[30], stage2_36[31], stage2_36[32]},
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11]},
      {stage3_40[1],stage3_39[10],stage3_38[12],stage3_37[12],stage3_36[14]}
   );
   gpc606_5 gpc4578 (
      {stage2_36[33], stage2_36[34], stage2_36[35], stage2_36[36], stage2_36[37], stage2_36[38]},
      {stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17]},
      {stage3_40[2],stage3_39[11],stage3_38[13],stage3_37[13],stage3_36[15]}
   );
   gpc606_5 gpc4579 (
      {stage2_36[39], stage2_36[40], stage2_36[41], stage2_36[42], stage2_36[43], stage2_36[44]},
      {stage2_38[18], stage2_38[19], stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23]},
      {stage3_40[3],stage3_39[12],stage3_38[14],stage3_37[14],stage3_36[16]}
   );
   gpc606_5 gpc4580 (
      {stage2_36[45], stage2_36[46], stage2_36[47], stage2_36[48], stage2_36[49], stage2_36[50]},
      {stage2_38[24], stage2_38[25], stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29]},
      {stage3_40[4],stage3_39[13],stage3_38[15],stage3_37[15],stage3_36[17]}
   );
   gpc606_5 gpc4581 (
      {stage2_36[51], stage2_36[52], stage2_36[53], stage2_36[54], stage2_36[55], stage2_36[56]},
      {stage2_38[30], stage2_38[31], stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35]},
      {stage3_40[5],stage3_39[14],stage3_38[16],stage3_37[16],stage3_36[18]}
   );
   gpc606_5 gpc4582 (
      {stage2_36[57], stage2_36[58], stage2_36[59], stage2_36[60], stage2_36[61], stage2_36[62]},
      {stage2_38[36], stage2_38[37], stage2_38[38], stage2_38[39], stage2_38[40], stage2_38[41]},
      {stage3_40[6],stage3_39[15],stage3_38[17],stage3_37[17],stage3_36[19]}
   );
   gpc2135_5 gpc4583 (
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4]},
      {stage2_40[0], stage2_40[1], stage2_40[2]},
      {stage2_41[0]},
      {stage2_42[0], stage2_42[1]},
      {stage3_43[0],stage3_42[0],stage3_41[0],stage3_40[7],stage3_39[16]}
   );
   gpc2135_5 gpc4584 (
      {stage2_39[5], stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9]},
      {stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage2_41[1]},
      {stage2_42[2], stage2_42[3]},
      {stage3_43[1],stage3_42[1],stage3_41[1],stage3_40[8],stage3_39[17]}
   );
   gpc2135_5 gpc4585 (
      {stage2_39[10], stage2_39[11], stage2_39[12], stage2_39[13], stage2_39[14]},
      {stage2_40[6], stage2_40[7], stage2_40[8]},
      {stage2_41[2]},
      {stage2_42[4], stage2_42[5]},
      {stage3_43[2],stage3_42[2],stage3_41[2],stage3_40[9],stage3_39[18]}
   );
   gpc2135_5 gpc4586 (
      {stage2_39[15], stage2_39[16], stage2_39[17], stage2_39[18], stage2_39[19]},
      {stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage2_41[3]},
      {stage2_42[6], stage2_42[7]},
      {stage3_43[3],stage3_42[3],stage3_41[3],stage3_40[10],stage3_39[19]}
   );
   gpc2135_5 gpc4587 (
      {stage2_39[20], stage2_39[21], stage2_39[22], stage2_39[23], stage2_39[24]},
      {stage2_40[12], stage2_40[13], stage2_40[14]},
      {stage2_41[4]},
      {stage2_42[8], stage2_42[9]},
      {stage3_43[4],stage3_42[4],stage3_41[4],stage3_40[11],stage3_39[20]}
   );
   gpc2135_5 gpc4588 (
      {stage2_39[25], stage2_39[26], stage2_39[27], stage2_39[28], stage2_39[29]},
      {stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage2_41[5]},
      {stage2_42[10], stage2_42[11]},
      {stage3_43[5],stage3_42[5],stage3_41[5],stage3_40[12],stage3_39[21]}
   );
   gpc2135_5 gpc4589 (
      {stage2_39[30], stage2_39[31], stage2_39[32], stage2_39[33], stage2_39[34]},
      {stage2_40[18], stage2_40[19], stage2_40[20]},
      {stage2_41[6]},
      {stage2_42[12], stage2_42[13]},
      {stage3_43[6],stage3_42[6],stage3_41[6],stage3_40[13],stage3_39[22]}
   );
   gpc2135_5 gpc4590 (
      {stage2_39[35], stage2_39[36], stage2_39[37], stage2_39[38], stage2_39[39]},
      {stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage2_41[7]},
      {stage2_42[14], stage2_42[15]},
      {stage3_43[7],stage3_42[7],stage3_41[7],stage3_40[14],stage3_39[23]}
   );
   gpc2135_5 gpc4591 (
      {stage2_39[40], stage2_39[41], stage2_39[42], stage2_39[43], stage2_39[44]},
      {stage2_40[24], stage2_40[25], stage2_40[26]},
      {stage2_41[8]},
      {stage2_42[16], stage2_42[17]},
      {stage3_43[8],stage3_42[8],stage3_41[8],stage3_40[15],stage3_39[24]}
   );
   gpc606_5 gpc4592 (
      {stage2_39[45], stage2_39[46], stage2_39[47], stage2_39[48], stage2_39[49], stage2_39[50]},
      {stage2_41[9], stage2_41[10], stage2_41[11], stage2_41[12], stage2_41[13], stage2_41[14]},
      {stage3_43[9],stage3_42[9],stage3_41[9],stage3_40[16],stage3_39[25]}
   );
   gpc606_5 gpc4593 (
      {stage2_39[51], stage2_39[52], stage2_39[53], stage2_39[54], stage2_39[55], stage2_39[56]},
      {stage2_41[15], stage2_41[16], stage2_41[17], stage2_41[18], stage2_41[19], stage2_41[20]},
      {stage3_43[10],stage3_42[10],stage3_41[10],stage3_40[17],stage3_39[26]}
   );
   gpc606_5 gpc4594 (
      {stage2_39[57], stage2_39[58], stage2_39[59], stage2_39[60], stage2_39[61], stage2_39[62]},
      {stage2_41[21], stage2_41[22], stage2_41[23], stage2_41[24], stage2_41[25], stage2_41[26]},
      {stage3_43[11],stage3_42[11],stage3_41[11],stage3_40[18],stage3_39[27]}
   );
   gpc606_5 gpc4595 (
      {stage2_39[63], stage2_39[64], stage2_39[65], stage2_39[66], stage2_39[67], stage2_39[68]},
      {stage2_41[27], stage2_41[28], stage2_41[29], stage2_41[30], stage2_41[31], stage2_41[32]},
      {stage3_43[12],stage3_42[12],stage3_41[12],stage3_40[19],stage3_39[28]}
   );
   gpc606_5 gpc4596 (
      {stage2_39[69], stage2_39[70], stage2_39[71], stage2_39[72], stage2_39[73], stage2_39[74]},
      {stage2_41[33], stage2_41[34], stage2_41[35], stage2_41[36], stage2_41[37], stage2_41[38]},
      {stage3_43[13],stage3_42[13],stage3_41[13],stage3_40[20],stage3_39[29]}
   );
   gpc606_5 gpc4597 (
      {stage2_39[75], stage2_39[76], stage2_39[77], stage2_39[78], stage2_39[79], stage2_39[80]},
      {stage2_41[39], stage2_41[40], stage2_41[41], stage2_41[42], stage2_41[43], stage2_41[44]},
      {stage3_43[14],stage3_42[14],stage3_41[14],stage3_40[21],stage3_39[30]}
   );
   gpc606_5 gpc4598 (
      {stage2_40[27], stage2_40[28], stage2_40[29], stage2_40[30], stage2_40[31], stage2_40[32]},
      {stage2_42[18], stage2_42[19], stage2_42[20], stage2_42[21], stage2_42[22], stage2_42[23]},
      {stage3_44[0],stage3_43[15],stage3_42[15],stage3_41[15],stage3_40[22]}
   );
   gpc606_5 gpc4599 (
      {stage2_40[33], stage2_40[34], stage2_40[35], stage2_40[36], stage2_40[37], stage2_40[38]},
      {stage2_42[24], stage2_42[25], stage2_42[26], stage2_42[27], stage2_42[28], stage2_42[29]},
      {stage3_44[1],stage3_43[16],stage3_42[16],stage3_41[16],stage3_40[23]}
   );
   gpc2135_5 gpc4600 (
      {stage2_41[45], stage2_41[46], stage2_41[47], stage2_41[48], stage2_41[49]},
      {stage2_42[30], stage2_42[31], stage2_42[32]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1]},
      {stage3_45[0],stage3_44[2],stage3_43[17],stage3_42[17],stage3_41[17]}
   );
   gpc1163_5 gpc4601 (
      {stage2_41[50], stage2_41[51], stage2_41[52]},
      {stage2_42[33], stage2_42[34], stage2_42[35], stage2_42[36], stage2_42[37], stage2_42[38]},
      {stage2_43[1]},
      {stage2_44[2]},
      {stage3_45[1],stage3_44[3],stage3_43[18],stage3_42[18],stage3_41[18]}
   );
   gpc1163_5 gpc4602 (
      {stage2_41[53], stage2_41[54], stage2_41[55]},
      {stage2_42[39], stage2_42[40], stage2_42[41], stage2_42[42], stage2_42[43], stage2_42[44]},
      {stage2_43[2]},
      {stage2_44[3]},
      {stage3_45[2],stage3_44[4],stage3_43[19],stage3_42[19],stage3_41[19]}
   );
   gpc1163_5 gpc4603 (
      {stage2_41[56], stage2_41[57], stage2_41[58]},
      {stage2_42[45], stage2_42[46], stage2_42[47], stage2_42[48], stage2_42[49], stage2_42[50]},
      {stage2_43[3]},
      {stage2_44[4]},
      {stage3_45[3],stage3_44[5],stage3_43[20],stage3_42[20],stage3_41[20]}
   );
   gpc606_5 gpc4604 (
      {stage2_41[59], stage2_41[60], stage2_41[61], stage2_41[62], stage2_41[63], stage2_41[64]},
      {stage2_43[4], stage2_43[5], stage2_43[6], stage2_43[7], stage2_43[8], stage2_43[9]},
      {stage3_45[4],stage3_44[6],stage3_43[21],stage3_42[21],stage3_41[21]}
   );
   gpc615_5 gpc4605 (
      {stage2_41[65], stage2_41[66], stage2_41[67], stage2_41[68], stage2_41[69]},
      {stage2_42[51]},
      {stage2_43[10], stage2_43[11], stage2_43[12], stage2_43[13], stage2_43[14], stage2_43[15]},
      {stage3_45[5],stage3_44[7],stage3_43[22],stage3_42[22],stage3_41[22]}
   );
   gpc615_5 gpc4606 (
      {stage2_41[70], stage2_41[71], stage2_41[72], stage2_41[73], stage2_41[74]},
      {stage2_42[52]},
      {stage2_43[16], stage2_43[17], stage2_43[18], stage2_43[19], stage2_43[20], stage2_43[21]},
      {stage3_45[6],stage3_44[8],stage3_43[23],stage3_42[23],stage3_41[23]}
   );
   gpc615_5 gpc4607 (
      {stage2_42[53], stage2_42[54], stage2_42[55], stage2_42[56], stage2_42[57]},
      {stage2_43[22]},
      {stage2_44[5], stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10]},
      {stage3_46[0],stage3_45[7],stage3_44[9],stage3_43[24],stage3_42[24]}
   );
   gpc606_5 gpc4608 (
      {stage2_43[23], stage2_43[24], stage2_43[25], stage2_43[26], stage2_43[27], stage2_43[28]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[1],stage3_45[8],stage3_44[10],stage3_43[25]}
   );
   gpc615_5 gpc4609 (
      {stage2_43[29], stage2_43[30], stage2_43[31], stage2_43[32], stage2_43[33]},
      {stage2_44[11]},
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage3_47[1],stage3_46[2],stage3_45[9],stage3_44[11],stage3_43[26]}
   );
   gpc615_5 gpc4610 (
      {stage2_43[34], stage2_43[35], stage2_43[36], stage2_43[37], stage2_43[38]},
      {stage2_44[12]},
      {stage2_45[12], stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage3_47[2],stage3_46[3],stage3_45[10],stage3_44[12],stage3_43[27]}
   );
   gpc615_5 gpc4611 (
      {stage2_43[39], stage2_43[40], stage2_43[41], stage2_43[42], stage2_43[43]},
      {stage2_44[13]},
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22], stage2_45[23]},
      {stage3_47[3],stage3_46[4],stage3_45[11],stage3_44[13],stage3_43[28]}
   );
   gpc615_5 gpc4612 (
      {stage2_43[44], stage2_43[45], stage2_43[46], stage2_43[47], stage2_43[48]},
      {stage2_44[14]},
      {stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27], stage2_45[28], stage2_45[29]},
      {stage3_47[4],stage3_46[5],stage3_45[12],stage3_44[14],stage3_43[29]}
   );
   gpc615_5 gpc4613 (
      {stage2_43[49], stage2_43[50], stage2_43[51], stage2_43[52], stage2_43[53]},
      {stage2_44[15]},
      {stage2_45[30], stage2_45[31], stage2_45[32], stage2_45[33], stage2_45[34], stage2_45[35]},
      {stage3_47[5],stage3_46[6],stage3_45[13],stage3_44[15],stage3_43[30]}
   );
   gpc606_5 gpc4614 (
      {stage2_44[16], stage2_44[17], stage2_44[18], stage2_44[19], stage2_44[20], stage2_44[21]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[6],stage3_46[7],stage3_45[14],stage3_44[16]}
   );
   gpc606_5 gpc4615 (
      {stage2_44[22], stage2_44[23], stage2_44[24], stage2_44[25], stage2_44[26], stage2_44[27]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[7],stage3_46[8],stage3_45[15],stage3_44[17]}
   );
   gpc606_5 gpc4616 (
      {stage2_44[28], stage2_44[29], stage2_44[30], stage2_44[31], stage2_44[32], stage2_44[33]},
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage3_48[2],stage3_47[8],stage3_46[9],stage3_45[16],stage3_44[18]}
   );
   gpc606_5 gpc4617 (
      {stage2_44[34], stage2_44[35], stage2_44[36], stage2_44[37], stage2_44[38], stage2_44[39]},
      {stage2_46[18], stage2_46[19], stage2_46[20], stage2_46[21], stage2_46[22], stage2_46[23]},
      {stage3_48[3],stage3_47[9],stage3_46[10],stage3_45[17],stage3_44[19]}
   );
   gpc606_5 gpc4618 (
      {stage2_44[40], stage2_44[41], stage2_44[42], stage2_44[43], stage2_44[44], stage2_44[45]},
      {stage2_46[24], stage2_46[25], stage2_46[26], stage2_46[27], stage2_46[28], stage2_46[29]},
      {stage3_48[4],stage3_47[10],stage3_46[11],stage3_45[18],stage3_44[20]}
   );
   gpc606_5 gpc4619 (
      {stage2_44[46], stage2_44[47], stage2_44[48], stage2_44[49], stage2_44[50], stage2_44[51]},
      {stage2_46[30], stage2_46[31], stage2_46[32], stage2_46[33], stage2_46[34], stage2_46[35]},
      {stage3_48[5],stage3_47[11],stage3_46[12],stage3_45[19],stage3_44[21]}
   );
   gpc615_5 gpc4620 (
      {stage2_45[36], stage2_45[37], stage2_45[38], stage2_45[39], stage2_45[40]},
      {stage2_46[36]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[6],stage3_47[12],stage3_46[13],stage3_45[20]}
   );
   gpc615_5 gpc4621 (
      {stage2_45[41], stage2_45[42], stage2_45[43], stage2_45[44], stage2_45[45]},
      {stage2_46[37]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[7],stage3_47[13],stage3_46[14],stage3_45[21]}
   );
   gpc615_5 gpc4622 (
      {stage2_45[46], stage2_45[47], stage2_45[48], stage2_45[49], stage2_45[50]},
      {stage2_46[38]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[8],stage3_47[14],stage3_46[15],stage3_45[22]}
   );
   gpc615_5 gpc4623 (
      {stage2_45[51], stage2_45[52], stage2_45[53], stage2_45[54], stage2_45[55]},
      {stage2_46[39]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[9],stage3_47[15],stage3_46[16],stage3_45[23]}
   );
   gpc615_5 gpc4624 (
      {stage2_45[56], stage2_45[57], stage2_45[58], stage2_45[59], stage2_45[60]},
      {stage2_46[40]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[10],stage3_47[16],stage3_46[17],stage3_45[24]}
   );
   gpc615_5 gpc4625 (
      {stage2_45[61], stage2_45[62], stage2_45[63], stage2_45[64], stage2_45[65]},
      {stage2_46[41]},
      {stage2_47[30], stage2_47[31], stage2_47[32], stage2_47[33], stage2_47[34], stage2_47[35]},
      {stage3_49[5],stage3_48[11],stage3_47[17],stage3_46[18],stage3_45[25]}
   );
   gpc615_5 gpc4626 (
      {stage2_47[36], stage2_47[37], stage2_47[38], stage2_47[39], stage2_47[40]},
      {stage2_48[0]},
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5]},
      {stage3_51[0],stage3_50[0],stage3_49[6],stage3_48[12],stage3_47[18]}
   );
   gpc615_5 gpc4627 (
      {stage2_47[41], stage2_47[42], stage2_47[43], stage2_47[44], stage2_47[45]},
      {stage2_48[1]},
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage3_51[1],stage3_50[1],stage3_49[7],stage3_48[13],stage3_47[19]}
   );
   gpc615_5 gpc4628 (
      {stage2_47[46], stage2_47[47], stage2_47[48], stage2_47[49], stage2_47[50]},
      {stage2_48[2]},
      {stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17]},
      {stage3_51[2],stage3_50[2],stage3_49[8],stage3_48[14],stage3_47[20]}
   );
   gpc615_5 gpc4629 (
      {stage2_47[51], stage2_47[52], stage2_47[53], stage2_47[54], stage2_47[55]},
      {stage2_48[3]},
      {stage2_49[18], stage2_49[19], stage2_49[20], stage2_49[21], stage2_49[22], stage2_49[23]},
      {stage3_51[3],stage3_50[3],stage3_49[9],stage3_48[15],stage3_47[21]}
   );
   gpc615_5 gpc4630 (
      {stage2_47[56], stage2_47[57], stage2_47[58], stage2_47[59], stage2_47[60]},
      {stage2_48[4]},
      {stage2_49[24], stage2_49[25], stage2_49[26], stage2_49[27], stage2_49[28], stage2_49[29]},
      {stage3_51[4],stage3_50[4],stage3_49[10],stage3_48[16],stage3_47[22]}
   );
   gpc606_5 gpc4631 (
      {stage2_48[5], stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10]},
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage3_52[0],stage3_51[5],stage3_50[5],stage3_49[11],stage3_48[17]}
   );
   gpc606_5 gpc4632 (
      {stage2_48[11], stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15], stage2_48[16]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[1],stage3_51[6],stage3_50[6],stage3_49[12],stage3_48[18]}
   );
   gpc615_5 gpc4633 (
      {stage2_48[17], stage2_48[18], stage2_48[19], stage2_48[20], stage2_48[21]},
      {stage2_49[30]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[2],stage3_51[7],stage3_50[7],stage3_49[13],stage3_48[19]}
   );
   gpc615_5 gpc4634 (
      {stage2_48[22], stage2_48[23], stage2_48[24], stage2_48[25], stage2_48[26]},
      {stage2_49[31]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[3],stage3_51[8],stage3_50[8],stage3_49[14],stage3_48[20]}
   );
   gpc615_5 gpc4635 (
      {stage2_48[27], stage2_48[28], stage2_48[29], stage2_48[30], stage2_48[31]},
      {stage2_49[32]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[4],stage3_51[9],stage3_50[9],stage3_49[15],stage3_48[21]}
   );
   gpc615_5 gpc4636 (
      {stage2_48[32], stage2_48[33], stage2_48[34], stage2_48[35], stage2_48[36]},
      {stage2_49[33]},
      {stage2_50[30], stage2_50[31], stage2_50[32], stage2_50[33], stage2_50[34], stage2_50[35]},
      {stage3_52[5],stage3_51[10],stage3_50[10],stage3_49[16],stage3_48[22]}
   );
   gpc615_5 gpc4637 (
      {stage2_48[37], stage2_48[38], stage2_48[39], stage2_48[40], stage2_48[41]},
      {stage2_49[34]},
      {stage2_50[36], stage2_50[37], stage2_50[38], stage2_50[39], stage2_50[40], stage2_50[41]},
      {stage3_52[6],stage3_51[11],stage3_50[11],stage3_49[17],stage3_48[23]}
   );
   gpc117_4 gpc4638 (
      {stage2_49[35], stage2_49[36], stage2_49[37], stage2_49[38], stage2_49[39], stage2_49[40], stage2_49[41]},
      {stage2_50[42]},
      {stage2_51[0]},
      {stage3_52[7],stage3_51[12],stage3_50[12],stage3_49[18]}
   );
   gpc117_4 gpc4639 (
      {stage2_49[42], stage2_49[43], stage2_49[44], stage2_49[45], stage2_49[46], stage2_49[47], stage2_49[48]},
      {stage2_50[43]},
      {stage2_51[1]},
      {stage3_52[8],stage3_51[13],stage3_50[13],stage3_49[19]}
   );
   gpc117_4 gpc4640 (
      {stage2_49[49], stage2_49[50], stage2_49[51], stage2_49[52], stage2_49[53], stage2_49[54], stage2_49[55]},
      {stage2_50[44]},
      {stage2_51[2]},
      {stage3_52[9],stage3_51[14],stage3_50[14],stage3_49[20]}
   );
   gpc117_4 gpc4641 (
      {stage2_49[56], stage2_49[57], stage2_49[58], stage2_49[59], stage2_49[60], stage2_49[61], stage2_49[62]},
      {stage2_50[45]},
      {stage2_51[3]},
      {stage3_52[10],stage3_51[15],stage3_50[15],stage3_49[21]}
   );
   gpc117_4 gpc4642 (
      {stage2_49[63], stage2_49[64], stage2_49[65], stage2_49[66], stage2_49[67], stage2_49[68], stage2_49[69]},
      {stage2_50[46]},
      {stage2_51[4]},
      {stage3_52[11],stage3_51[16],stage3_50[16],stage3_49[22]}
   );
   gpc615_5 gpc4643 (
      {stage2_50[47], stage2_50[48], stage2_50[49], stage2_50[50], stage2_50[51]},
      {stage2_51[5]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[0],stage3_52[12],stage3_51[17],stage3_50[17]}
   );
   gpc615_5 gpc4644 (
      {stage2_50[52], stage2_50[53], stage2_50[54], stage2_50[55], stage2_50[56]},
      {stage2_51[6]},
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11]},
      {stage3_54[1],stage3_53[1],stage3_52[13],stage3_51[18],stage3_50[18]}
   );
   gpc606_5 gpc4645 (
      {stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11], stage2_51[12]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[2],stage3_53[2],stage3_52[14],stage3_51[19]}
   );
   gpc606_5 gpc4646 (
      {stage2_51[13], stage2_51[14], stage2_51[15], stage2_51[16], stage2_51[17], stage2_51[18]},
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage3_55[1],stage3_54[3],stage3_53[3],stage3_52[15],stage3_51[20]}
   );
   gpc606_5 gpc4647 (
      {stage2_51[19], stage2_51[20], stage2_51[21], stage2_51[22], stage2_51[23], stage2_51[24]},
      {stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage3_55[2],stage3_54[4],stage3_53[4],stage3_52[16],stage3_51[21]}
   );
   gpc606_5 gpc4648 (
      {stage2_51[25], stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29], stage2_51[30]},
      {stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22], stage2_53[23]},
      {stage3_55[3],stage3_54[5],stage3_53[5],stage3_52[17],stage3_51[22]}
   );
   gpc606_5 gpc4649 (
      {stage2_51[31], stage2_51[32], stage2_51[33], stage2_51[34], stage2_51[35], stage2_51[36]},
      {stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28], stage2_53[29]},
      {stage3_55[4],stage3_54[6],stage3_53[6],stage3_52[18],stage3_51[23]}
   );
   gpc615_5 gpc4650 (
      {stage2_51[37], stage2_51[38], stage2_51[39], stage2_51[40], stage2_51[41]},
      {stage2_52[12]},
      {stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34], stage2_53[35]},
      {stage3_55[5],stage3_54[7],stage3_53[7],stage3_52[19],stage3_51[24]}
   );
   gpc615_5 gpc4651 (
      {stage2_51[42], stage2_51[43], stage2_51[44], stage2_51[45], stage2_51[46]},
      {stage2_52[13]},
      {stage2_53[36], stage2_53[37], stage2_53[38], stage2_53[39], stage2_53[40], stage2_53[41]},
      {stage3_55[6],stage3_54[8],stage3_53[8],stage3_52[20],stage3_51[25]}
   );
   gpc615_5 gpc4652 (
      {stage2_51[47], stage2_51[48], stage2_51[49], stage2_51[50], stage2_51[51]},
      {stage2_52[14]},
      {stage2_53[42], stage2_53[43], stage2_53[44], stage2_53[45], stage2_53[46], stage2_53[47]},
      {stage3_55[7],stage3_54[9],stage3_53[9],stage3_52[21],stage3_51[26]}
   );
   gpc623_5 gpc4653 (
      {stage2_51[52], stage2_51[53], stage2_51[54]},
      {stage2_52[15], stage2_52[16]},
      {stage2_53[48], stage2_53[49], stage2_53[50], stage2_53[51], stage2_53[52], stage2_53[53]},
      {stage3_55[8],stage3_54[10],stage3_53[10],stage3_52[22],stage3_51[27]}
   );
   gpc623_5 gpc4654 (
      {stage2_51[55], stage2_51[56], stage2_51[57]},
      {stage2_52[17], stage2_52[18]},
      {stage2_53[54], stage2_53[55], stage2_53[56], stage2_53[57], stage2_53[58], stage2_53[59]},
      {stage3_55[9],stage3_54[11],stage3_53[11],stage3_52[23],stage3_51[28]}
   );
   gpc623_5 gpc4655 (
      {stage2_51[58], stage2_51[59], stage2_51[60]},
      {stage2_52[19], stage2_52[20]},
      {stage2_53[60], stage2_53[61], stage2_53[62], stage2_53[63], stage2_53[64], stage2_53[65]},
      {stage3_55[10],stage3_54[12],stage3_53[12],stage3_52[24],stage3_51[29]}
   );
   gpc606_5 gpc4656 (
      {stage2_52[21], stage2_52[22], stage2_52[23], stage2_52[24], stage2_52[25], stage2_52[26]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[11],stage3_54[13],stage3_53[13],stage3_52[25]}
   );
   gpc606_5 gpc4657 (
      {stage2_52[27], stage2_52[28], stage2_52[29], stage2_52[30], stage2_52[31], stage2_52[32]},
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage3_56[1],stage3_55[12],stage3_54[14],stage3_53[14],stage3_52[26]}
   );
   gpc606_5 gpc4658 (
      {stage2_52[33], stage2_52[34], stage2_52[35], stage2_52[36], stage2_52[37], stage2_52[38]},
      {stage2_54[12], stage2_54[13], stage2_54[14], stage2_54[15], stage2_54[16], stage2_54[17]},
      {stage3_56[2],stage3_55[13],stage3_54[15],stage3_53[15],stage3_52[27]}
   );
   gpc606_5 gpc4659 (
      {stage2_54[18], stage2_54[19], stage2_54[20], stage2_54[21], stage2_54[22], stage2_54[23]},
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5]},
      {stage3_58[0],stage3_57[0],stage3_56[3],stage3_55[14],stage3_54[16]}
   );
   gpc606_5 gpc4660 (
      {stage2_54[24], stage2_54[25], stage2_54[26], stage2_54[27], stage2_54[28], stage2_54[29]},
      {stage2_56[6], stage2_56[7], stage2_56[8], stage2_56[9], stage2_56[10], stage2_56[11]},
      {stage3_58[1],stage3_57[1],stage3_56[4],stage3_55[15],stage3_54[17]}
   );
   gpc606_5 gpc4661 (
      {stage2_54[30], stage2_54[31], stage2_54[32], stage2_54[33], stage2_54[34], stage2_54[35]},
      {stage2_56[12], stage2_56[13], stage2_56[14], stage2_56[15], stage2_56[16], stage2_56[17]},
      {stage3_58[2],stage3_57[2],stage3_56[5],stage3_55[16],stage3_54[18]}
   );
   gpc606_5 gpc4662 (
      {stage2_54[36], stage2_54[37], stage2_54[38], stage2_54[39], stage2_54[40], stage2_54[41]},
      {stage2_56[18], stage2_56[19], stage2_56[20], stage2_56[21], stage2_56[22], stage2_56[23]},
      {stage3_58[3],stage3_57[3],stage3_56[6],stage3_55[17],stage3_54[19]}
   );
   gpc606_5 gpc4663 (
      {stage2_54[42], stage2_54[43], stage2_54[44], stage2_54[45], stage2_54[46], stage2_54[47]},
      {stage2_56[24], stage2_56[25], stage2_56[26], stage2_56[27], stage2_56[28], stage2_56[29]},
      {stage3_58[4],stage3_57[4],stage3_56[7],stage3_55[18],stage3_54[20]}
   );
   gpc606_5 gpc4664 (
      {stage2_54[48], stage2_54[49], stage2_54[50], stage2_54[51], stage2_54[52], stage2_54[53]},
      {stage2_56[30], stage2_56[31], stage2_56[32], stage2_56[33], stage2_56[34], stage2_56[35]},
      {stage3_58[5],stage3_57[5],stage3_56[8],stage3_55[19],stage3_54[21]}
   );
   gpc606_5 gpc4665 (
      {stage2_54[54], stage2_54[55], stage2_54[56], stage2_54[57], stage2_54[58], stage2_54[59]},
      {stage2_56[36], stage2_56[37], stage2_56[38], stage2_56[39], stage2_56[40], stage2_56[41]},
      {stage3_58[6],stage3_57[6],stage3_56[9],stage3_55[20],stage3_54[22]}
   );
   gpc606_5 gpc4666 (
      {stage2_54[60], stage2_54[61], stage2_54[62], stage2_54[63], stage2_54[64], stage2_54[65]},
      {stage2_56[42], stage2_56[43], stage2_56[44], stage2_56[45], stage2_56[46], stage2_56[47]},
      {stage3_58[7],stage3_57[7],stage3_56[10],stage3_55[21],stage3_54[23]}
   );
   gpc606_5 gpc4667 (
      {stage2_54[66], stage2_54[67], stage2_54[68], stage2_54[69], stage2_54[70], stage2_54[71]},
      {stage2_56[48], stage2_56[49], stage2_56[50], stage2_56[51], stage2_56[52], stage2_56[53]},
      {stage3_58[8],stage3_57[8],stage3_56[11],stage3_55[22],stage3_54[24]}
   );
   gpc615_5 gpc4668 (
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4]},
      {stage2_56[54]},
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4], stage2_57[5]},
      {stage3_59[0],stage3_58[9],stage3_57[9],stage3_56[12],stage3_55[23]}
   );
   gpc615_5 gpc4669 (
      {stage2_55[5], stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9]},
      {stage2_56[55]},
      {stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9], stage2_57[10], stage2_57[11]},
      {stage3_59[1],stage3_58[10],stage3_57[10],stage3_56[13],stage3_55[24]}
   );
   gpc615_5 gpc4670 (
      {stage2_55[10], stage2_55[11], stage2_55[12], stage2_55[13], stage2_55[14]},
      {stage2_56[56]},
      {stage2_57[12], stage2_57[13], stage2_57[14], stage2_57[15], stage2_57[16], stage2_57[17]},
      {stage3_59[2],stage3_58[11],stage3_57[11],stage3_56[14],stage3_55[25]}
   );
   gpc615_5 gpc4671 (
      {stage2_55[15], stage2_55[16], stage2_55[17], stage2_55[18], stage2_55[19]},
      {stage2_56[57]},
      {stage2_57[18], stage2_57[19], stage2_57[20], stage2_57[21], stage2_57[22], stage2_57[23]},
      {stage3_59[3],stage3_58[12],stage3_57[12],stage3_56[15],stage3_55[26]}
   );
   gpc615_5 gpc4672 (
      {stage2_55[20], stage2_55[21], stage2_55[22], stage2_55[23], stage2_55[24]},
      {stage2_56[58]},
      {stage2_57[24], stage2_57[25], stage2_57[26], stage2_57[27], stage2_57[28], stage2_57[29]},
      {stage3_59[4],stage3_58[13],stage3_57[13],stage3_56[16],stage3_55[27]}
   );
   gpc615_5 gpc4673 (
      {stage2_55[25], stage2_55[26], stage2_55[27], stage2_55[28], stage2_55[29]},
      {stage2_56[59]},
      {stage2_57[30], stage2_57[31], stage2_57[32], stage2_57[33], stage2_57[34], stage2_57[35]},
      {stage3_59[5],stage3_58[14],stage3_57[14],stage3_56[17],stage3_55[28]}
   );
   gpc615_5 gpc4674 (
      {stage2_55[30], stage2_55[31], stage2_55[32], stage2_55[33], stage2_55[34]},
      {stage2_56[60]},
      {stage2_57[36], stage2_57[37], stage2_57[38], stage2_57[39], stage2_57[40], stage2_57[41]},
      {stage3_59[6],stage3_58[15],stage3_57[15],stage3_56[18],stage3_55[29]}
   );
   gpc606_5 gpc4675 (
      {stage2_56[61], stage2_56[62], stage2_56[63], stage2_56[64], stage2_56[65], stage2_56[66]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[7],stage3_58[16],stage3_57[16],stage3_56[19]}
   );
   gpc606_5 gpc4676 (
      {stage2_57[42], stage2_57[43], stage2_57[44], stage2_57[45], stage2_57[46], stage2_57[47]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[1],stage3_59[8],stage3_58[17],stage3_57[17]}
   );
   gpc606_5 gpc4677 (
      {stage2_57[48], stage2_57[49], stage2_57[50], stage2_57[51], stage2_57[52], stage2_57[53]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[2],stage3_59[9],stage3_58[18],stage3_57[18]}
   );
   gpc606_5 gpc4678 (
      {stage2_57[54], stage2_57[55], stage2_57[56], stage2_57[57], stage2_57[58], stage2_57[59]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage3_61[2],stage3_60[3],stage3_59[10],stage3_58[19],stage3_57[19]}
   );
   gpc606_5 gpc4679 (
      {stage2_57[60], stage2_57[61], stage2_57[62], stage2_57[63], stage2_57[64], stage2_57[65]},
      {stage2_59[18], stage2_59[19], stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23]},
      {stage3_61[3],stage3_60[4],stage3_59[11],stage3_58[20],stage3_57[20]}
   );
   gpc606_5 gpc4680 (
      {stage2_57[66], stage2_57[67], stage2_57[68], stage2_57[69], stage2_57[70], stage2_57[71]},
      {stage2_59[24], stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29]},
      {stage3_61[4],stage3_60[5],stage3_59[12],stage3_58[21],stage3_57[21]}
   );
   gpc606_5 gpc4681 (
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage2_60[0], stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage3_62[0],stage3_61[5],stage3_60[6],stage3_59[13],stage3_58[22]}
   );
   gpc606_5 gpc4682 (
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage2_60[6], stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11]},
      {stage3_62[1],stage3_61[6],stage3_60[7],stage3_59[14],stage3_58[23]}
   );
   gpc606_5 gpc4683 (
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23]},
      {stage2_60[12], stage2_60[13], stage2_60[14], stage2_60[15], stage2_60[16], stage2_60[17]},
      {stage3_62[2],stage3_61[7],stage3_60[8],stage3_59[15],stage3_58[24]}
   );
   gpc606_5 gpc4684 (
      {stage2_58[24], stage2_58[25], stage2_58[26], stage2_58[27], stage2_58[28], stage2_58[29]},
      {stage2_60[18], stage2_60[19], stage2_60[20], stage2_60[21], stage2_60[22], stage2_60[23]},
      {stage3_62[3],stage3_61[8],stage3_60[9],stage3_59[16],stage3_58[25]}
   );
   gpc606_5 gpc4685 (
      {stage2_58[30], stage2_58[31], stage2_58[32], stage2_58[33], stage2_58[34], stage2_58[35]},
      {stage2_60[24], stage2_60[25], stage2_60[26], stage2_60[27], stage2_60[28], stage2_60[29]},
      {stage3_62[4],stage3_61[9],stage3_60[10],stage3_59[17],stage3_58[26]}
   );
   gpc606_5 gpc4686 (
      {stage2_58[36], stage2_58[37], stage2_58[38], stage2_58[39], stage2_58[40], stage2_58[41]},
      {stage2_60[30], stage2_60[31], stage2_60[32], stage2_60[33], stage2_60[34], stage2_60[35]},
      {stage3_62[5],stage3_61[10],stage3_60[11],stage3_59[18],stage3_58[27]}
   );
   gpc606_5 gpc4687 (
      {stage2_58[42], stage2_58[43], stage2_58[44], stage2_58[45], stage2_58[46], stage2_58[47]},
      {stage2_60[36], stage2_60[37], stage2_60[38], stage2_60[39], stage2_60[40], stage2_60[41]},
      {stage3_62[6],stage3_61[11],stage3_60[12],stage3_59[19],stage3_58[28]}
   );
   gpc606_5 gpc4688 (
      {stage2_59[30], stage2_59[31], stage2_59[32], stage2_59[33], stage2_59[34], stage2_59[35]},
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage3_63[0],stage3_62[7],stage3_61[12],stage3_60[13],stage3_59[20]}
   );
   gpc606_5 gpc4689 (
      {stage2_61[6], stage2_61[7], stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[0],stage3_63[1],stage3_62[8],stage3_61[13]}
   );
   gpc606_5 gpc4690 (
      {stage2_61[12], stage2_61[13], stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17]},
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage3_65[1],stage3_64[1],stage3_63[2],stage3_62[9],stage3_61[14]}
   );
   gpc606_5 gpc4691 (
      {stage2_61[18], stage2_61[19], stage2_61[20], stage2_61[21], stage2_61[22], stage2_61[23]},
      {stage2_63[12], stage2_63[13], stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17]},
      {stage3_65[2],stage3_64[2],stage3_63[3],stage3_62[10],stage3_61[15]}
   );
   gpc606_5 gpc4692 (
      {stage2_61[24], stage2_61[25], stage2_61[26], stage2_61[27], stage2_61[28], stage2_61[29]},
      {stage2_63[18], stage2_63[19], stage2_63[20], stage2_63[21], stage2_63[22], stage2_63[23]},
      {stage3_65[3],stage3_64[3],stage3_63[4],stage3_62[11],stage3_61[16]}
   );
   gpc606_5 gpc4693 (
      {stage2_61[30], stage2_61[31], stage2_61[32], stage2_61[33], stage2_61[34], stage2_61[35]},
      {stage2_63[24], stage2_63[25], stage2_63[26], stage2_63[27], stage2_63[28], stage2_63[29]},
      {stage3_65[4],stage3_64[4],stage3_63[5],stage3_62[12],stage3_61[17]}
   );
   gpc606_5 gpc4694 (
      {stage2_61[36], stage2_61[37], stage2_61[38], stage2_61[39], stage2_61[40], stage2_61[41]},
      {stage2_63[30], stage2_63[31], stage2_63[32], stage2_63[33], stage2_63[34], stage2_63[35]},
      {stage3_65[5],stage3_64[5],stage3_63[6],stage3_62[13],stage3_61[18]}
   );
   gpc606_5 gpc4695 (
      {stage2_61[42], stage2_61[43], stage2_61[44], stage2_61[45], stage2_61[46], stage2_61[47]},
      {stage2_63[36], stage2_63[37], stage2_63[38], stage2_63[39], stage2_63[40], stage2_63[41]},
      {stage3_65[6],stage3_64[6],stage3_63[7],stage3_62[14],stage3_61[19]}
   );
   gpc606_5 gpc4696 (
      {stage2_61[48], stage2_61[49], stage2_61[50], stage2_61[51], stage2_61[52], stage2_61[53]},
      {stage2_63[42], stage2_63[43], stage2_63[44], stage2_63[45], stage2_63[46], stage2_63[47]},
      {stage3_65[7],stage3_64[7],stage3_63[8],stage3_62[15],stage3_61[20]}
   );
   gpc1163_5 gpc4697 (
      {stage2_62[0], stage2_62[1], stage2_62[2]},
      {stage2_63[48], stage2_63[49], stage2_63[50], stage2_63[51], stage2_63[52], stage2_63[53]},
      {stage2_64[0]},
      {stage2_65[0]},
      {stage3_66[0],stage3_65[8],stage3_64[8],stage3_63[9],stage3_62[16]}
   );
   gpc1163_5 gpc4698 (
      {stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage2_63[54], stage2_63[55], stage2_63[56], stage2_63[57], stage2_63[58], stage2_63[59]},
      {stage2_64[1]},
      {stage2_65[1]},
      {stage3_66[1],stage3_65[9],stage3_64[9],stage3_63[10],stage3_62[17]}
   );
   gpc1163_5 gpc4699 (
      {stage2_62[6], stage2_62[7], stage2_62[8]},
      {stage2_63[60], stage2_63[61], stage2_63[62], stage2_63[63], stage2_63[64], stage2_63[65]},
      {stage2_64[2]},
      {stage2_65[2]},
      {stage3_66[2],stage3_65[10],stage3_64[10],stage3_63[11],stage3_62[18]}
   );
   gpc606_5 gpc4700 (
      {stage2_62[9], stage2_62[10], stage2_62[11], stage2_62[12], stage2_62[13], stage2_62[14]},
      {stage2_64[3], stage2_64[4], stage2_64[5], stage2_64[6], stage2_64[7], stage2_64[8]},
      {stage3_66[3],stage3_65[11],stage3_64[11],stage3_63[12],stage3_62[19]}
   );
   gpc606_5 gpc4701 (
      {stage2_62[15], stage2_62[16], stage2_62[17], stage2_62[18], stage2_62[19], stage2_62[20]},
      {stage2_64[9], stage2_64[10], stage2_64[11], stage2_64[12], stage2_64[13], stage2_64[14]},
      {stage3_66[4],stage3_65[12],stage3_64[12],stage3_63[13],stage3_62[20]}
   );
   gpc606_5 gpc4702 (
      {stage2_62[21], stage2_62[22], stage2_62[23], stage2_62[24], stage2_62[25], stage2_62[26]},
      {stage2_64[15], stage2_64[16], stage2_64[17], stage2_64[18], stage2_64[19], stage2_64[20]},
      {stage3_66[5],stage3_65[13],stage3_64[13],stage3_63[14],stage3_62[21]}
   );
   gpc606_5 gpc4703 (
      {stage2_62[27], stage2_62[28], stage2_62[29], stage2_62[30], stage2_62[31], stage2_62[32]},
      {stage2_64[21], stage2_64[22], stage2_64[23], stage2_64[24], stage2_64[25], stage2_64[26]},
      {stage3_66[6],stage3_65[14],stage3_64[14],stage3_63[15],stage3_62[22]}
   );
   gpc606_5 gpc4704 (
      {stage2_62[33], stage2_62[34], stage2_62[35], stage2_62[36], stage2_62[37], stage2_62[38]},
      {stage2_64[27], stage2_64[28], stage2_64[29], stage2_64[30], stage2_64[31], stage2_64[32]},
      {stage3_66[7],stage3_65[15],stage3_64[15],stage3_63[16],stage3_62[23]}
   );
   gpc606_5 gpc4705 (
      {stage2_62[39], stage2_62[40], stage2_62[41], stage2_62[42], stage2_62[43], stage2_62[44]},
      {stage2_64[33], stage2_64[34], stage2_64[35], stage2_64[36], stage2_64[37], stage2_64[38]},
      {stage3_66[8],stage3_65[16],stage3_64[16],stage3_63[17],stage3_62[24]}
   );
   gpc606_5 gpc4706 (
      {stage2_62[45], stage2_62[46], stage2_62[47], stage2_62[48], stage2_62[49], stage2_62[50]},
      {stage2_64[39], stage2_64[40], stage2_64[41], stage2_64[42], stage2_64[43], stage2_64[44]},
      {stage3_66[9],stage3_65[17],stage3_64[17],stage3_63[18],stage3_62[25]}
   );
   gpc606_5 gpc4707 (
      {stage2_65[3], stage2_65[4], stage2_65[5], stage2_65[6], stage2_65[7], stage2_65[8]},
      {stage2_67[0], stage2_67[1], stage2_67[2], stage2_67[3], stage2_67[4], stage2_67[5]},
      {stage3_69[0],stage3_68[0],stage3_67[0],stage3_66[10],stage3_65[18]}
   );
   gpc1_1 gpc4708 (
      {stage2_0[20]},
      {stage3_0[4]}
   );
   gpc1_1 gpc4709 (
      {stage2_0[21]},
      {stage3_0[5]}
   );
   gpc1_1 gpc4710 (
      {stage2_0[22]},
      {stage3_0[6]}
   );
   gpc1_1 gpc4711 (
      {stage2_0[23]},
      {stage3_0[7]}
   );
   gpc1_1 gpc4712 (
      {stage2_0[24]},
      {stage3_0[8]}
   );
   gpc1_1 gpc4713 (
      {stage2_0[25]},
      {stage3_0[9]}
   );
   gpc1_1 gpc4714 (
      {stage2_0[26]},
      {stage3_0[10]}
   );
   gpc1_1 gpc4715 (
      {stage2_0[27]},
      {stage3_0[11]}
   );
   gpc1_1 gpc4716 (
      {stage2_0[28]},
      {stage3_0[12]}
   );
   gpc1_1 gpc4717 (
      {stage2_0[29]},
      {stage3_0[13]}
   );
   gpc1_1 gpc4718 (
      {stage2_1[35]},
      {stage3_1[9]}
   );
   gpc1_1 gpc4719 (
      {stage2_1[36]},
      {stage3_1[10]}
   );
   gpc1_1 gpc4720 (
      {stage2_2[29]},
      {stage3_2[10]}
   );
   gpc1_1 gpc4721 (
      {stage2_2[30]},
      {stage3_2[11]}
   );
   gpc1_1 gpc4722 (
      {stage2_2[31]},
      {stage3_2[12]}
   );
   gpc1_1 gpc4723 (
      {stage2_2[32]},
      {stage3_2[13]}
   );
   gpc1_1 gpc4724 (
      {stage2_2[33]},
      {stage3_2[14]}
   );
   gpc1_1 gpc4725 (
      {stage2_2[34]},
      {stage3_2[15]}
   );
   gpc1_1 gpc4726 (
      {stage2_2[35]},
      {stage3_2[16]}
   );
   gpc1_1 gpc4727 (
      {stage2_2[36]},
      {stage3_2[17]}
   );
   gpc1_1 gpc4728 (
      {stage2_3[50]},
      {stage3_3[15]}
   );
   gpc1_1 gpc4729 (
      {stage2_3[51]},
      {stage3_3[16]}
   );
   gpc1_1 gpc4730 (
      {stage2_3[52]},
      {stage3_3[17]}
   );
   gpc1_1 gpc4731 (
      {stage2_3[53]},
      {stage3_3[18]}
   );
   gpc1_1 gpc4732 (
      {stage2_4[43]},
      {stage3_4[19]}
   );
   gpc1_1 gpc4733 (
      {stage2_4[44]},
      {stage3_4[20]}
   );
   gpc1_1 gpc4734 (
      {stage2_5[26]},
      {stage3_5[15]}
   );
   gpc1_1 gpc4735 (
      {stage2_5[27]},
      {stage3_5[16]}
   );
   gpc1_1 gpc4736 (
      {stage2_5[28]},
      {stage3_5[17]}
   );
   gpc1_1 gpc4737 (
      {stage2_5[29]},
      {stage3_5[18]}
   );
   gpc1_1 gpc4738 (
      {stage2_5[30]},
      {stage3_5[19]}
   );
   gpc1_1 gpc4739 (
      {stage2_5[31]},
      {stage3_5[20]}
   );
   gpc1_1 gpc4740 (
      {stage2_5[32]},
      {stage3_5[21]}
   );
   gpc1_1 gpc4741 (
      {stage2_5[33]},
      {stage3_5[22]}
   );
   gpc1_1 gpc4742 (
      {stage2_5[34]},
      {stage3_5[23]}
   );
   gpc1_1 gpc4743 (
      {stage2_5[35]},
      {stage3_5[24]}
   );
   gpc1_1 gpc4744 (
      {stage2_5[36]},
      {stage3_5[25]}
   );
   gpc1_1 gpc4745 (
      {stage2_5[37]},
      {stage3_5[26]}
   );
   gpc1_1 gpc4746 (
      {stage2_5[38]},
      {stage3_5[27]}
   );
   gpc1_1 gpc4747 (
      {stage2_5[39]},
      {stage3_5[28]}
   );
   gpc1_1 gpc4748 (
      {stage2_5[40]},
      {stage3_5[29]}
   );
   gpc1_1 gpc4749 (
      {stage2_5[41]},
      {stage3_5[30]}
   );
   gpc1_1 gpc4750 (
      {stage2_5[42]},
      {stage3_5[31]}
   );
   gpc1_1 gpc4751 (
      {stage2_5[43]},
      {stage3_5[32]}
   );
   gpc1_1 gpc4752 (
      {stage2_5[44]},
      {stage3_5[33]}
   );
   gpc1_1 gpc4753 (
      {stage2_5[45]},
      {stage3_5[34]}
   );
   gpc1_1 gpc4754 (
      {stage2_6[49]},
      {stage3_6[14]}
   );
   gpc1_1 gpc4755 (
      {stage2_6[50]},
      {stage3_6[15]}
   );
   gpc1_1 gpc4756 (
      {stage2_6[51]},
      {stage3_6[16]}
   );
   gpc1_1 gpc4757 (
      {stage2_7[35]},
      {stage3_7[20]}
   );
   gpc1_1 gpc4758 (
      {stage2_7[36]},
      {stage3_7[21]}
   );
   gpc1_1 gpc4759 (
      {stage2_7[37]},
      {stage3_7[22]}
   );
   gpc1_1 gpc4760 (
      {stage2_7[38]},
      {stage3_7[23]}
   );
   gpc1_1 gpc4761 (
      {stage2_7[39]},
      {stage3_7[24]}
   );
   gpc1_1 gpc4762 (
      {stage2_7[40]},
      {stage3_7[25]}
   );
   gpc1_1 gpc4763 (
      {stage2_7[41]},
      {stage3_7[26]}
   );
   gpc1_1 gpc4764 (
      {stage2_7[42]},
      {stage3_7[27]}
   );
   gpc1_1 gpc4765 (
      {stage2_10[60]},
      {stage3_10[23]}
   );
   gpc1_1 gpc4766 (
      {stage2_10[61]},
      {stage3_10[24]}
   );
   gpc1_1 gpc4767 (
      {stage2_10[62]},
      {stage3_10[25]}
   );
   gpc1_1 gpc4768 (
      {stage2_10[63]},
      {stage3_10[26]}
   );
   gpc1_1 gpc4769 (
      {stage2_10[64]},
      {stage3_10[27]}
   );
   gpc1_1 gpc4770 (
      {stage2_10[65]},
      {stage3_10[28]}
   );
   gpc1_1 gpc4771 (
      {stage2_10[66]},
      {stage3_10[29]}
   );
   gpc1_1 gpc4772 (
      {stage2_10[67]},
      {stage3_10[30]}
   );
   gpc1_1 gpc4773 (
      {stage2_10[68]},
      {stage3_10[31]}
   );
   gpc1_1 gpc4774 (
      {stage2_10[69]},
      {stage3_10[32]}
   );
   gpc1_1 gpc4775 (
      {stage2_11[43]},
      {stage3_11[25]}
   );
   gpc1_1 gpc4776 (
      {stage2_11[44]},
      {stage3_11[26]}
   );
   gpc1_1 gpc4777 (
      {stage2_11[45]},
      {stage3_11[27]}
   );
   gpc1_1 gpc4778 (
      {stage2_11[46]},
      {stage3_11[28]}
   );
   gpc1_1 gpc4779 (
      {stage2_11[47]},
      {stage3_11[29]}
   );
   gpc1_1 gpc4780 (
      {stage2_11[48]},
      {stage3_11[30]}
   );
   gpc1_1 gpc4781 (
      {stage2_12[47]},
      {stage3_12[18]}
   );
   gpc1_1 gpc4782 (
      {stage2_12[48]},
      {stage3_12[19]}
   );
   gpc1_1 gpc4783 (
      {stage2_12[49]},
      {stage3_12[20]}
   );
   gpc1_1 gpc4784 (
      {stage2_12[50]},
      {stage3_12[21]}
   );
   gpc1_1 gpc4785 (
      {stage2_12[51]},
      {stage3_12[22]}
   );
   gpc1_1 gpc4786 (
      {stage2_12[52]},
      {stage3_12[23]}
   );
   gpc1_1 gpc4787 (
      {stage2_12[53]},
      {stage3_12[24]}
   );
   gpc1_1 gpc4788 (
      {stage2_13[60]},
      {stage3_13[20]}
   );
   gpc1_1 gpc4789 (
      {stage2_13[61]},
      {stage3_13[21]}
   );
   gpc1_1 gpc4790 (
      {stage2_13[62]},
      {stage3_13[22]}
   );
   gpc1_1 gpc4791 (
      {stage2_13[63]},
      {stage3_13[23]}
   );
   gpc1_1 gpc4792 (
      {stage2_14[42]},
      {stage3_14[24]}
   );
   gpc1_1 gpc4793 (
      {stage2_14[43]},
      {stage3_14[25]}
   );
   gpc1_1 gpc4794 (
      {stage2_14[44]},
      {stage3_14[26]}
   );
   gpc1_1 gpc4795 (
      {stage2_15[55]},
      {stage3_15[22]}
   );
   gpc1_1 gpc4796 (
      {stage2_15[56]},
      {stage3_15[23]}
   );
   gpc1_1 gpc4797 (
      {stage2_15[57]},
      {stage3_15[24]}
   );
   gpc1_1 gpc4798 (
      {stage2_15[58]},
      {stage3_15[25]}
   );
   gpc1_1 gpc4799 (
      {stage2_15[59]},
      {stage3_15[26]}
   );
   gpc1_1 gpc4800 (
      {stage2_15[60]},
      {stage3_15[27]}
   );
   gpc1_1 gpc4801 (
      {stage2_15[61]},
      {stage3_15[28]}
   );
   gpc1_1 gpc4802 (
      {stage2_15[62]},
      {stage3_15[29]}
   );
   gpc1_1 gpc4803 (
      {stage2_15[63]},
      {stage3_15[30]}
   );
   gpc1_1 gpc4804 (
      {stage2_15[64]},
      {stage3_15[31]}
   );
   gpc1_1 gpc4805 (
      {stage2_15[65]},
      {stage3_15[32]}
   );
   gpc1_1 gpc4806 (
      {stage2_15[66]},
      {stage3_15[33]}
   );
   gpc1_1 gpc4807 (
      {stage2_15[67]},
      {stage3_15[34]}
   );
   gpc1_1 gpc4808 (
      {stage2_15[68]},
      {stage3_15[35]}
   );
   gpc1_1 gpc4809 (
      {stage2_15[69]},
      {stage3_15[36]}
   );
   gpc1_1 gpc4810 (
      {stage2_15[70]},
      {stage3_15[37]}
   );
   gpc1_1 gpc4811 (
      {stage2_15[71]},
      {stage3_15[38]}
   );
   gpc1_1 gpc4812 (
      {stage2_15[72]},
      {stage3_15[39]}
   );
   gpc1_1 gpc4813 (
      {stage2_15[73]},
      {stage3_15[40]}
   );
   gpc1_1 gpc4814 (
      {stage2_16[53]},
      {stage3_16[18]}
   );
   gpc1_1 gpc4815 (
      {stage2_16[54]},
      {stage3_16[19]}
   );
   gpc1_1 gpc4816 (
      {stage2_17[48]},
      {stage3_17[21]}
   );
   gpc1_1 gpc4817 (
      {stage2_17[49]},
      {stage3_17[22]}
   );
   gpc1_1 gpc4818 (
      {stage2_17[50]},
      {stage3_17[23]}
   );
   gpc1_1 gpc4819 (
      {stage2_17[51]},
      {stage3_17[24]}
   );
   gpc1_1 gpc4820 (
      {stage2_17[52]},
      {stage3_17[25]}
   );
   gpc1_1 gpc4821 (
      {stage2_17[53]},
      {stage3_17[26]}
   );
   gpc1_1 gpc4822 (
      {stage2_17[54]},
      {stage3_17[27]}
   );
   gpc1_1 gpc4823 (
      {stage2_17[55]},
      {stage3_17[28]}
   );
   gpc1_1 gpc4824 (
      {stage2_17[56]},
      {stage3_17[29]}
   );
   gpc1_1 gpc4825 (
      {stage2_19[30]},
      {stage3_19[21]}
   );
   gpc1_1 gpc4826 (
      {stage2_19[31]},
      {stage3_19[22]}
   );
   gpc1_1 gpc4827 (
      {stage2_19[32]},
      {stage3_19[23]}
   );
   gpc1_1 gpc4828 (
      {stage2_19[33]},
      {stage3_19[24]}
   );
   gpc1_1 gpc4829 (
      {stage2_19[34]},
      {stage3_19[25]}
   );
   gpc1_1 gpc4830 (
      {stage2_19[35]},
      {stage3_19[26]}
   );
   gpc1_1 gpc4831 (
      {stage2_19[36]},
      {stage3_19[27]}
   );
   gpc1_1 gpc4832 (
      {stage2_20[72]},
      {stage3_20[16]}
   );
   gpc1_1 gpc4833 (
      {stage2_20[73]},
      {stage3_20[17]}
   );
   gpc1_1 gpc4834 (
      {stage2_20[74]},
      {stage3_20[18]}
   );
   gpc1_1 gpc4835 (
      {stage2_20[75]},
      {stage3_20[19]}
   );
   gpc1_1 gpc4836 (
      {stage2_20[76]},
      {stage3_20[20]}
   );
   gpc1_1 gpc4837 (
      {stage2_20[77]},
      {stage3_20[21]}
   );
   gpc1_1 gpc4838 (
      {stage2_20[78]},
      {stage3_20[22]}
   );
   gpc1_1 gpc4839 (
      {stage2_20[79]},
      {stage3_20[23]}
   );
   gpc1_1 gpc4840 (
      {stage2_22[40]},
      {stage3_22[28]}
   );
   gpc1_1 gpc4841 (
      {stage2_24[72]},
      {stage3_24[21]}
   );
   gpc1_1 gpc4842 (
      {stage2_24[73]},
      {stage3_24[22]}
   );
   gpc1_1 gpc4843 (
      {stage2_24[74]},
      {stage3_24[23]}
   );
   gpc1_1 gpc4844 (
      {stage2_24[75]},
      {stage3_24[24]}
   );
   gpc1_1 gpc4845 (
      {stage2_24[76]},
      {stage3_24[25]}
   );
   gpc1_1 gpc4846 (
      {stage2_24[77]},
      {stage3_24[26]}
   );
   gpc1_1 gpc4847 (
      {stage2_24[78]},
      {stage3_24[27]}
   );
   gpc1_1 gpc4848 (
      {stage2_24[79]},
      {stage3_24[28]}
   );
   gpc1_1 gpc4849 (
      {stage2_24[80]},
      {stage3_24[29]}
   );
   gpc1_1 gpc4850 (
      {stage2_24[81]},
      {stage3_24[30]}
   );
   gpc1_1 gpc4851 (
      {stage2_25[46]},
      {stage3_25[29]}
   );
   gpc1_1 gpc4852 (
      {stage2_25[47]},
      {stage3_25[30]}
   );
   gpc1_1 gpc4853 (
      {stage2_25[48]},
      {stage3_25[31]}
   );
   gpc1_1 gpc4854 (
      {stage2_25[49]},
      {stage3_25[32]}
   );
   gpc1_1 gpc4855 (
      {stage2_25[50]},
      {stage3_25[33]}
   );
   gpc1_1 gpc4856 (
      {stage2_29[36]},
      {stage3_29[25]}
   );
   gpc1_1 gpc4857 (
      {stage2_29[37]},
      {stage3_29[26]}
   );
   gpc1_1 gpc4858 (
      {stage2_29[38]},
      {stage3_29[27]}
   );
   gpc1_1 gpc4859 (
      {stage2_29[39]},
      {stage3_29[28]}
   );
   gpc1_1 gpc4860 (
      {stage2_29[40]},
      {stage3_29[29]}
   );
   gpc1_1 gpc4861 (
      {stage2_29[41]},
      {stage3_29[30]}
   );
   gpc1_1 gpc4862 (
      {stage2_29[42]},
      {stage3_29[31]}
   );
   gpc1_1 gpc4863 (
      {stage2_29[43]},
      {stage3_29[32]}
   );
   gpc1_1 gpc4864 (
      {stage2_29[44]},
      {stage3_29[33]}
   );
   gpc1_1 gpc4865 (
      {stage2_29[45]},
      {stage3_29[34]}
   );
   gpc1_1 gpc4866 (
      {stage2_30[52]},
      {stage3_30[19]}
   );
   gpc1_1 gpc4867 (
      {stage2_30[53]},
      {stage3_30[20]}
   );
   gpc1_1 gpc4868 (
      {stage2_30[54]},
      {stage3_30[21]}
   );
   gpc1_1 gpc4869 (
      {stage2_30[55]},
      {stage3_30[22]}
   );
   gpc1_1 gpc4870 (
      {stage2_30[56]},
      {stage3_30[23]}
   );
   gpc1_1 gpc4871 (
      {stage2_30[57]},
      {stage3_30[24]}
   );
   gpc1_1 gpc4872 (
      {stage2_30[58]},
      {stage3_30[25]}
   );
   gpc1_1 gpc4873 (
      {stage2_31[43]},
      {stage3_31[21]}
   );
   gpc1_1 gpc4874 (
      {stage2_31[44]},
      {stage3_31[22]}
   );
   gpc1_1 gpc4875 (
      {stage2_31[45]},
      {stage3_31[23]}
   );
   gpc1_1 gpc4876 (
      {stage2_31[46]},
      {stage3_31[24]}
   );
   gpc1_1 gpc4877 (
      {stage2_31[47]},
      {stage3_31[25]}
   );
   gpc1_1 gpc4878 (
      {stage2_31[48]},
      {stage3_31[26]}
   );
   gpc1_1 gpc4879 (
      {stage2_31[49]},
      {stage3_31[27]}
   );
   gpc1_1 gpc4880 (
      {stage2_31[50]},
      {stage3_31[28]}
   );
   gpc1_1 gpc4881 (
      {stage2_31[51]},
      {stage3_31[29]}
   );
   gpc1_1 gpc4882 (
      {stage2_31[52]},
      {stage3_31[30]}
   );
   gpc1_1 gpc4883 (
      {stage2_31[53]},
      {stage3_31[31]}
   );
   gpc1_1 gpc4884 (
      {stage2_32[39]},
      {stage3_32[20]}
   );
   gpc1_1 gpc4885 (
      {stage2_32[40]},
      {stage3_32[21]}
   );
   gpc1_1 gpc4886 (
      {stage2_32[41]},
      {stage3_32[22]}
   );
   gpc1_1 gpc4887 (
      {stage2_32[42]},
      {stage3_32[23]}
   );
   gpc1_1 gpc4888 (
      {stage2_32[43]},
      {stage3_32[24]}
   );
   gpc1_1 gpc4889 (
      {stage2_32[44]},
      {stage3_32[25]}
   );
   gpc1_1 gpc4890 (
      {stage2_32[45]},
      {stage3_32[26]}
   );
   gpc1_1 gpc4891 (
      {stage2_32[46]},
      {stage3_32[27]}
   );
   gpc1_1 gpc4892 (
      {stage2_33[38]},
      {stage3_33[13]}
   );
   gpc1_1 gpc4893 (
      {stage2_33[39]},
      {stage3_33[14]}
   );
   gpc1_1 gpc4894 (
      {stage2_33[40]},
      {stage3_33[15]}
   );
   gpc1_1 gpc4895 (
      {stage2_33[41]},
      {stage3_33[16]}
   );
   gpc1_1 gpc4896 (
      {stage2_33[42]},
      {stage3_33[17]}
   );
   gpc1_1 gpc4897 (
      {stage2_33[43]},
      {stage3_33[18]}
   );
   gpc1_1 gpc4898 (
      {stage2_33[44]},
      {stage3_33[19]}
   );
   gpc1_1 gpc4899 (
      {stage2_33[45]},
      {stage3_33[20]}
   );
   gpc1_1 gpc4900 (
      {stage2_33[46]},
      {stage3_33[21]}
   );
   gpc1_1 gpc4901 (
      {stage2_33[47]},
      {stage3_33[22]}
   );
   gpc1_1 gpc4902 (
      {stage2_33[48]},
      {stage3_33[23]}
   );
   gpc1_1 gpc4903 (
      {stage2_33[49]},
      {stage3_33[24]}
   );
   gpc1_1 gpc4904 (
      {stage2_33[50]},
      {stage3_33[25]}
   );
   gpc1_1 gpc4905 (
      {stage2_33[51]},
      {stage3_33[26]}
   );
   gpc1_1 gpc4906 (
      {stage2_34[24]},
      {stage3_34[14]}
   );
   gpc1_1 gpc4907 (
      {stage2_34[25]},
      {stage3_34[15]}
   );
   gpc1_1 gpc4908 (
      {stage2_34[26]},
      {stage3_34[16]}
   );
   gpc1_1 gpc4909 (
      {stage2_34[27]},
      {stage3_34[17]}
   );
   gpc1_1 gpc4910 (
      {stage2_34[28]},
      {stage3_34[18]}
   );
   gpc1_1 gpc4911 (
      {stage2_34[29]},
      {stage3_34[19]}
   );
   gpc1_1 gpc4912 (
      {stage2_34[30]},
      {stage3_34[20]}
   );
   gpc1_1 gpc4913 (
      {stage2_34[31]},
      {stage3_34[21]}
   );
   gpc1_1 gpc4914 (
      {stage2_34[32]},
      {stage3_34[22]}
   );
   gpc1_1 gpc4915 (
      {stage2_34[33]},
      {stage3_34[23]}
   );
   gpc1_1 gpc4916 (
      {stage2_34[34]},
      {stage3_34[24]}
   );
   gpc1_1 gpc4917 (
      {stage2_34[35]},
      {stage3_34[25]}
   );
   gpc1_1 gpc4918 (
      {stage2_34[36]},
      {stage3_34[26]}
   );
   gpc1_1 gpc4919 (
      {stage2_35[47]},
      {stage3_35[21]}
   );
   gpc1_1 gpc4920 (
      {stage2_35[48]},
      {stage3_35[22]}
   );
   gpc1_1 gpc4921 (
      {stage2_35[49]},
      {stage3_35[23]}
   );
   gpc1_1 gpc4922 (
      {stage2_35[50]},
      {stage3_35[24]}
   );
   gpc1_1 gpc4923 (
      {stage2_35[51]},
      {stage3_35[25]}
   );
   gpc1_1 gpc4924 (
      {stage2_35[52]},
      {stage3_35[26]}
   );
   gpc1_1 gpc4925 (
      {stage2_35[53]},
      {stage3_35[27]}
   );
   gpc1_1 gpc4926 (
      {stage2_35[54]},
      {stage3_35[28]}
   );
   gpc1_1 gpc4927 (
      {stage2_35[55]},
      {stage3_35[29]}
   );
   gpc1_1 gpc4928 (
      {stage2_35[56]},
      {stage3_35[30]}
   );
   gpc1_1 gpc4929 (
      {stage2_35[57]},
      {stage3_35[31]}
   );
   gpc1_1 gpc4930 (
      {stage2_35[58]},
      {stage3_35[32]}
   );
   gpc1_1 gpc4931 (
      {stage2_37[54]},
      {stage3_37[18]}
   );
   gpc1_1 gpc4932 (
      {stage2_38[42]},
      {stage3_38[18]}
   );
   gpc1_1 gpc4933 (
      {stage2_38[43]},
      {stage3_38[19]}
   );
   gpc1_1 gpc4934 (
      {stage2_38[44]},
      {stage3_38[20]}
   );
   gpc1_1 gpc4935 (
      {stage2_38[45]},
      {stage3_38[21]}
   );
   gpc1_1 gpc4936 (
      {stage2_38[46]},
      {stage3_38[22]}
   );
   gpc1_1 gpc4937 (
      {stage2_40[39]},
      {stage3_40[24]}
   );
   gpc1_1 gpc4938 (
      {stage2_40[40]},
      {stage3_40[25]}
   );
   gpc1_1 gpc4939 (
      {stage2_40[41]},
      {stage3_40[26]}
   );
   gpc1_1 gpc4940 (
      {stage2_40[42]},
      {stage3_40[27]}
   );
   gpc1_1 gpc4941 (
      {stage2_40[43]},
      {stage3_40[28]}
   );
   gpc1_1 gpc4942 (
      {stage2_40[44]},
      {stage3_40[29]}
   );
   gpc1_1 gpc4943 (
      {stage2_42[58]},
      {stage3_42[25]}
   );
   gpc1_1 gpc4944 (
      {stage2_42[59]},
      {stage3_42[26]}
   );
   gpc1_1 gpc4945 (
      {stage2_42[60]},
      {stage3_42[27]}
   );
   gpc1_1 gpc4946 (
      {stage2_42[61]},
      {stage3_42[28]}
   );
   gpc1_1 gpc4947 (
      {stage2_42[62]},
      {stage3_42[29]}
   );
   gpc1_1 gpc4948 (
      {stage2_43[54]},
      {stage3_43[31]}
   );
   gpc1_1 gpc4949 (
      {stage2_43[55]},
      {stage3_43[32]}
   );
   gpc1_1 gpc4950 (
      {stage2_43[56]},
      {stage3_43[33]}
   );
   gpc1_1 gpc4951 (
      {stage2_43[57]},
      {stage3_43[34]}
   );
   gpc1_1 gpc4952 (
      {stage2_43[58]},
      {stage3_43[35]}
   );
   gpc1_1 gpc4953 (
      {stage2_43[59]},
      {stage3_43[36]}
   );
   gpc1_1 gpc4954 (
      {stage2_43[60]},
      {stage3_43[37]}
   );
   gpc1_1 gpc4955 (
      {stage2_43[61]},
      {stage3_43[38]}
   );
   gpc1_1 gpc4956 (
      {stage2_45[66]},
      {stage3_45[26]}
   );
   gpc1_1 gpc4957 (
      {stage2_45[67]},
      {stage3_45[27]}
   );
   gpc1_1 gpc4958 (
      {stage2_45[68]},
      {stage3_45[28]}
   );
   gpc1_1 gpc4959 (
      {stage2_45[69]},
      {stage3_45[29]}
   );
   gpc1_1 gpc4960 (
      {stage2_45[70]},
      {stage3_45[30]}
   );
   gpc1_1 gpc4961 (
      {stage2_45[71]},
      {stage3_45[31]}
   );
   gpc1_1 gpc4962 (
      {stage2_45[72]},
      {stage3_45[32]}
   );
   gpc1_1 gpc4963 (
      {stage2_45[73]},
      {stage3_45[33]}
   );
   gpc1_1 gpc4964 (
      {stage2_45[74]},
      {stage3_45[34]}
   );
   gpc1_1 gpc4965 (
      {stage2_45[75]},
      {stage3_45[35]}
   );
   gpc1_1 gpc4966 (
      {stage2_45[76]},
      {stage3_45[36]}
   );
   gpc1_1 gpc4967 (
      {stage2_45[77]},
      {stage3_45[37]}
   );
   gpc1_1 gpc4968 (
      {stage2_45[78]},
      {stage3_45[38]}
   );
   gpc1_1 gpc4969 (
      {stage2_46[42]},
      {stage3_46[19]}
   );
   gpc1_1 gpc4970 (
      {stage2_46[43]},
      {stage3_46[20]}
   );
   gpc1_1 gpc4971 (
      {stage2_46[44]},
      {stage3_46[21]}
   );
   gpc1_1 gpc4972 (
      {stage2_46[45]},
      {stage3_46[22]}
   );
   gpc1_1 gpc4973 (
      {stage2_46[46]},
      {stage3_46[23]}
   );
   gpc1_1 gpc4974 (
      {stage2_46[47]},
      {stage3_46[24]}
   );
   gpc1_1 gpc4975 (
      {stage2_46[48]},
      {stage3_46[25]}
   );
   gpc1_1 gpc4976 (
      {stage2_46[49]},
      {stage3_46[26]}
   );
   gpc1_1 gpc4977 (
      {stage2_46[50]},
      {stage3_46[27]}
   );
   gpc1_1 gpc4978 (
      {stage2_46[51]},
      {stage3_46[28]}
   );
   gpc1_1 gpc4979 (
      {stage2_46[52]},
      {stage3_46[29]}
   );
   gpc1_1 gpc4980 (
      {stage2_46[53]},
      {stage3_46[30]}
   );
   gpc1_1 gpc4981 (
      {stage2_46[54]},
      {stage3_46[31]}
   );
   gpc1_1 gpc4982 (
      {stage2_46[55]},
      {stage3_46[32]}
   );
   gpc1_1 gpc4983 (
      {stage2_46[56]},
      {stage3_46[33]}
   );
   gpc1_1 gpc4984 (
      {stage2_46[57]},
      {stage3_46[34]}
   );
   gpc1_1 gpc4985 (
      {stage2_46[58]},
      {stage3_46[35]}
   );
   gpc1_1 gpc4986 (
      {stage2_46[59]},
      {stage3_46[36]}
   );
   gpc1_1 gpc4987 (
      {stage2_46[60]},
      {stage3_46[37]}
   );
   gpc1_1 gpc4988 (
      {stage2_46[61]},
      {stage3_46[38]}
   );
   gpc1_1 gpc4989 (
      {stage2_46[62]},
      {stage3_46[39]}
   );
   gpc1_1 gpc4990 (
      {stage2_47[61]},
      {stage3_47[23]}
   );
   gpc1_1 gpc4991 (
      {stage2_47[62]},
      {stage3_47[24]}
   );
   gpc1_1 gpc4992 (
      {stage2_47[63]},
      {stage3_47[25]}
   );
   gpc1_1 gpc4993 (
      {stage2_47[64]},
      {stage3_47[26]}
   );
   gpc1_1 gpc4994 (
      {stage2_47[65]},
      {stage3_47[27]}
   );
   gpc1_1 gpc4995 (
      {stage2_47[66]},
      {stage3_47[28]}
   );
   gpc1_1 gpc4996 (
      {stage2_47[67]},
      {stage3_47[29]}
   );
   gpc1_1 gpc4997 (
      {stage2_47[68]},
      {stage3_47[30]}
   );
   gpc1_1 gpc4998 (
      {stage2_47[69]},
      {stage3_47[31]}
   );
   gpc1_1 gpc4999 (
      {stage2_47[70]},
      {stage3_47[32]}
   );
   gpc1_1 gpc5000 (
      {stage2_49[70]},
      {stage3_49[23]}
   );
   gpc1_1 gpc5001 (
      {stage2_49[71]},
      {stage3_49[24]}
   );
   gpc1_1 gpc5002 (
      {stage2_49[72]},
      {stage3_49[25]}
   );
   gpc1_1 gpc5003 (
      {stage2_49[73]},
      {stage3_49[26]}
   );
   gpc1_1 gpc5004 (
      {stage2_49[74]},
      {stage3_49[27]}
   );
   gpc1_1 gpc5005 (
      {stage2_49[75]},
      {stage3_49[28]}
   );
   gpc1_1 gpc5006 (
      {stage2_49[76]},
      {stage3_49[29]}
   );
   gpc1_1 gpc5007 (
      {stage2_49[77]},
      {stage3_49[30]}
   );
   gpc1_1 gpc5008 (
      {stage2_49[78]},
      {stage3_49[31]}
   );
   gpc1_1 gpc5009 (
      {stage2_49[79]},
      {stage3_49[32]}
   );
   gpc1_1 gpc5010 (
      {stage2_49[80]},
      {stage3_49[33]}
   );
   gpc1_1 gpc5011 (
      {stage2_49[81]},
      {stage3_49[34]}
   );
   gpc1_1 gpc5012 (
      {stage2_49[82]},
      {stage3_49[35]}
   );
   gpc1_1 gpc5013 (
      {stage2_49[83]},
      {stage3_49[36]}
   );
   gpc1_1 gpc5014 (
      {stage2_49[84]},
      {stage3_49[37]}
   );
   gpc1_1 gpc5015 (
      {stage2_49[85]},
      {stage3_49[38]}
   );
   gpc1_1 gpc5016 (
      {stage2_49[86]},
      {stage3_49[39]}
   );
   gpc1_1 gpc5017 (
      {stage2_49[87]},
      {stage3_49[40]}
   );
   gpc1_1 gpc5018 (
      {stage2_49[88]},
      {stage3_49[41]}
   );
   gpc1_1 gpc5019 (
      {stage2_49[89]},
      {stage3_49[42]}
   );
   gpc1_1 gpc5020 (
      {stage2_49[90]},
      {stage3_49[43]}
   );
   gpc1_1 gpc5021 (
      {stage2_49[91]},
      {stage3_49[44]}
   );
   gpc1_1 gpc5022 (
      {stage2_49[92]},
      {stage3_49[45]}
   );
   gpc1_1 gpc5023 (
      {stage2_49[93]},
      {stage3_49[46]}
   );
   gpc1_1 gpc5024 (
      {stage2_49[94]},
      {stage3_49[47]}
   );
   gpc1_1 gpc5025 (
      {stage2_49[95]},
      {stage3_49[48]}
   );
   gpc1_1 gpc5026 (
      {stage2_49[96]},
      {stage3_49[49]}
   );
   gpc1_1 gpc5027 (
      {stage2_49[97]},
      {stage3_49[50]}
   );
   gpc1_1 gpc5028 (
      {stage2_49[98]},
      {stage3_49[51]}
   );
   gpc1_1 gpc5029 (
      {stage2_49[99]},
      {stage3_49[52]}
   );
   gpc1_1 gpc5030 (
      {stage2_49[100]},
      {stage3_49[53]}
   );
   gpc1_1 gpc5031 (
      {stage2_49[101]},
      {stage3_49[54]}
   );
   gpc1_1 gpc5032 (
      {stage2_49[102]},
      {stage3_49[55]}
   );
   gpc1_1 gpc5033 (
      {stage2_49[103]},
      {stage3_49[56]}
   );
   gpc1_1 gpc5034 (
      {stage2_49[104]},
      {stage3_49[57]}
   );
   gpc1_1 gpc5035 (
      {stage2_49[105]},
      {stage3_49[58]}
   );
   gpc1_1 gpc5036 (
      {stage2_49[106]},
      {stage3_49[59]}
   );
   gpc1_1 gpc5037 (
      {stage2_49[107]},
      {stage3_49[60]}
   );
   gpc1_1 gpc5038 (
      {stage2_49[108]},
      {stage3_49[61]}
   );
   gpc1_1 gpc5039 (
      {stage2_49[109]},
      {stage3_49[62]}
   );
   gpc1_1 gpc5040 (
      {stage2_49[110]},
      {stage3_49[63]}
   );
   gpc1_1 gpc5041 (
      {stage2_49[111]},
      {stage3_49[64]}
   );
   gpc1_1 gpc5042 (
      {stage2_49[112]},
      {stage3_49[65]}
   );
   gpc1_1 gpc5043 (
      {stage2_49[113]},
      {stage3_49[66]}
   );
   gpc1_1 gpc5044 (
      {stage2_49[114]},
      {stage3_49[67]}
   );
   gpc1_1 gpc5045 (
      {stage2_50[57]},
      {stage3_50[19]}
   );
   gpc1_1 gpc5046 (
      {stage2_50[58]},
      {stage3_50[20]}
   );
   gpc1_1 gpc5047 (
      {stage2_50[59]},
      {stage3_50[21]}
   );
   gpc1_1 gpc5048 (
      {stage2_50[60]},
      {stage3_50[22]}
   );
   gpc1_1 gpc5049 (
      {stage2_50[61]},
      {stage3_50[23]}
   );
   gpc1_1 gpc5050 (
      {stage2_50[62]},
      {stage3_50[24]}
   );
   gpc1_1 gpc5051 (
      {stage2_50[63]},
      {stage3_50[25]}
   );
   gpc1_1 gpc5052 (
      {stage2_50[64]},
      {stage3_50[26]}
   );
   gpc1_1 gpc5053 (
      {stage2_50[65]},
      {stage3_50[27]}
   );
   gpc1_1 gpc5054 (
      {stage2_50[66]},
      {stage3_50[28]}
   );
   gpc1_1 gpc5055 (
      {stage2_50[67]},
      {stage3_50[29]}
   );
   gpc1_1 gpc5056 (
      {stage2_51[61]},
      {stage3_51[30]}
   );
   gpc1_1 gpc5057 (
      {stage2_51[62]},
      {stage3_51[31]}
   );
   gpc1_1 gpc5058 (
      {stage2_51[63]},
      {stage3_51[32]}
   );
   gpc1_1 gpc5059 (
      {stage2_51[64]},
      {stage3_51[33]}
   );
   gpc1_1 gpc5060 (
      {stage2_51[65]},
      {stage3_51[34]}
   );
   gpc1_1 gpc5061 (
      {stage2_51[66]},
      {stage3_51[35]}
   );
   gpc1_1 gpc5062 (
      {stage2_51[67]},
      {stage3_51[36]}
   );
   gpc1_1 gpc5063 (
      {stage2_51[68]},
      {stage3_51[37]}
   );
   gpc1_1 gpc5064 (
      {stage2_51[69]},
      {stage3_51[38]}
   );
   gpc1_1 gpc5065 (
      {stage2_51[70]},
      {stage3_51[39]}
   );
   gpc1_1 gpc5066 (
      {stage2_51[71]},
      {stage3_51[40]}
   );
   gpc1_1 gpc5067 (
      {stage2_51[72]},
      {stage3_51[41]}
   );
   gpc1_1 gpc5068 (
      {stage2_51[73]},
      {stage3_51[42]}
   );
   gpc1_1 gpc5069 (
      {stage2_51[74]},
      {stage3_51[43]}
   );
   gpc1_1 gpc5070 (
      {stage2_51[75]},
      {stage3_51[44]}
   );
   gpc1_1 gpc5071 (
      {stage2_51[76]},
      {stage3_51[45]}
   );
   gpc1_1 gpc5072 (
      {stage2_51[77]},
      {stage3_51[46]}
   );
   gpc1_1 gpc5073 (
      {stage2_51[78]},
      {stage3_51[47]}
   );
   gpc1_1 gpc5074 (
      {stage2_52[39]},
      {stage3_52[28]}
   );
   gpc1_1 gpc5075 (
      {stage2_52[40]},
      {stage3_52[29]}
   );
   gpc1_1 gpc5076 (
      {stage2_52[41]},
      {stage3_52[30]}
   );
   gpc1_1 gpc5077 (
      {stage2_52[42]},
      {stage3_52[31]}
   );
   gpc1_1 gpc5078 (
      {stage2_52[43]},
      {stage3_52[32]}
   );
   gpc1_1 gpc5079 (
      {stage2_52[44]},
      {stage3_52[33]}
   );
   gpc1_1 gpc5080 (
      {stage2_52[45]},
      {stage3_52[34]}
   );
   gpc1_1 gpc5081 (
      {stage2_52[46]},
      {stage3_52[35]}
   );
   gpc1_1 gpc5082 (
      {stage2_52[47]},
      {stage3_52[36]}
   );
   gpc1_1 gpc5083 (
      {stage2_52[48]},
      {stage3_52[37]}
   );
   gpc1_1 gpc5084 (
      {stage2_52[49]},
      {stage3_52[38]}
   );
   gpc1_1 gpc5085 (
      {stage2_52[50]},
      {stage3_52[39]}
   );
   gpc1_1 gpc5086 (
      {stage2_53[66]},
      {stage3_53[16]}
   );
   gpc1_1 gpc5087 (
      {stage2_53[67]},
      {stage3_53[17]}
   );
   gpc1_1 gpc5088 (
      {stage2_53[68]},
      {stage3_53[18]}
   );
   gpc1_1 gpc5089 (
      {stage2_53[69]},
      {stage3_53[19]}
   );
   gpc1_1 gpc5090 (
      {stage2_53[70]},
      {stage3_53[20]}
   );
   gpc1_1 gpc5091 (
      {stage2_53[71]},
      {stage3_53[21]}
   );
   gpc1_1 gpc5092 (
      {stage2_53[72]},
      {stage3_53[22]}
   );
   gpc1_1 gpc5093 (
      {stage2_53[73]},
      {stage3_53[23]}
   );
   gpc1_1 gpc5094 (
      {stage2_53[74]},
      {stage3_53[24]}
   );
   gpc1_1 gpc5095 (
      {stage2_53[75]},
      {stage3_53[25]}
   );
   gpc1_1 gpc5096 (
      {stage2_53[76]},
      {stage3_53[26]}
   );
   gpc1_1 gpc5097 (
      {stage2_53[77]},
      {stage3_53[27]}
   );
   gpc1_1 gpc5098 (
      {stage2_54[72]},
      {stage3_54[25]}
   );
   gpc1_1 gpc5099 (
      {stage2_54[73]},
      {stage3_54[26]}
   );
   gpc1_1 gpc5100 (
      {stage2_54[74]},
      {stage3_54[27]}
   );
   gpc1_1 gpc5101 (
      {stage2_56[67]},
      {stage3_56[20]}
   );
   gpc1_1 gpc5102 (
      {stage2_56[68]},
      {stage3_56[21]}
   );
   gpc1_1 gpc5103 (
      {stage2_56[69]},
      {stage3_56[22]}
   );
   gpc1_1 gpc5104 (
      {stage2_56[70]},
      {stage3_56[23]}
   );
   gpc1_1 gpc5105 (
      {stage2_56[71]},
      {stage3_56[24]}
   );
   gpc1_1 gpc5106 (
      {stage2_56[72]},
      {stage3_56[25]}
   );
   gpc1_1 gpc5107 (
      {stage2_57[72]},
      {stage3_57[22]}
   );
   gpc1_1 gpc5108 (
      {stage2_57[73]},
      {stage3_57[23]}
   );
   gpc1_1 gpc5109 (
      {stage2_57[74]},
      {stage3_57[24]}
   );
   gpc1_1 gpc5110 (
      {stage2_57[75]},
      {stage3_57[25]}
   );
   gpc1_1 gpc5111 (
      {stage2_57[76]},
      {stage3_57[26]}
   );
   gpc1_1 gpc5112 (
      {stage2_57[77]},
      {stage3_57[27]}
   );
   gpc1_1 gpc5113 (
      {stage2_57[78]},
      {stage3_57[28]}
   );
   gpc1_1 gpc5114 (
      {stage2_57[79]},
      {stage3_57[29]}
   );
   gpc1_1 gpc5115 (
      {stage2_57[80]},
      {stage3_57[30]}
   );
   gpc1_1 gpc5116 (
      {stage2_57[81]},
      {stage3_57[31]}
   );
   gpc1_1 gpc5117 (
      {stage2_57[82]},
      {stage3_57[32]}
   );
   gpc1_1 gpc5118 (
      {stage2_59[36]},
      {stage3_59[21]}
   );
   gpc1_1 gpc5119 (
      {stage2_59[37]},
      {stage3_59[22]}
   );
   gpc1_1 gpc5120 (
      {stage2_59[38]},
      {stage3_59[23]}
   );
   gpc1_1 gpc5121 (
      {stage2_59[39]},
      {stage3_59[24]}
   );
   gpc1_1 gpc5122 (
      {stage2_59[40]},
      {stage3_59[25]}
   );
   gpc1_1 gpc5123 (
      {stage2_59[41]},
      {stage3_59[26]}
   );
   gpc1_1 gpc5124 (
      {stage2_59[42]},
      {stage3_59[27]}
   );
   gpc1_1 gpc5125 (
      {stage2_59[43]},
      {stage3_59[28]}
   );
   gpc1_1 gpc5126 (
      {stage2_59[44]},
      {stage3_59[29]}
   );
   gpc1_1 gpc5127 (
      {stage2_59[45]},
      {stage3_59[30]}
   );
   gpc1_1 gpc5128 (
      {stage2_59[46]},
      {stage3_59[31]}
   );
   gpc1_1 gpc5129 (
      {stage2_59[47]},
      {stage3_59[32]}
   );
   gpc1_1 gpc5130 (
      {stage2_60[42]},
      {stage3_60[14]}
   );
   gpc1_1 gpc5131 (
      {stage2_60[43]},
      {stage3_60[15]}
   );
   gpc1_1 gpc5132 (
      {stage2_60[44]},
      {stage3_60[16]}
   );
   gpc1_1 gpc5133 (
      {stage2_60[45]},
      {stage3_60[17]}
   );
   gpc1_1 gpc5134 (
      {stage2_60[46]},
      {stage3_60[18]}
   );
   gpc1_1 gpc5135 (
      {stage2_60[47]},
      {stage3_60[19]}
   );
   gpc1_1 gpc5136 (
      {stage2_60[48]},
      {stage3_60[20]}
   );
   gpc1_1 gpc5137 (
      {stage2_60[49]},
      {stage3_60[21]}
   );
   gpc1_1 gpc5138 (
      {stage2_60[50]},
      {stage3_60[22]}
   );
   gpc1_1 gpc5139 (
      {stage2_60[51]},
      {stage3_60[23]}
   );
   gpc1_1 gpc5140 (
      {stage2_60[52]},
      {stage3_60[24]}
   );
   gpc1_1 gpc5141 (
      {stage2_60[53]},
      {stage3_60[25]}
   );
   gpc1_1 gpc5142 (
      {stage2_60[54]},
      {stage3_60[26]}
   );
   gpc1_1 gpc5143 (
      {stage2_60[55]},
      {stage3_60[27]}
   );
   gpc1_1 gpc5144 (
      {stage2_60[56]},
      {stage3_60[28]}
   );
   gpc1_1 gpc5145 (
      {stage2_60[57]},
      {stage3_60[29]}
   );
   gpc1_1 gpc5146 (
      {stage2_60[58]},
      {stage3_60[30]}
   );
   gpc1_1 gpc5147 (
      {stage2_60[59]},
      {stage3_60[31]}
   );
   gpc1_1 gpc5148 (
      {stage2_60[60]},
      {stage3_60[32]}
   );
   gpc1_1 gpc5149 (
      {stage2_60[61]},
      {stage3_60[33]}
   );
   gpc1_1 gpc5150 (
      {stage2_60[62]},
      {stage3_60[34]}
   );
   gpc1_1 gpc5151 (
      {stage2_61[54]},
      {stage3_61[21]}
   );
   gpc1_1 gpc5152 (
      {stage2_61[55]},
      {stage3_61[22]}
   );
   gpc1_1 gpc5153 (
      {stage2_61[56]},
      {stage3_61[23]}
   );
   gpc1_1 gpc5154 (
      {stage2_62[51]},
      {stage3_62[26]}
   );
   gpc1_1 gpc5155 (
      {stage2_62[52]},
      {stage3_62[27]}
   );
   gpc1_1 gpc5156 (
      {stage2_63[66]},
      {stage3_63[19]}
   );
   gpc1_1 gpc5157 (
      {stage2_63[67]},
      {stage3_63[20]}
   );
   gpc1_1 gpc5158 (
      {stage2_63[68]},
      {stage3_63[21]}
   );
   gpc1_1 gpc5159 (
      {stage2_63[69]},
      {stage3_63[22]}
   );
   gpc1_1 gpc5160 (
      {stage2_63[70]},
      {stage3_63[23]}
   );
   gpc1_1 gpc5161 (
      {stage2_63[71]},
      {stage3_63[24]}
   );
   gpc1_1 gpc5162 (
      {stage2_63[72]},
      {stage3_63[25]}
   );
   gpc1_1 gpc5163 (
      {stage2_63[73]},
      {stage3_63[26]}
   );
   gpc1_1 gpc5164 (
      {stage2_63[74]},
      {stage3_63[27]}
   );
   gpc1_1 gpc5165 (
      {stage2_65[9]},
      {stage3_65[19]}
   );
   gpc1_1 gpc5166 (
      {stage2_65[10]},
      {stage3_65[20]}
   );
   gpc1_1 gpc5167 (
      {stage2_65[11]},
      {stage3_65[21]}
   );
   gpc1_1 gpc5168 (
      {stage2_65[12]},
      {stage3_65[22]}
   );
   gpc1_1 gpc5169 (
      {stage2_65[13]},
      {stage3_65[23]}
   );
   gpc1_1 gpc5170 (
      {stage2_65[14]},
      {stage3_65[24]}
   );
   gpc1_1 gpc5171 (
      {stage2_65[15]},
      {stage3_65[25]}
   );
   gpc1_1 gpc5172 (
      {stage2_65[16]},
      {stage3_65[26]}
   );
   gpc1_1 gpc5173 (
      {stage2_65[17]},
      {stage3_65[27]}
   );
   gpc1_1 gpc5174 (
      {stage2_66[0]},
      {stage3_66[11]}
   );
   gpc1_1 gpc5175 (
      {stage2_66[1]},
      {stage3_66[12]}
   );
   gpc1_1 gpc5176 (
      {stage2_66[2]},
      {stage3_66[13]}
   );
   gpc1_1 gpc5177 (
      {stage2_66[3]},
      {stage3_66[14]}
   );
   gpc1_1 gpc5178 (
      {stage2_66[4]},
      {stage3_66[15]}
   );
   gpc1_1 gpc5179 (
      {stage2_66[5]},
      {stage3_66[16]}
   );
   gpc1_1 gpc5180 (
      {stage2_66[6]},
      {stage3_66[17]}
   );
   gpc1_1 gpc5181 (
      {stage2_66[7]},
      {stage3_66[18]}
   );
   gpc1_1 gpc5182 (
      {stage2_66[8]},
      {stage3_66[19]}
   );
   gpc1_1 gpc5183 (
      {stage2_66[9]},
      {stage3_66[20]}
   );
   gpc1_1 gpc5184 (
      {stage2_66[10]},
      {stage3_66[21]}
   );
   gpc1_1 gpc5185 (
      {stage2_66[11]},
      {stage3_66[22]}
   );
   gpc1_1 gpc5186 (
      {stage2_66[12]},
      {stage3_66[23]}
   );
   gpc1_1 gpc5187 (
      {stage2_66[13]},
      {stage3_66[24]}
   );
   gpc1_1 gpc5188 (
      {stage2_66[14]},
      {stage3_66[25]}
   );
   gpc1_1 gpc5189 (
      {stage2_66[15]},
      {stage3_66[26]}
   );
   gpc1_1 gpc5190 (
      {stage2_66[16]},
      {stage3_66[27]}
   );
   gpc1_1 gpc5191 (
      {stage2_67[6]},
      {stage3_67[1]}
   );
   gpc2135_5 gpc5192 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4]},
      {stage3_2[0], stage3_2[1], stage3_2[2]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc1163_5 gpc5193 (
      {stage3_1[5], stage3_1[6], stage3_1[7]},
      {stage3_2[3], stage3_2[4], stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8]},
      {stage3_3[1]},
      {stage3_4[2]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc5194 (
      {stage3_2[9], stage3_2[10], stage3_2[11], stage3_2[12], stage3_2[13]},
      {stage3_3[2]},
      {stage3_4[3], stage3_4[4], stage3_4[5], stage3_4[6], stage3_4[7], stage3_4[8]},
      {stage4_6[0],stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc606_5 gpc5195 (
      {stage3_4[9], stage3_4[10], stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[3],stage4_4[3]}
   );
   gpc1343_5 gpc5196 (
      {stage3_5[0], stage3_5[1], stage3_5[2]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[0], stage3_7[1], stage3_7[2]},
      {stage3_8[0]},
      {stage4_9[0],stage4_8[1],stage4_7[1],stage4_6[2],stage4_5[4]}
   );
   gpc1343_5 gpc5197 (
      {stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_6[10], stage3_6[11], stage3_6[12], stage3_6[13]},
      {stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[1]},
      {stage4_9[1],stage4_8[2],stage4_7[2],stage4_6[3],stage4_5[5]}
   );
   gpc606_5 gpc5198 (
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[2],stage4_8[3],stage4_7[3],stage4_6[4],stage4_5[6]}
   );
   gpc606_5 gpc5199 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[3],stage4_8[4],stage4_7[4],stage4_6[5],stage4_5[7]}
   );
   gpc606_5 gpc5200 (
      {stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21], stage3_5[22], stage3_5[23]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[4],stage4_8[5],stage4_7[5],stage4_6[6],stage4_5[8]}
   );
   gpc606_5 gpc5201 (
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[0],stage4_9[5]}
   );
   gpc615_5 gpc5202 (
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10]},
      {stage3_10[0]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[1],stage4_11[1],stage4_10[1],stage4_9[6]}
   );
   gpc615_5 gpc5203 (
      {stage3_9[11], stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15]},
      {stage3_10[1]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[2],stage4_11[2],stage4_10[2],stage4_9[7]}
   );
   gpc2135_5 gpc5204 (
      {stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage3_11[18], stage3_11[19], stage3_11[20]},
      {stage3_12[0]},
      {stage3_13[0], stage3_13[1]},
      {stage4_14[0],stage4_13[3],stage4_12[3],stage4_11[3],stage4_10[3]}
   );
   gpc2135_5 gpc5205 (
      {stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage3_12[1]},
      {stage3_13[2], stage3_13[3]},
      {stage4_14[1],stage4_13[4],stage4_12[4],stage4_11[4],stage4_10[4]}
   );
   gpc117_4 gpc5206 (
      {stage3_10[12], stage3_10[13], stage3_10[14], stage3_10[15], stage3_10[16], stage3_10[17], stage3_10[18]},
      {stage3_11[24]},
      {stage3_12[2]},
      {stage4_13[5],stage4_12[5],stage4_11[5],stage4_10[5]}
   );
   gpc117_4 gpc5207 (
      {stage3_10[19], stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage3_11[25]},
      {stage3_12[3]},
      {stage4_13[6],stage4_12[6],stage4_11[6],stage4_10[6]}
   );
   gpc606_5 gpc5208 (
      {stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[2],stage4_13[7],stage4_12[7]}
   );
   gpc606_5 gpc5209 (
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[1],stage4_14[3],stage4_13[8],stage4_12[8]}
   );
   gpc606_5 gpc5210 (
      {stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[2],stage4_15[2],stage4_14[4],stage4_13[9]}
   );
   gpc606_5 gpc5211 (
      {stage3_13[10], stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15]},
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11]},
      {stage4_17[1],stage4_16[3],stage4_15[3],stage4_14[5],stage4_13[10]}
   );
   gpc606_5 gpc5212 (
      {stage3_13[16], stage3_13[17], stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21]},
      {stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17]},
      {stage4_17[2],stage4_16[4],stage4_15[4],stage4_14[6],stage4_13[11]}
   );
   gpc117_4 gpc5213 (
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17], stage3_14[18]},
      {stage3_15[18]},
      {stage3_16[0]},
      {stage4_17[3],stage4_16[5],stage4_15[5],stage4_14[7]}
   );
   gpc615_5 gpc5214 (
      {stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage3_15[19]},
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage4_18[0],stage4_17[4],stage4_16[6],stage4_15[6],stage4_14[8]}
   );
   gpc615_5 gpc5215 (
      {stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24]},
      {stage3_16[7]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[1],stage4_17[5],stage4_16[7],stage4_15[7]}
   );
   gpc615_5 gpc5216 (
      {stage3_15[25], stage3_15[26], stage3_15[27], stage3_15[28], stage3_15[29]},
      {stage3_16[8]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[2],stage4_17[6],stage4_16[8],stage4_15[8]}
   );
   gpc615_5 gpc5217 (
      {stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33], stage3_15[34]},
      {stage3_16[9]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[3],stage4_17[7],stage4_16[9],stage4_15[9]}
   );
   gpc615_5 gpc5218 (
      {stage3_15[35], stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39]},
      {stage3_16[10]},
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage4_19[3],stage4_18[4],stage4_17[8],stage4_16[10],stage4_15[10]}
   );
   gpc615_5 gpc5219 (
      {stage3_16[11], stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15]},
      {stage3_17[24]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[4],stage4_18[5],stage4_17[9],stage4_16[11]}
   );
   gpc615_5 gpc5220 (
      {stage3_16[16], stage3_16[17], stage3_16[18], stage3_16[19], 1'b0},
      {stage3_17[25]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[5],stage4_18[6],stage4_17[10],stage4_16[12]}
   );
   gpc615_5 gpc5221 (
      {stage3_18[12], stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16]},
      {stage3_19[0]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[0],stage4_20[2],stage4_19[6],stage4_18[7]}
   );
   gpc615_5 gpc5222 (
      {stage3_18[17], stage3_18[18], stage3_18[19], stage3_18[20], stage3_18[21]},
      {stage3_19[1]},
      {stage3_20[6], stage3_20[7], stage3_20[8], stage3_20[9], stage3_20[10], stage3_20[11]},
      {stage4_22[1],stage4_21[1],stage4_20[3],stage4_19[7],stage4_18[8]}
   );
   gpc615_5 gpc5223 (
      {stage3_18[22], stage3_18[23], stage3_18[24], stage3_18[25], stage3_18[26]},
      {stage3_19[2]},
      {stage3_20[12], stage3_20[13], stage3_20[14], stage3_20[15], stage3_20[16], stage3_20[17]},
      {stage4_22[2],stage4_21[2],stage4_20[4],stage4_19[8],stage4_18[9]}
   );
   gpc215_4 gpc5224 (
      {stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6], stage3_19[7]},
      {stage3_20[18]},
      {stage3_21[0], stage3_21[1]},
      {stage4_22[3],stage4_21[3],stage4_20[5],stage4_19[9]}
   );
   gpc223_4 gpc5225 (
      {stage3_19[8], stage3_19[9], stage3_19[10]},
      {stage3_20[19], stage3_20[20]},
      {stage3_21[2], stage3_21[3]},
      {stage4_22[4],stage4_21[4],stage4_20[6],stage4_19[10]}
   );
   gpc207_4 gpc5226 (
      {stage3_19[11], stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage3_21[4], stage3_21[5]},
      {stage4_22[5],stage4_21[5],stage4_20[7],stage4_19[11]}
   );
   gpc615_5 gpc5227 (
      {stage3_19[18], stage3_19[19], stage3_19[20], stage3_19[21], stage3_19[22]},
      {stage3_20[21]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[0],stage4_22[6],stage4_21[6],stage4_20[8],stage4_19[12]}
   );
   gpc615_5 gpc5228 (
      {stage3_19[23], stage3_19[24], stage3_19[25], stage3_19[26], stage3_19[27]},
      {stage3_20[22]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[1],stage4_22[7],stage4_21[7],stage4_20[9],stage4_19[13]}
   );
   gpc606_5 gpc5229 (
      {stage3_21[18], stage3_21[19], stage3_21[20], stage3_21[21], stage3_21[22], stage3_21[23]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[0],stage4_23[2],stage4_22[8],stage4_21[8]}
   );
   gpc2135_5 gpc5230 (
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4]},
      {stage3_23[6], stage3_23[7], stage3_23[8]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1]},
      {stage4_26[0],stage4_25[1],stage4_24[1],stage4_23[3],stage4_22[9]}
   );
   gpc2135_5 gpc5231 (
      {stage3_22[5], stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9]},
      {stage3_23[9], stage3_23[10], stage3_23[11]},
      {stage3_24[1]},
      {stage3_25[2], stage3_25[3]},
      {stage4_26[1],stage4_25[2],stage4_24[2],stage4_23[4],stage4_22[10]}
   );
   gpc615_5 gpc5232 (
      {stage3_22[10], stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14]},
      {stage3_23[12]},
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6], stage3_24[7]},
      {stage4_26[2],stage4_25[3],stage4_24[3],stage4_23[5],stage4_22[11]}
   );
   gpc615_5 gpc5233 (
      {stage3_22[15], stage3_22[16], stage3_22[17], stage3_22[18], stage3_22[19]},
      {stage3_23[13]},
      {stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11], stage3_24[12], stage3_24[13]},
      {stage4_26[3],stage4_25[4],stage4_24[4],stage4_23[6],stage4_22[12]}
   );
   gpc615_5 gpc5234 (
      {stage3_22[20], stage3_22[21], stage3_22[22], stage3_22[23], stage3_22[24]},
      {stage3_23[14]},
      {stage3_24[14], stage3_24[15], stage3_24[16], stage3_24[17], stage3_24[18], stage3_24[19]},
      {stage4_26[4],stage4_25[5],stage4_24[5],stage4_23[7],stage4_22[13]}
   );
   gpc615_5 gpc5235 (
      {stage3_22[25], stage3_22[26], stage3_22[27], stage3_22[28], 1'b0},
      {stage3_23[15]},
      {stage3_24[20], stage3_24[21], stage3_24[22], stage3_24[23], stage3_24[24], stage3_24[25]},
      {stage4_26[5],stage4_25[6],stage4_24[6],stage4_23[8],stage4_22[14]}
   );
   gpc1163_5 gpc5236 (
      {stage3_25[4], stage3_25[5], stage3_25[6]},
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4], stage3_26[5]},
      {stage3_27[0]},
      {stage3_28[0]},
      {stage4_29[0],stage4_28[0],stage4_27[0],stage4_26[6],stage4_25[7]}
   );
   gpc1163_5 gpc5237 (
      {stage3_25[7], stage3_25[8], stage3_25[9]},
      {stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage3_27[1]},
      {stage3_28[1]},
      {stage4_29[1],stage4_28[1],stage4_27[1],stage4_26[7],stage4_25[8]}
   );
   gpc1163_5 gpc5238 (
      {stage3_25[10], stage3_25[11], stage3_25[12]},
      {stage3_26[12], stage3_26[13], stage3_26[14], stage3_26[15], stage3_26[16], stage3_26[17]},
      {stage3_27[2]},
      {stage3_28[2]},
      {stage4_29[2],stage4_28[2],stage4_27[2],stage4_26[8],stage4_25[9]}
   );
   gpc1163_5 gpc5239 (
      {stage3_25[13], stage3_25[14], stage3_25[15]},
      {stage3_26[18], stage3_26[19], stage3_26[20], stage3_26[21], stage3_26[22], stage3_26[23]},
      {stage3_27[3]},
      {stage3_28[3]},
      {stage4_29[3],stage4_28[3],stage4_27[3],stage4_26[9],stage4_25[10]}
   );
   gpc606_5 gpc5240 (
      {stage3_25[16], stage3_25[17], stage3_25[18], stage3_25[19], stage3_25[20], stage3_25[21]},
      {stage3_27[4], stage3_27[5], stage3_27[6], stage3_27[7], stage3_27[8], stage3_27[9]},
      {stage4_29[4],stage4_28[4],stage4_27[4],stage4_26[10],stage4_25[11]}
   );
   gpc606_5 gpc5241 (
      {stage3_25[22], stage3_25[23], stage3_25[24], stage3_25[25], stage3_25[26], stage3_25[27]},
      {stage3_27[10], stage3_27[11], stage3_27[12], stage3_27[13], stage3_27[14], stage3_27[15]},
      {stage4_29[5],stage4_28[5],stage4_27[5],stage4_26[11],stage4_25[12]}
   );
   gpc606_5 gpc5242 (
      {stage3_25[28], stage3_25[29], stage3_25[30], stage3_25[31], stage3_25[32], stage3_25[33]},
      {stage3_27[16], stage3_27[17], stage3_27[18], stage3_27[19], stage3_27[20], stage3_27[21]},
      {stage4_29[6],stage4_28[6],stage4_27[6],stage4_26[12],stage4_25[13]}
   );
   gpc606_5 gpc5243 (
      {stage3_28[4], stage3_28[5], stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage4_32[0],stage4_31[0],stage4_30[0],stage4_29[7],stage4_28[7]}
   );
   gpc606_5 gpc5244 (
      {stage3_28[10], stage3_28[11], stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15]},
      {stage3_30[6], stage3_30[7], stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11]},
      {stage4_32[1],stage4_31[1],stage4_30[1],stage4_29[8],stage4_28[8]}
   );
   gpc606_5 gpc5245 (
      {stage3_28[16], stage3_28[17], stage3_28[18], stage3_28[19], stage3_28[20], stage3_28[21]},
      {stage3_30[12], stage3_30[13], stage3_30[14], stage3_30[15], stage3_30[16], stage3_30[17]},
      {stage4_32[2],stage4_31[2],stage4_30[2],stage4_29[9],stage4_28[9]}
   );
   gpc606_5 gpc5246 (
      {stage3_28[22], stage3_28[23], stage3_28[24], stage3_28[25], stage3_28[26], stage3_28[27]},
      {stage3_30[18], stage3_30[19], stage3_30[20], stage3_30[21], stage3_30[22], stage3_30[23]},
      {stage4_32[3],stage4_31[3],stage4_30[3],stage4_29[10],stage4_28[10]}
   );
   gpc606_5 gpc5247 (
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5]},
      {stage4_33[0],stage4_32[4],stage4_31[4],stage4_30[4],stage4_29[11]}
   );
   gpc606_5 gpc5248 (
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_31[6], stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11]},
      {stage4_33[1],stage4_32[5],stage4_31[5],stage4_30[5],stage4_29[12]}
   );
   gpc606_5 gpc5249 (
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_31[12], stage3_31[13], stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17]},
      {stage4_33[2],stage4_32[6],stage4_31[6],stage4_30[6],stage4_29[13]}
   );
   gpc606_5 gpc5250 (
      {stage3_29[18], stage3_29[19], stage3_29[20], stage3_29[21], stage3_29[22], stage3_29[23]},
      {stage3_31[18], stage3_31[19], stage3_31[20], stage3_31[21], stage3_31[22], stage3_31[23]},
      {stage4_33[3],stage4_32[7],stage4_31[7],stage4_30[7],stage4_29[14]}
   );
   gpc606_5 gpc5251 (
      {stage3_29[24], stage3_29[25], stage3_29[26], stage3_29[27], stage3_29[28], stage3_29[29]},
      {stage3_31[24], stage3_31[25], stage3_31[26], stage3_31[27], stage3_31[28], stage3_31[29]},
      {stage4_33[4],stage4_32[8],stage4_31[8],stage4_30[8],stage4_29[15]}
   );
   gpc606_5 gpc5252 (
      {stage3_29[30], stage3_29[31], stage3_29[32], stage3_29[33], stage3_29[34], 1'b0},
      {stage3_31[30], stage3_31[31], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage4_33[5],stage4_32[9],stage4_31[9],stage4_30[9],stage4_29[16]}
   );
   gpc606_5 gpc5253 (
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[6],stage4_32[10]}
   );
   gpc606_5 gpc5254 (
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[1],stage4_34[1],stage4_33[7],stage4_32[11]}
   );
   gpc606_5 gpc5255 (
      {stage3_32[12], stage3_32[13], stage3_32[14], stage3_32[15], stage3_32[16], stage3_32[17]},
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage4_36[2],stage4_35[2],stage4_34[2],stage4_33[8],stage4_32[12]}
   );
   gpc606_5 gpc5256 (
      {stage3_32[18], stage3_32[19], stage3_32[20], stage3_32[21], stage3_32[22], stage3_32[23]},
      {stage3_34[18], stage3_34[19], stage3_34[20], stage3_34[21], stage3_34[22], stage3_34[23]},
      {stage4_36[3],stage4_35[3],stage4_34[3],stage4_33[9],stage4_32[13]}
   );
   gpc606_5 gpc5257 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5]},
      {stage4_37[0],stage4_36[4],stage4_35[4],stage4_34[4],stage4_33[10]}
   );
   gpc606_5 gpc5258 (
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_35[6], stage3_35[7], stage3_35[8], stage3_35[9], stage3_35[10], stage3_35[11]},
      {stage4_37[1],stage4_36[5],stage4_35[5],stage4_34[5],stage4_33[11]}
   );
   gpc606_5 gpc5259 (
      {stage3_33[12], stage3_33[13], stage3_33[14], stage3_33[15], stage3_33[16], stage3_33[17]},
      {stage3_35[12], stage3_35[13], stage3_35[14], stage3_35[15], stage3_35[16], stage3_35[17]},
      {stage4_37[2],stage4_36[6],stage4_35[6],stage4_34[6],stage4_33[12]}
   );
   gpc606_5 gpc5260 (
      {stage3_33[18], stage3_33[19], stage3_33[20], stage3_33[21], stage3_33[22], stage3_33[23]},
      {stage3_35[18], stage3_35[19], stage3_35[20], stage3_35[21], stage3_35[22], stage3_35[23]},
      {stage4_37[3],stage4_36[7],stage4_35[7],stage4_34[7],stage4_33[13]}
   );
   gpc606_5 gpc5261 (
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3], stage3_36[4], stage3_36[5]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5]},
      {stage4_40[0],stage4_39[0],stage4_38[0],stage4_37[4],stage4_36[8]}
   );
   gpc606_5 gpc5262 (
      {stage3_36[6], stage3_36[7], stage3_36[8], stage3_36[9], stage3_36[10], stage3_36[11]},
      {stage3_38[6], stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11]},
      {stage4_40[1],stage4_39[1],stage4_38[1],stage4_37[5],stage4_36[9]}
   );
   gpc606_5 gpc5263 (
      {stage3_36[12], stage3_36[13], stage3_36[14], stage3_36[15], stage3_36[16], stage3_36[17]},
      {stage3_38[12], stage3_38[13], stage3_38[14], stage3_38[15], stage3_38[16], stage3_38[17]},
      {stage4_40[2],stage4_39[2],stage4_38[2],stage4_37[6],stage4_36[10]}
   );
   gpc606_5 gpc5264 (
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4], stage3_37[5]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[3],stage4_39[3],stage4_38[3],stage4_37[7]}
   );
   gpc606_5 gpc5265 (
      {stage3_37[6], stage3_37[7], stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11]},
      {stage3_39[6], stage3_39[7], stage3_39[8], stage3_39[9], stage3_39[10], stage3_39[11]},
      {stage4_41[1],stage4_40[4],stage4_39[4],stage4_38[4],stage4_37[8]}
   );
   gpc615_5 gpc5266 (
      {stage3_37[12], stage3_37[13], stage3_37[14], stage3_37[15], stage3_37[16]},
      {stage3_38[18]},
      {stage3_39[12], stage3_39[13], stage3_39[14], stage3_39[15], stage3_39[16], stage3_39[17]},
      {stage4_41[2],stage4_40[5],stage4_39[5],stage4_38[5],stage4_37[9]}
   );
   gpc615_5 gpc5267 (
      {stage3_38[19], stage3_38[20], stage3_38[21], stage3_38[22], 1'b0},
      {stage3_39[18]},
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage4_42[0],stage4_41[3],stage4_40[6],stage4_39[6],stage4_38[6]}
   );
   gpc606_5 gpc5268 (
      {stage3_39[19], stage3_39[20], stage3_39[21], stage3_39[22], stage3_39[23], stage3_39[24]},
      {stage3_41[0], stage3_41[1], stage3_41[2], stage3_41[3], stage3_41[4], stage3_41[5]},
      {stage4_43[0],stage4_42[1],stage4_41[4],stage4_40[7],stage4_39[7]}
   );
   gpc606_5 gpc5269 (
      {stage3_39[25], stage3_39[26], stage3_39[27], stage3_39[28], stage3_39[29], stage3_39[30]},
      {stage3_41[6], stage3_41[7], stage3_41[8], stage3_41[9], stage3_41[10], stage3_41[11]},
      {stage4_43[1],stage4_42[2],stage4_41[5],stage4_40[8],stage4_39[8]}
   );
   gpc606_5 gpc5270 (
      {stage3_40[6], stage3_40[7], stage3_40[8], stage3_40[9], stage3_40[10], stage3_40[11]},
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5]},
      {stage4_44[0],stage4_43[2],stage4_42[3],stage4_41[6],stage4_40[9]}
   );
   gpc606_5 gpc5271 (
      {stage3_40[12], stage3_40[13], stage3_40[14], stage3_40[15], stage3_40[16], stage3_40[17]},
      {stage3_42[6], stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11]},
      {stage4_44[1],stage4_43[3],stage4_42[4],stage4_41[7],stage4_40[10]}
   );
   gpc606_5 gpc5272 (
      {stage3_40[18], stage3_40[19], stage3_40[20], stage3_40[21], stage3_40[22], stage3_40[23]},
      {stage3_42[12], stage3_42[13], stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17]},
      {stage4_44[2],stage4_43[4],stage4_42[5],stage4_41[8],stage4_40[11]}
   );
   gpc606_5 gpc5273 (
      {stage3_40[24], stage3_40[25], stage3_40[26], stage3_40[27], stage3_40[28], stage3_40[29]},
      {stage3_42[18], stage3_42[19], stage3_42[20], stage3_42[21], stage3_42[22], stage3_42[23]},
      {stage4_44[3],stage4_43[5],stage4_42[6],stage4_41[9],stage4_40[12]}
   );
   gpc606_5 gpc5274 (
      {stage3_41[12], stage3_41[13], stage3_41[14], stage3_41[15], stage3_41[16], stage3_41[17]},
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4], stage3_43[5]},
      {stage4_45[0],stage4_44[4],stage4_43[6],stage4_42[7],stage4_41[10]}
   );
   gpc606_5 gpc5275 (
      {stage3_41[18], stage3_41[19], stage3_41[20], stage3_41[21], stage3_41[22], stage3_41[23]},
      {stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9], stage3_43[10], stage3_43[11]},
      {stage4_45[1],stage4_44[5],stage4_43[7],stage4_42[8],stage4_41[11]}
   );
   gpc606_5 gpc5276 (
      {stage3_43[12], stage3_43[13], stage3_43[14], stage3_43[15], stage3_43[16], stage3_43[17]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[0],stage4_45[2],stage4_44[6],stage4_43[8]}
   );
   gpc606_5 gpc5277 (
      {stage3_43[18], stage3_43[19], stage3_43[20], stage3_43[21], stage3_43[22], stage3_43[23]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage4_47[1],stage4_46[1],stage4_45[3],stage4_44[7],stage4_43[9]}
   );
   gpc606_5 gpc5278 (
      {stage3_43[24], stage3_43[25], stage3_43[26], stage3_43[27], stage3_43[28], stage3_43[29]},
      {stage3_45[12], stage3_45[13], stage3_45[14], stage3_45[15], stage3_45[16], stage3_45[17]},
      {stage4_47[2],stage4_46[2],stage4_45[4],stage4_44[8],stage4_43[10]}
   );
   gpc606_5 gpc5279 (
      {stage3_44[0], stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage3_46[0], stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage4_48[0],stage4_47[3],stage4_46[3],stage4_45[5],stage4_44[9]}
   );
   gpc615_5 gpc5280 (
      {stage3_44[6], stage3_44[7], stage3_44[8], stage3_44[9], stage3_44[10]},
      {stage3_45[18]},
      {stage3_46[6], stage3_46[7], stage3_46[8], stage3_46[9], stage3_46[10], stage3_46[11]},
      {stage4_48[1],stage4_47[4],stage4_46[4],stage4_45[6],stage4_44[10]}
   );
   gpc615_5 gpc5281 (
      {stage3_44[11], stage3_44[12], stage3_44[13], stage3_44[14], stage3_44[15]},
      {stage3_45[19]},
      {stage3_46[12], stage3_46[13], stage3_46[14], stage3_46[15], stage3_46[16], stage3_46[17]},
      {stage4_48[2],stage4_47[5],stage4_46[5],stage4_45[7],stage4_44[11]}
   );
   gpc615_5 gpc5282 (
      {stage3_44[16], stage3_44[17], stage3_44[18], stage3_44[19], stage3_44[20]},
      {stage3_45[20]},
      {stage3_46[18], stage3_46[19], stage3_46[20], stage3_46[21], stage3_46[22], stage3_46[23]},
      {stage4_48[3],stage4_47[6],stage4_46[6],stage4_45[8],stage4_44[12]}
   );
   gpc606_5 gpc5283 (
      {stage3_45[21], stage3_45[22], stage3_45[23], stage3_45[24], stage3_45[25], stage3_45[26]},
      {stage3_47[0], stage3_47[1], stage3_47[2], stage3_47[3], stage3_47[4], stage3_47[5]},
      {stage4_49[0],stage4_48[4],stage4_47[7],stage4_46[7],stage4_45[9]}
   );
   gpc606_5 gpc5284 (
      {stage3_45[27], stage3_45[28], stage3_45[29], stage3_45[30], stage3_45[31], stage3_45[32]},
      {stage3_47[6], stage3_47[7], stage3_47[8], stage3_47[9], stage3_47[10], stage3_47[11]},
      {stage4_49[1],stage4_48[5],stage4_47[8],stage4_46[8],stage4_45[10]}
   );
   gpc606_5 gpc5285 (
      {stage3_45[33], stage3_45[34], stage3_45[35], stage3_45[36], stage3_45[37], stage3_45[38]},
      {stage3_47[12], stage3_47[13], stage3_47[14], stage3_47[15], stage3_47[16], stage3_47[17]},
      {stage4_49[2],stage4_48[6],stage4_47[9],stage4_46[9],stage4_45[11]}
   );
   gpc1406_5 gpc5286 (
      {stage3_46[24], stage3_46[25], stage3_46[26], stage3_46[27], stage3_46[28], stage3_46[29]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3]},
      {stage3_49[0]},
      {stage4_50[0],stage4_49[3],stage4_48[7],stage4_47[10],stage4_46[10]}
   );
   gpc207_4 gpc5287 (
      {stage3_46[30], stage3_46[31], stage3_46[32], stage3_46[33], stage3_46[34], stage3_46[35], stage3_46[36]},
      {stage3_48[4], stage3_48[5]},
      {stage4_49[4],stage4_48[8],stage4_47[11],stage4_46[11]}
   );
   gpc615_5 gpc5288 (
      {stage3_47[18], stage3_47[19], stage3_47[20], stage3_47[21], stage3_47[22]},
      {stage3_48[6]},
      {stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5], stage3_49[6]},
      {stage4_51[0],stage4_50[1],stage4_49[5],stage4_48[9],stage4_47[12]}
   );
   gpc615_5 gpc5289 (
      {stage3_47[23], stage3_47[24], stage3_47[25], stage3_47[26], stage3_47[27]},
      {stage3_48[7]},
      {stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11], stage3_49[12]},
      {stage4_51[1],stage4_50[2],stage4_49[6],stage4_48[10],stage4_47[13]}
   );
   gpc615_5 gpc5290 (
      {stage3_47[28], stage3_47[29], stage3_47[30], stage3_47[31], stage3_47[32]},
      {stage3_48[8]},
      {stage3_49[13], stage3_49[14], stage3_49[15], stage3_49[16], stage3_49[17], stage3_49[18]},
      {stage4_51[2],stage4_50[3],stage4_49[7],stage4_48[11],stage4_47[14]}
   );
   gpc135_4 gpc5291 (
      {stage3_48[9], stage3_48[10], stage3_48[11], stage3_48[12], stage3_48[13]},
      {stage3_49[19], stage3_49[20], stage3_49[21]},
      {stage3_50[0]},
      {stage4_51[3],stage4_50[4],stage4_49[8],stage4_48[12]}
   );
   gpc135_4 gpc5292 (
      {stage3_48[14], stage3_48[15], stage3_48[16], stage3_48[17], stage3_48[18]},
      {stage3_49[22], stage3_49[23], stage3_49[24]},
      {stage3_50[1]},
      {stage4_51[4],stage4_50[5],stage4_49[9],stage4_48[13]}
   );
   gpc135_4 gpc5293 (
      {stage3_48[19], stage3_48[20], stage3_48[21], stage3_48[22], stage3_48[23]},
      {stage3_49[25], stage3_49[26], stage3_49[27]},
      {stage3_50[2]},
      {stage4_51[5],stage4_50[6],stage4_49[10],stage4_48[14]}
   );
   gpc606_5 gpc5294 (
      {stage3_49[28], stage3_49[29], stage3_49[30], stage3_49[31], stage3_49[32], stage3_49[33]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[0],stage4_51[6],stage4_50[7],stage4_49[11]}
   );
   gpc606_5 gpc5295 (
      {stage3_49[34], stage3_49[35], stage3_49[36], stage3_49[37], stage3_49[38], stage3_49[39]},
      {stage3_51[6], stage3_51[7], stage3_51[8], stage3_51[9], stage3_51[10], stage3_51[11]},
      {stage4_53[1],stage4_52[1],stage4_51[7],stage4_50[8],stage4_49[12]}
   );
   gpc606_5 gpc5296 (
      {stage3_49[40], stage3_49[41], stage3_49[42], stage3_49[43], stage3_49[44], stage3_49[45]},
      {stage3_51[12], stage3_51[13], stage3_51[14], stage3_51[15], stage3_51[16], stage3_51[17]},
      {stage4_53[2],stage4_52[2],stage4_51[8],stage4_50[9],stage4_49[13]}
   );
   gpc615_5 gpc5297 (
      {stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6], stage3_50[7]},
      {stage3_51[18]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[3],stage4_52[3],stage4_51[9],stage4_50[10]}
   );
   gpc615_5 gpc5298 (
      {stage3_50[8], stage3_50[9], stage3_50[10], stage3_50[11], stage3_50[12]},
      {stage3_51[19]},
      {stage3_52[6], stage3_52[7], stage3_52[8], stage3_52[9], stage3_52[10], stage3_52[11]},
      {stage4_54[1],stage4_53[4],stage4_52[4],stage4_51[10],stage4_50[11]}
   );
   gpc615_5 gpc5299 (
      {stage3_50[13], stage3_50[14], stage3_50[15], stage3_50[16], stage3_50[17]},
      {stage3_51[20]},
      {stage3_52[12], stage3_52[13], stage3_52[14], stage3_52[15], stage3_52[16], stage3_52[17]},
      {stage4_54[2],stage4_53[5],stage4_52[5],stage4_51[11],stage4_50[12]}
   );
   gpc615_5 gpc5300 (
      {stage3_50[18], stage3_50[19], stage3_50[20], stage3_50[21], stage3_50[22]},
      {stage3_51[21]},
      {stage3_52[18], stage3_52[19], stage3_52[20], stage3_52[21], stage3_52[22], stage3_52[23]},
      {stage4_54[3],stage4_53[6],stage4_52[6],stage4_51[12],stage4_50[13]}
   );
   gpc615_5 gpc5301 (
      {stage3_50[23], stage3_50[24], stage3_50[25], stage3_50[26], stage3_50[27]},
      {stage3_51[22]},
      {stage3_52[24], stage3_52[25], stage3_52[26], stage3_52[27], stage3_52[28], stage3_52[29]},
      {stage4_54[4],stage4_53[7],stage4_52[7],stage4_51[13],stage4_50[14]}
   );
   gpc215_4 gpc5302 (
      {stage3_51[23], stage3_51[24], stage3_51[25], stage3_51[26], stage3_51[27]},
      {stage3_52[30]},
      {stage3_53[0], stage3_53[1]},
      {stage4_54[5],stage4_53[8],stage4_52[8],stage4_51[14]}
   );
   gpc215_4 gpc5303 (
      {stage3_51[28], stage3_51[29], stage3_51[30], stage3_51[31], stage3_51[32]},
      {stage3_52[31]},
      {stage3_53[2], stage3_53[3]},
      {stage4_54[6],stage4_53[9],stage4_52[9],stage4_51[15]}
   );
   gpc606_5 gpc5304 (
      {stage3_51[33], stage3_51[34], stage3_51[35], stage3_51[36], stage3_51[37], stage3_51[38]},
      {stage3_53[4], stage3_53[5], stage3_53[6], stage3_53[7], stage3_53[8], stage3_53[9]},
      {stage4_55[0],stage4_54[7],stage4_53[10],stage4_52[10],stage4_51[16]}
   );
   gpc615_5 gpc5305 (
      {stage3_51[39], stage3_51[40], stage3_51[41], stage3_51[42], stage3_51[43]},
      {stage3_52[32]},
      {stage3_53[10], stage3_53[11], stage3_53[12], stage3_53[13], stage3_53[14], stage3_53[15]},
      {stage4_55[1],stage4_54[8],stage4_53[11],stage4_52[11],stage4_51[17]}
   );
   gpc623_5 gpc5306 (
      {stage3_51[44], stage3_51[45], stage3_51[46]},
      {stage3_52[33], stage3_52[34]},
      {stage3_53[16], stage3_53[17], stage3_53[18], stage3_53[19], stage3_53[20], stage3_53[21]},
      {stage4_55[2],stage4_54[9],stage4_53[12],stage4_52[12],stage4_51[18]}
   );
   gpc606_5 gpc5307 (
      {stage3_52[35], stage3_52[36], stage3_52[37], stage3_52[38], stage3_52[39], 1'b0},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage4_56[0],stage4_55[3],stage4_54[10],stage4_53[13],stage4_52[13]}
   );
   gpc606_5 gpc5308 (
      {stage3_53[22], stage3_53[23], stage3_53[24], stage3_53[25], stage3_53[26], stage3_53[27]},
      {stage3_55[0], stage3_55[1], stage3_55[2], stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage4_57[0],stage4_56[1],stage4_55[4],stage4_54[11],stage4_53[14]}
   );
   gpc2135_5 gpc5309 (
      {stage3_54[6], stage3_54[7], stage3_54[8], stage3_54[9], stage3_54[10]},
      {stage3_55[6], stage3_55[7], stage3_55[8]},
      {stage3_56[0]},
      {stage3_57[0], stage3_57[1]},
      {stage4_58[0],stage4_57[1],stage4_56[2],stage4_55[5],stage4_54[12]}
   );
   gpc615_5 gpc5310 (
      {stage3_54[11], stage3_54[12], stage3_54[13], stage3_54[14], stage3_54[15]},
      {stage3_55[9]},
      {stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5], stage3_56[6]},
      {stage4_58[1],stage4_57[2],stage4_56[3],stage4_55[6],stage4_54[13]}
   );
   gpc615_5 gpc5311 (
      {stage3_54[16], stage3_54[17], stage3_54[18], stage3_54[19], stage3_54[20]},
      {stage3_55[10]},
      {stage3_56[7], stage3_56[8], stage3_56[9], stage3_56[10], stage3_56[11], stage3_56[12]},
      {stage4_58[2],stage4_57[3],stage4_56[4],stage4_55[7],stage4_54[14]}
   );
   gpc615_5 gpc5312 (
      {stage3_54[21], stage3_54[22], stage3_54[23], stage3_54[24], stage3_54[25]},
      {stage3_55[11]},
      {stage3_56[13], stage3_56[14], stage3_56[15], stage3_56[16], stage3_56[17], stage3_56[18]},
      {stage4_58[3],stage4_57[4],stage4_56[5],stage4_55[8],stage4_54[15]}
   );
   gpc615_5 gpc5313 (
      {stage3_55[12], stage3_55[13], stage3_55[14], stage3_55[15], stage3_55[16]},
      {stage3_56[19]},
      {stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5], stage3_57[6], stage3_57[7]},
      {stage4_59[0],stage4_58[4],stage4_57[5],stage4_56[6],stage4_55[9]}
   );
   gpc615_5 gpc5314 (
      {stage3_55[17], stage3_55[18], stage3_55[19], stage3_55[20], stage3_55[21]},
      {stage3_56[20]},
      {stage3_57[8], stage3_57[9], stage3_57[10], stage3_57[11], stage3_57[12], stage3_57[13]},
      {stage4_59[1],stage4_58[5],stage4_57[6],stage4_56[7],stage4_55[10]}
   );
   gpc615_5 gpc5315 (
      {stage3_55[22], stage3_55[23], stage3_55[24], stage3_55[25], stage3_55[26]},
      {stage3_56[21]},
      {stage3_57[14], stage3_57[15], stage3_57[16], stage3_57[17], stage3_57[18], stage3_57[19]},
      {stage4_59[2],stage4_58[6],stage4_57[7],stage4_56[8],stage4_55[11]}
   );
   gpc623_5 gpc5316 (
      {stage3_55[27], stage3_55[28], stage3_55[29]},
      {stage3_56[22], stage3_56[23]},
      {stage3_57[20], stage3_57[21], stage3_57[22], stage3_57[23], stage3_57[24], stage3_57[25]},
      {stage4_59[3],stage4_58[7],stage4_57[8],stage4_56[9],stage4_55[12]}
   );
   gpc615_5 gpc5317 (
      {stage3_57[26], stage3_57[27], stage3_57[28], stage3_57[29], stage3_57[30]},
      {stage3_58[0]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[0],stage4_59[4],stage4_58[8],stage4_57[9]}
   );
   gpc2135_5 gpc5318 (
      {stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5]},
      {stage3_59[6], stage3_59[7], stage3_59[8]},
      {stage3_60[0]},
      {stage3_61[0], stage3_61[1]},
      {stage4_62[0],stage4_61[1],stage4_60[1],stage4_59[5],stage4_58[9]}
   );
   gpc2135_5 gpc5319 (
      {stage3_58[6], stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10]},
      {stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage3_60[1]},
      {stage3_61[2], stage3_61[3]},
      {stage4_62[1],stage4_61[2],stage4_60[2],stage4_59[6],stage4_58[10]}
   );
   gpc2135_5 gpc5320 (
      {stage3_58[11], stage3_58[12], stage3_58[13], stage3_58[14], stage3_58[15]},
      {stage3_59[12], stage3_59[13], stage3_59[14]},
      {stage3_60[2]},
      {stage3_61[4], stage3_61[5]},
      {stage4_62[2],stage4_61[3],stage4_60[3],stage4_59[7],stage4_58[11]}
   );
   gpc606_5 gpc5321 (
      {stage3_58[16], stage3_58[17], stage3_58[18], stage3_58[19], stage3_58[20], stage3_58[21]},
      {stage3_60[3], stage3_60[4], stage3_60[5], stage3_60[6], stage3_60[7], stage3_60[8]},
      {stage4_62[3],stage4_61[4],stage4_60[4],stage4_59[8],stage4_58[12]}
   );
   gpc606_5 gpc5322 (
      {stage3_59[15], stage3_59[16], stage3_59[17], stage3_59[18], stage3_59[19], stage3_59[20]},
      {stage3_61[6], stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11]},
      {stage4_63[0],stage4_62[4],stage4_61[5],stage4_60[5],stage4_59[9]}
   );
   gpc606_5 gpc5323 (
      {stage3_59[21], stage3_59[22], stage3_59[23], stage3_59[24], stage3_59[25], stage3_59[26]},
      {stage3_61[12], stage3_61[13], stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17]},
      {stage4_63[1],stage4_62[5],stage4_61[6],stage4_60[6],stage4_59[10]}
   );
   gpc606_5 gpc5324 (
      {stage3_59[27], stage3_59[28], stage3_59[29], stage3_59[30], stage3_59[31], stage3_59[32]},
      {stage3_61[18], stage3_61[19], stage3_61[20], stage3_61[21], stage3_61[22], stage3_61[23]},
      {stage4_63[2],stage4_62[6],stage4_61[7],stage4_60[7],stage4_59[11]}
   );
   gpc606_5 gpc5325 (
      {stage3_60[9], stage3_60[10], stage3_60[11], stage3_60[12], stage3_60[13], stage3_60[14]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[3],stage4_62[7],stage4_61[8],stage4_60[8]}
   );
   gpc606_5 gpc5326 (
      {stage3_60[15], stage3_60[16], stage3_60[17], stage3_60[18], stage3_60[19], stage3_60[20]},
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage4_64[1],stage4_63[4],stage4_62[8],stage4_61[9],stage4_60[9]}
   );
   gpc606_5 gpc5327 (
      {stage3_60[21], stage3_60[22], stage3_60[23], stage3_60[24], stage3_60[25], stage3_60[26]},
      {stage3_62[12], stage3_62[13], stage3_62[14], stage3_62[15], stage3_62[16], stage3_62[17]},
      {stage4_64[2],stage4_63[5],stage4_62[9],stage4_61[10],stage4_60[10]}
   );
   gpc606_5 gpc5328 (
      {stage3_60[27], stage3_60[28], stage3_60[29], stage3_60[30], stage3_60[31], stage3_60[32]},
      {stage3_62[18], stage3_62[19], stage3_62[20], stage3_62[21], stage3_62[22], stage3_62[23]},
      {stage4_64[3],stage4_63[6],stage4_62[10],stage4_61[11],stage4_60[11]}
   );
   gpc606_5 gpc5329 (
      {stage3_62[24], stage3_62[25], stage3_62[26], stage3_62[27], 1'b0, 1'b0},
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage4_66[0],stage4_65[0],stage4_64[4],stage4_63[7],stage4_62[11]}
   );
   gpc606_5 gpc5330 (
      {stage3_63[0], stage3_63[1], stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[1],stage4_65[1],stage4_64[5],stage4_63[8]}
   );
   gpc606_5 gpc5331 (
      {stage3_63[6], stage3_63[7], stage3_63[8], stage3_63[9], stage3_63[10], stage3_63[11]},
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage4_67[1],stage4_66[2],stage4_65[2],stage4_64[6],stage4_63[9]}
   );
   gpc606_5 gpc5332 (
      {stage3_63[12], stage3_63[13], stage3_63[14], stage3_63[15], stage3_63[16], stage3_63[17]},
      {stage3_65[12], stage3_65[13], stage3_65[14], stage3_65[15], stage3_65[16], stage3_65[17]},
      {stage4_67[2],stage4_66[3],stage4_65[3],stage4_64[7],stage4_63[10]}
   );
   gpc606_5 gpc5333 (
      {stage3_63[18], stage3_63[19], stage3_63[20], stage3_63[21], stage3_63[22], stage3_63[23]},
      {stage3_65[18], stage3_65[19], stage3_65[20], stage3_65[21], stage3_65[22], stage3_65[23]},
      {stage4_67[3],stage4_66[4],stage4_65[4],stage4_64[8],stage4_63[11]}
   );
   gpc606_5 gpc5334 (
      {stage3_63[24], stage3_63[25], stage3_63[26], stage3_63[27], 1'b0, 1'b0},
      {stage3_65[24], stage3_65[25], stage3_65[26], stage3_65[27], 1'b0, 1'b0},
      {stage4_67[4],stage4_66[5],stage4_65[5],stage4_64[9],stage4_63[12]}
   );
   gpc606_5 gpc5335 (
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[5],stage4_66[6],stage4_65[6],stage4_64[10]}
   );
   gpc606_5 gpc5336 (
      {stage3_64[12], stage3_64[13], stage3_64[14], stage3_64[15], stage3_64[16], stage3_64[17]},
      {stage3_66[6], stage3_66[7], stage3_66[8], stage3_66[9], stage3_66[10], stage3_66[11]},
      {stage4_68[1],stage4_67[6],stage4_66[7],stage4_65[7],stage4_64[11]}
   );
   gpc1_1 gpc5337 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc5338 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc5339 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc5340 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc5341 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc5342 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc5343 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc5344 (
      {stage3_0[7]},
      {stage4_0[7]}
   );
   gpc1_1 gpc5345 (
      {stage3_0[8]},
      {stage4_0[8]}
   );
   gpc1_1 gpc5346 (
      {stage3_0[9]},
      {stage4_0[9]}
   );
   gpc1_1 gpc5347 (
      {stage3_0[10]},
      {stage4_0[10]}
   );
   gpc1_1 gpc5348 (
      {stage3_0[11]},
      {stage4_0[11]}
   );
   gpc1_1 gpc5349 (
      {stage3_0[12]},
      {stage4_0[12]}
   );
   gpc1_1 gpc5350 (
      {stage3_0[13]},
      {stage4_0[13]}
   );
   gpc1_1 gpc5351 (
      {stage3_1[8]},
      {stage4_1[2]}
   );
   gpc1_1 gpc5352 (
      {stage3_1[9]},
      {stage4_1[3]}
   );
   gpc1_1 gpc5353 (
      {stage3_1[10]},
      {stage4_1[4]}
   );
   gpc1_1 gpc5354 (
      {stage3_2[14]},
      {stage4_2[3]}
   );
   gpc1_1 gpc5355 (
      {stage3_2[15]},
      {stage4_2[4]}
   );
   gpc1_1 gpc5356 (
      {stage3_2[16]},
      {stage4_2[5]}
   );
   gpc1_1 gpc5357 (
      {stage3_2[17]},
      {stage4_2[6]}
   );
   gpc1_1 gpc5358 (
      {stage3_3[3]},
      {stage4_3[3]}
   );
   gpc1_1 gpc5359 (
      {stage3_3[4]},
      {stage4_3[4]}
   );
   gpc1_1 gpc5360 (
      {stage3_3[5]},
      {stage4_3[5]}
   );
   gpc1_1 gpc5361 (
      {stage3_3[6]},
      {stage4_3[6]}
   );
   gpc1_1 gpc5362 (
      {stage3_3[7]},
      {stage4_3[7]}
   );
   gpc1_1 gpc5363 (
      {stage3_3[8]},
      {stage4_3[8]}
   );
   gpc1_1 gpc5364 (
      {stage3_3[9]},
      {stage4_3[9]}
   );
   gpc1_1 gpc5365 (
      {stage3_3[10]},
      {stage4_3[10]}
   );
   gpc1_1 gpc5366 (
      {stage3_3[11]},
      {stage4_3[11]}
   );
   gpc1_1 gpc5367 (
      {stage3_3[12]},
      {stage4_3[12]}
   );
   gpc1_1 gpc5368 (
      {stage3_3[13]},
      {stage4_3[13]}
   );
   gpc1_1 gpc5369 (
      {stage3_3[14]},
      {stage4_3[14]}
   );
   gpc1_1 gpc5370 (
      {stage3_3[15]},
      {stage4_3[15]}
   );
   gpc1_1 gpc5371 (
      {stage3_3[16]},
      {stage4_3[16]}
   );
   gpc1_1 gpc5372 (
      {stage3_3[17]},
      {stage4_3[17]}
   );
   gpc1_1 gpc5373 (
      {stage3_3[18]},
      {stage4_3[18]}
   );
   gpc1_1 gpc5374 (
      {stage3_4[15]},
      {stage4_4[4]}
   );
   gpc1_1 gpc5375 (
      {stage3_4[16]},
      {stage4_4[5]}
   );
   gpc1_1 gpc5376 (
      {stage3_4[17]},
      {stage4_4[6]}
   );
   gpc1_1 gpc5377 (
      {stage3_4[18]},
      {stage4_4[7]}
   );
   gpc1_1 gpc5378 (
      {stage3_4[19]},
      {stage4_4[8]}
   );
   gpc1_1 gpc5379 (
      {stage3_4[20]},
      {stage4_4[9]}
   );
   gpc1_1 gpc5380 (
      {stage3_5[24]},
      {stage4_5[9]}
   );
   gpc1_1 gpc5381 (
      {stage3_5[25]},
      {stage4_5[10]}
   );
   gpc1_1 gpc5382 (
      {stage3_5[26]},
      {stage4_5[11]}
   );
   gpc1_1 gpc5383 (
      {stage3_5[27]},
      {stage4_5[12]}
   );
   gpc1_1 gpc5384 (
      {stage3_5[28]},
      {stage4_5[13]}
   );
   gpc1_1 gpc5385 (
      {stage3_5[29]},
      {stage4_5[14]}
   );
   gpc1_1 gpc5386 (
      {stage3_5[30]},
      {stage4_5[15]}
   );
   gpc1_1 gpc5387 (
      {stage3_5[31]},
      {stage4_5[16]}
   );
   gpc1_1 gpc5388 (
      {stage3_5[32]},
      {stage4_5[17]}
   );
   gpc1_1 gpc5389 (
      {stage3_5[33]},
      {stage4_5[18]}
   );
   gpc1_1 gpc5390 (
      {stage3_5[34]},
      {stage4_5[19]}
   );
   gpc1_1 gpc5391 (
      {stage3_6[14]},
      {stage4_6[7]}
   );
   gpc1_1 gpc5392 (
      {stage3_6[15]},
      {stage4_6[8]}
   );
   gpc1_1 gpc5393 (
      {stage3_6[16]},
      {stage4_6[9]}
   );
   gpc1_1 gpc5394 (
      {stage3_7[24]},
      {stage4_7[6]}
   );
   gpc1_1 gpc5395 (
      {stage3_7[25]},
      {stage4_7[7]}
   );
   gpc1_1 gpc5396 (
      {stage3_7[26]},
      {stage4_7[8]}
   );
   gpc1_1 gpc5397 (
      {stage3_7[27]},
      {stage4_7[9]}
   );
   gpc1_1 gpc5398 (
      {stage3_8[2]},
      {stage4_8[6]}
   );
   gpc1_1 gpc5399 (
      {stage3_8[3]},
      {stage4_8[7]}
   );
   gpc1_1 gpc5400 (
      {stage3_8[4]},
      {stage4_8[8]}
   );
   gpc1_1 gpc5401 (
      {stage3_8[5]},
      {stage4_8[9]}
   );
   gpc1_1 gpc5402 (
      {stage3_8[6]},
      {stage4_8[10]}
   );
   gpc1_1 gpc5403 (
      {stage3_8[7]},
      {stage4_8[11]}
   );
   gpc1_1 gpc5404 (
      {stage3_8[8]},
      {stage4_8[12]}
   );
   gpc1_1 gpc5405 (
      {stage3_8[9]},
      {stage4_8[13]}
   );
   gpc1_1 gpc5406 (
      {stage3_8[10]},
      {stage4_8[14]}
   );
   gpc1_1 gpc5407 (
      {stage3_8[11]},
      {stage4_8[15]}
   );
   gpc1_1 gpc5408 (
      {stage3_8[12]},
      {stage4_8[16]}
   );
   gpc1_1 gpc5409 (
      {stage3_8[13]},
      {stage4_8[17]}
   );
   gpc1_1 gpc5410 (
      {stage3_8[14]},
      {stage4_8[18]}
   );
   gpc1_1 gpc5411 (
      {stage3_8[15]},
      {stage4_8[19]}
   );
   gpc1_1 gpc5412 (
      {stage3_8[16]},
      {stage4_8[20]}
   );
   gpc1_1 gpc5413 (
      {stage3_8[17]},
      {stage4_8[21]}
   );
   gpc1_1 gpc5414 (
      {stage3_10[26]},
      {stage4_10[7]}
   );
   gpc1_1 gpc5415 (
      {stage3_10[27]},
      {stage4_10[8]}
   );
   gpc1_1 gpc5416 (
      {stage3_10[28]},
      {stage4_10[9]}
   );
   gpc1_1 gpc5417 (
      {stage3_10[29]},
      {stage4_10[10]}
   );
   gpc1_1 gpc5418 (
      {stage3_10[30]},
      {stage4_10[11]}
   );
   gpc1_1 gpc5419 (
      {stage3_10[31]},
      {stage4_10[12]}
   );
   gpc1_1 gpc5420 (
      {stage3_10[32]},
      {stage4_10[13]}
   );
   gpc1_1 gpc5421 (
      {stage3_11[26]},
      {stage4_11[7]}
   );
   gpc1_1 gpc5422 (
      {stage3_11[27]},
      {stage4_11[8]}
   );
   gpc1_1 gpc5423 (
      {stage3_11[28]},
      {stage4_11[9]}
   );
   gpc1_1 gpc5424 (
      {stage3_11[29]},
      {stage4_11[10]}
   );
   gpc1_1 gpc5425 (
      {stage3_11[30]},
      {stage4_11[11]}
   );
   gpc1_1 gpc5426 (
      {stage3_12[16]},
      {stage4_12[9]}
   );
   gpc1_1 gpc5427 (
      {stage3_12[17]},
      {stage4_12[10]}
   );
   gpc1_1 gpc5428 (
      {stage3_12[18]},
      {stage4_12[11]}
   );
   gpc1_1 gpc5429 (
      {stage3_12[19]},
      {stage4_12[12]}
   );
   gpc1_1 gpc5430 (
      {stage3_12[20]},
      {stage4_12[13]}
   );
   gpc1_1 gpc5431 (
      {stage3_12[21]},
      {stage4_12[14]}
   );
   gpc1_1 gpc5432 (
      {stage3_12[22]},
      {stage4_12[15]}
   );
   gpc1_1 gpc5433 (
      {stage3_12[23]},
      {stage4_12[16]}
   );
   gpc1_1 gpc5434 (
      {stage3_12[24]},
      {stage4_12[17]}
   );
   gpc1_1 gpc5435 (
      {stage3_13[22]},
      {stage4_13[12]}
   );
   gpc1_1 gpc5436 (
      {stage3_13[23]},
      {stage4_13[13]}
   );
   gpc1_1 gpc5437 (
      {stage3_14[24]},
      {stage4_14[9]}
   );
   gpc1_1 gpc5438 (
      {stage3_14[25]},
      {stage4_14[10]}
   );
   gpc1_1 gpc5439 (
      {stage3_14[26]},
      {stage4_14[11]}
   );
   gpc1_1 gpc5440 (
      {stage3_15[40]},
      {stage4_15[11]}
   );
   gpc1_1 gpc5441 (
      {stage3_17[26]},
      {stage4_17[11]}
   );
   gpc1_1 gpc5442 (
      {stage3_17[27]},
      {stage4_17[12]}
   );
   gpc1_1 gpc5443 (
      {stage3_17[28]},
      {stage4_17[13]}
   );
   gpc1_1 gpc5444 (
      {stage3_17[29]},
      {stage4_17[14]}
   );
   gpc1_1 gpc5445 (
      {stage3_18[27]},
      {stage4_18[10]}
   );
   gpc1_1 gpc5446 (
      {stage3_20[23]},
      {stage4_20[10]}
   );
   gpc1_1 gpc5447 (
      {stage3_24[26]},
      {stage4_24[7]}
   );
   gpc1_1 gpc5448 (
      {stage3_24[27]},
      {stage4_24[8]}
   );
   gpc1_1 gpc5449 (
      {stage3_24[28]},
      {stage4_24[9]}
   );
   gpc1_1 gpc5450 (
      {stage3_24[29]},
      {stage4_24[10]}
   );
   gpc1_1 gpc5451 (
      {stage3_24[30]},
      {stage4_24[11]}
   );
   gpc1_1 gpc5452 (
      {stage3_28[28]},
      {stage4_28[11]}
   );
   gpc1_1 gpc5453 (
      {stage3_30[24]},
      {stage4_30[10]}
   );
   gpc1_1 gpc5454 (
      {stage3_30[25]},
      {stage4_30[11]}
   );
   gpc1_1 gpc5455 (
      {stage3_32[24]},
      {stage4_32[14]}
   );
   gpc1_1 gpc5456 (
      {stage3_32[25]},
      {stage4_32[15]}
   );
   gpc1_1 gpc5457 (
      {stage3_32[26]},
      {stage4_32[16]}
   );
   gpc1_1 gpc5458 (
      {stage3_32[27]},
      {stage4_32[17]}
   );
   gpc1_1 gpc5459 (
      {stage3_33[24]},
      {stage4_33[14]}
   );
   gpc1_1 gpc5460 (
      {stage3_33[25]},
      {stage4_33[15]}
   );
   gpc1_1 gpc5461 (
      {stage3_33[26]},
      {stage4_33[16]}
   );
   gpc1_1 gpc5462 (
      {stage3_34[24]},
      {stage4_34[8]}
   );
   gpc1_1 gpc5463 (
      {stage3_34[25]},
      {stage4_34[9]}
   );
   gpc1_1 gpc5464 (
      {stage3_34[26]},
      {stage4_34[10]}
   );
   gpc1_1 gpc5465 (
      {stage3_35[24]},
      {stage4_35[8]}
   );
   gpc1_1 gpc5466 (
      {stage3_35[25]},
      {stage4_35[9]}
   );
   gpc1_1 gpc5467 (
      {stage3_35[26]},
      {stage4_35[10]}
   );
   gpc1_1 gpc5468 (
      {stage3_35[27]},
      {stage4_35[11]}
   );
   gpc1_1 gpc5469 (
      {stage3_35[28]},
      {stage4_35[12]}
   );
   gpc1_1 gpc5470 (
      {stage3_35[29]},
      {stage4_35[13]}
   );
   gpc1_1 gpc5471 (
      {stage3_35[30]},
      {stage4_35[14]}
   );
   gpc1_1 gpc5472 (
      {stage3_35[31]},
      {stage4_35[15]}
   );
   gpc1_1 gpc5473 (
      {stage3_35[32]},
      {stage4_35[16]}
   );
   gpc1_1 gpc5474 (
      {stage3_36[18]},
      {stage4_36[11]}
   );
   gpc1_1 gpc5475 (
      {stage3_36[19]},
      {stage4_36[12]}
   );
   gpc1_1 gpc5476 (
      {stage3_37[17]},
      {stage4_37[10]}
   );
   gpc1_1 gpc5477 (
      {stage3_37[18]},
      {stage4_37[11]}
   );
   gpc1_1 gpc5478 (
      {stage3_42[24]},
      {stage4_42[9]}
   );
   gpc1_1 gpc5479 (
      {stage3_42[25]},
      {stage4_42[10]}
   );
   gpc1_1 gpc5480 (
      {stage3_42[26]},
      {stage4_42[11]}
   );
   gpc1_1 gpc5481 (
      {stage3_42[27]},
      {stage4_42[12]}
   );
   gpc1_1 gpc5482 (
      {stage3_42[28]},
      {stage4_42[13]}
   );
   gpc1_1 gpc5483 (
      {stage3_42[29]},
      {stage4_42[14]}
   );
   gpc1_1 gpc5484 (
      {stage3_43[30]},
      {stage4_43[11]}
   );
   gpc1_1 gpc5485 (
      {stage3_43[31]},
      {stage4_43[12]}
   );
   gpc1_1 gpc5486 (
      {stage3_43[32]},
      {stage4_43[13]}
   );
   gpc1_1 gpc5487 (
      {stage3_43[33]},
      {stage4_43[14]}
   );
   gpc1_1 gpc5488 (
      {stage3_43[34]},
      {stage4_43[15]}
   );
   gpc1_1 gpc5489 (
      {stage3_43[35]},
      {stage4_43[16]}
   );
   gpc1_1 gpc5490 (
      {stage3_43[36]},
      {stage4_43[17]}
   );
   gpc1_1 gpc5491 (
      {stage3_43[37]},
      {stage4_43[18]}
   );
   gpc1_1 gpc5492 (
      {stage3_43[38]},
      {stage4_43[19]}
   );
   gpc1_1 gpc5493 (
      {stage3_44[21]},
      {stage4_44[13]}
   );
   gpc1_1 gpc5494 (
      {stage3_46[37]},
      {stage4_46[12]}
   );
   gpc1_1 gpc5495 (
      {stage3_46[38]},
      {stage4_46[13]}
   );
   gpc1_1 gpc5496 (
      {stage3_46[39]},
      {stage4_46[14]}
   );
   gpc1_1 gpc5497 (
      {stage3_49[46]},
      {stage4_49[14]}
   );
   gpc1_1 gpc5498 (
      {stage3_49[47]},
      {stage4_49[15]}
   );
   gpc1_1 gpc5499 (
      {stage3_49[48]},
      {stage4_49[16]}
   );
   gpc1_1 gpc5500 (
      {stage3_49[49]},
      {stage4_49[17]}
   );
   gpc1_1 gpc5501 (
      {stage3_49[50]},
      {stage4_49[18]}
   );
   gpc1_1 gpc5502 (
      {stage3_49[51]},
      {stage4_49[19]}
   );
   gpc1_1 gpc5503 (
      {stage3_49[52]},
      {stage4_49[20]}
   );
   gpc1_1 gpc5504 (
      {stage3_49[53]},
      {stage4_49[21]}
   );
   gpc1_1 gpc5505 (
      {stage3_49[54]},
      {stage4_49[22]}
   );
   gpc1_1 gpc5506 (
      {stage3_49[55]},
      {stage4_49[23]}
   );
   gpc1_1 gpc5507 (
      {stage3_49[56]},
      {stage4_49[24]}
   );
   gpc1_1 gpc5508 (
      {stage3_49[57]},
      {stage4_49[25]}
   );
   gpc1_1 gpc5509 (
      {stage3_49[58]},
      {stage4_49[26]}
   );
   gpc1_1 gpc5510 (
      {stage3_49[59]},
      {stage4_49[27]}
   );
   gpc1_1 gpc5511 (
      {stage3_49[60]},
      {stage4_49[28]}
   );
   gpc1_1 gpc5512 (
      {stage3_49[61]},
      {stage4_49[29]}
   );
   gpc1_1 gpc5513 (
      {stage3_49[62]},
      {stage4_49[30]}
   );
   gpc1_1 gpc5514 (
      {stage3_49[63]},
      {stage4_49[31]}
   );
   gpc1_1 gpc5515 (
      {stage3_49[64]},
      {stage4_49[32]}
   );
   gpc1_1 gpc5516 (
      {stage3_49[65]},
      {stage4_49[33]}
   );
   gpc1_1 gpc5517 (
      {stage3_49[66]},
      {stage4_49[34]}
   );
   gpc1_1 gpc5518 (
      {stage3_49[67]},
      {stage4_49[35]}
   );
   gpc1_1 gpc5519 (
      {stage3_50[28]},
      {stage4_50[15]}
   );
   gpc1_1 gpc5520 (
      {stage3_50[29]},
      {stage4_50[16]}
   );
   gpc1_1 gpc5521 (
      {stage3_51[47]},
      {stage4_51[19]}
   );
   gpc1_1 gpc5522 (
      {stage3_54[26]},
      {stage4_54[16]}
   );
   gpc1_1 gpc5523 (
      {stage3_54[27]},
      {stage4_54[17]}
   );
   gpc1_1 gpc5524 (
      {stage3_56[24]},
      {stage4_56[10]}
   );
   gpc1_1 gpc5525 (
      {stage3_56[25]},
      {stage4_56[11]}
   );
   gpc1_1 gpc5526 (
      {stage3_57[31]},
      {stage4_57[10]}
   );
   gpc1_1 gpc5527 (
      {stage3_57[32]},
      {stage4_57[11]}
   );
   gpc1_1 gpc5528 (
      {stage3_58[22]},
      {stage4_58[13]}
   );
   gpc1_1 gpc5529 (
      {stage3_58[23]},
      {stage4_58[14]}
   );
   gpc1_1 gpc5530 (
      {stage3_58[24]},
      {stage4_58[15]}
   );
   gpc1_1 gpc5531 (
      {stage3_58[25]},
      {stage4_58[16]}
   );
   gpc1_1 gpc5532 (
      {stage3_58[26]},
      {stage4_58[17]}
   );
   gpc1_1 gpc5533 (
      {stage3_58[27]},
      {stage4_58[18]}
   );
   gpc1_1 gpc5534 (
      {stage3_58[28]},
      {stage4_58[19]}
   );
   gpc1_1 gpc5535 (
      {stage3_60[33]},
      {stage4_60[12]}
   );
   gpc1_1 gpc5536 (
      {stage3_60[34]},
      {stage4_60[13]}
   );
   gpc1_1 gpc5537 (
      {stage3_66[12]},
      {stage4_66[8]}
   );
   gpc1_1 gpc5538 (
      {stage3_66[13]},
      {stage4_66[9]}
   );
   gpc1_1 gpc5539 (
      {stage3_66[14]},
      {stage4_66[10]}
   );
   gpc1_1 gpc5540 (
      {stage3_66[15]},
      {stage4_66[11]}
   );
   gpc1_1 gpc5541 (
      {stage3_66[16]},
      {stage4_66[12]}
   );
   gpc1_1 gpc5542 (
      {stage3_66[17]},
      {stage4_66[13]}
   );
   gpc1_1 gpc5543 (
      {stage3_66[18]},
      {stage4_66[14]}
   );
   gpc1_1 gpc5544 (
      {stage3_66[19]},
      {stage4_66[15]}
   );
   gpc1_1 gpc5545 (
      {stage3_66[20]},
      {stage4_66[16]}
   );
   gpc1_1 gpc5546 (
      {stage3_66[21]},
      {stage4_66[17]}
   );
   gpc1_1 gpc5547 (
      {stage3_66[22]},
      {stage4_66[18]}
   );
   gpc1_1 gpc5548 (
      {stage3_66[23]},
      {stage4_66[19]}
   );
   gpc1_1 gpc5549 (
      {stage3_66[24]},
      {stage4_66[20]}
   );
   gpc1_1 gpc5550 (
      {stage3_66[25]},
      {stage4_66[21]}
   );
   gpc1_1 gpc5551 (
      {stage3_66[26]},
      {stage4_66[22]}
   );
   gpc1_1 gpc5552 (
      {stage3_66[27]},
      {stage4_66[23]}
   );
   gpc1_1 gpc5553 (
      {stage3_67[0]},
      {stage4_67[7]}
   );
   gpc1_1 gpc5554 (
      {stage3_67[1]},
      {stage4_67[8]}
   );
   gpc1_1 gpc5555 (
      {stage3_68[0]},
      {stage4_68[2]}
   );
   gpc1_1 gpc5556 (
      {stage3_69[0]},
      {stage4_69[0]}
   );
   gpc2135_5 gpc5557 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4]},
      {stage4_1[0], stage4_1[1], stage4_1[2]},
      {stage4_2[0]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc606_5 gpc5558 (
      {stage4_0[5], stage4_0[6], stage4_0[7], stage4_0[8], stage4_0[9], stage4_0[10]},
      {stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5], stage4_2[6]},
      {stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1],stage5_0[1]}
   );
   gpc2135_5 gpc5559 (
      {stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5], stage4_3[6]},
      {stage4_4[0], stage4_4[1], stage4_4[2]},
      {stage4_5[0]},
      {stage4_6[0], stage4_6[1]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[2],stage5_3[2]}
   );
   gpc615_5 gpc5560 (
      {stage4_3[7], stage4_3[8], stage4_3[9], stage4_3[10], stage4_3[11]},
      {stage4_4[3]},
      {stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6]},
      {stage5_7[1],stage5_6[1],stage5_5[1],stage5_4[3],stage5_3[3]}
   );
   gpc615_5 gpc5561 (
      {stage4_3[12], stage4_3[13], stage4_3[14], stage4_3[15], stage4_3[16]},
      {stage4_4[4]},
      {stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11], stage4_5[12]},
      {stage5_7[2],stage5_6[2],stage5_5[2],stage5_4[4],stage5_3[4]}
   );
   gpc1163_5 gpc5562 (
      {stage4_5[13], stage4_5[14], stage4_5[15]},
      {stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5], stage4_6[6], stage4_6[7]},
      {stage4_7[0]},
      {stage4_8[0]},
      {stage5_9[0],stage5_8[0],stage5_7[3],stage5_6[3],stage5_5[3]}
   );
   gpc117_4 gpc5563 (
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[1]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[1],stage5_8[1],stage5_7[4]}
   );
   gpc117_4 gpc5564 (
      {stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5], stage4_8[6], stage4_8[7], stage4_8[8]},
      {stage4_9[1]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[1],stage5_9[2],stage5_8[2]}
   );
   gpc117_4 gpc5565 (
      {stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12], stage4_8[13], stage4_8[14], stage4_8[15]},
      {stage4_9[2]},
      {stage4_10[1]},
      {stage5_11[1],stage5_10[2],stage5_9[3],stage5_8[3]}
   );
   gpc606_5 gpc5566 (
      {stage4_8[16], stage4_8[17], stage4_8[18], stage4_8[19], stage4_8[20], stage4_8[21]},
      {stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage5_12[0],stage5_11[2],stage5_10[3],stage5_9[4],stage5_8[4]}
   );
   gpc615_5 gpc5567 (
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12]},
      {stage4_11[0]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[0],stage5_12[1],stage5_11[3],stage5_10[4]}
   );
   gpc606_5 gpc5568 (
      {stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[1],stage5_13[1],stage5_12[2],stage5_11[4]}
   );
   gpc606_5 gpc5569 (
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[1],stage5_14[2],stage5_13[2],stage5_12[3]}
   );
   gpc615_5 gpc5570 (
      {stage4_12[12], stage4_12[13], stage4_12[14], stage4_12[15], stage4_12[16]},
      {stage4_13[6]},
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10], stage4_14[11]},
      {stage5_16[1],stage5_15[2],stage5_14[3],stage5_13[3],stage5_12[4]}
   );
   gpc606_5 gpc5571 (
      {stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11], stage4_13[12]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {stage5_17[0],stage5_16[2],stage5_15[3],stage5_14[4],stage5_13[4]}
   );
   gpc615_5 gpc5572 (
      {stage4_15[6], stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10]},
      {stage4_16[0]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[0],stage5_17[1],stage5_16[3],stage5_15[4]}
   );
   gpc207_4 gpc5573 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6], stage4_16[7]},
      {stage4_18[0], stage4_18[1]},
      {stage5_19[1],stage5_18[1],stage5_17[2],stage5_16[4]}
   );
   gpc207_4 gpc5574 (
      {stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11], stage4_16[12], 1'b0, 1'b0},
      {stage4_18[2], stage4_18[3]},
      {stage5_19[2],stage5_18[2],stage5_17[3],stage5_16[5]}
   );
   gpc606_5 gpc5575 (
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[0],stage5_19[3],stage5_18[3],stage5_17[4]}
   );
   gpc615_5 gpc5576 (
      {stage4_18[4], stage4_18[5], stage4_18[6], stage4_18[7], stage4_18[8]},
      {stage4_19[6]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[1],stage5_19[4],stage5_18[4]}
   );
   gpc623_5 gpc5577 (
      {stage4_18[9], stage4_18[10], 1'b0},
      {stage4_19[7], stage4_19[8]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9], stage4_20[10], 1'b0},
      {stage5_22[1],stage5_21[2],stage5_20[2],stage5_19[5],stage5_18[5]}
   );
   gpc135_4 gpc5578 (
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4]},
      {stage4_23[0], stage4_23[1], stage4_23[2]},
      {stage4_24[0]},
      {stage5_25[0],stage5_24[0],stage5_23[0],stage5_22[2]}
   );
   gpc2135_5 gpc5579 (
      {stage4_22[5], stage4_22[6], stage4_22[7], stage4_22[8], stage4_22[9]},
      {stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[1]},
      {stage4_25[0], stage4_25[1]},
      {stage5_26[0],stage5_25[1],stage5_24[1],stage5_23[1],stage5_22[3]}
   );
   gpc2135_5 gpc5580 (
      {stage4_22[10], stage4_22[11], stage4_22[12], stage4_22[13], stage4_22[14]},
      {stage4_23[6], stage4_23[7], stage4_23[8]},
      {stage4_24[2]},
      {stage4_25[2], stage4_25[3]},
      {stage5_26[1],stage5_25[2],stage5_24[2],stage5_23[2],stage5_22[4]}
   );
   gpc606_5 gpc5581 (
      {stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6], stage4_24[7], stage4_24[8]},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage5_28[0],stage5_27[0],stage5_26[2],stage5_25[3],stage5_24[3]}
   );
   gpc23_3 gpc5582 (
      {stage4_25[4], stage4_25[5], stage4_25[6]},
      {stage4_26[6], stage4_26[7]},
      {stage5_27[1],stage5_26[3],stage5_25[4]}
   );
   gpc7_3 gpc5583 (
      {stage4_25[7], stage4_25[8], stage4_25[9], stage4_25[10], stage4_25[11], stage4_25[12], stage4_25[13]},
      {stage5_27[2],stage5_26[4],stage5_25[5]}
   );
   gpc615_5 gpc5584 (
      {stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11], stage4_26[12]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[3],stage5_26[5]}
   );
   gpc1343_5 gpc5585 (
      {stage4_27[1], stage4_27[2], stage4_27[3]},
      {stage4_28[6], stage4_28[7], stage4_28[8], stage4_28[9]},
      {stage4_29[0], stage4_29[1], stage4_29[2]},
      {stage4_30[0]},
      {stage5_31[0],stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[4]}
   );
   gpc1423_5 gpc5586 (
      {stage4_27[4], stage4_27[5], stage4_27[6]},
      {stage4_28[10], stage4_28[11]},
      {stage4_29[3], stage4_29[4], stage4_29[5], stage4_29[6]},
      {stage4_30[1]},
      {stage5_31[1],stage5_30[2],stage5_29[2],stage5_28[3],stage5_27[5]}
   );
   gpc606_5 gpc5587 (
      {stage4_29[7], stage4_29[8], stage4_29[9], stage4_29[10], stage4_29[11], stage4_29[12]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[2],stage5_30[3],stage5_29[3]}
   );
   gpc615_5 gpc5588 (
      {stage4_30[2], stage4_30[3], stage4_30[4], stage4_30[5], stage4_30[6]},
      {stage4_31[6]},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[3],stage5_30[4]}
   );
   gpc615_5 gpc5589 (
      {stage4_30[7], stage4_30[8], stage4_30[9], stage4_30[10], stage4_30[11]},
      {stage4_31[7]},
      {stage4_32[6], stage4_32[7], stage4_32[8], stage4_32[9], stage4_32[10], stage4_32[11]},
      {stage5_34[1],stage5_33[2],stage5_32[2],stage5_31[4],stage5_30[5]}
   );
   gpc606_5 gpc5590 (
      {stage4_32[12], stage4_32[13], stage4_32[14], stage4_32[15], stage4_32[16], stage4_32[17]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[0],stage5_34[2],stage5_33[3],stage5_32[3]}
   );
   gpc606_5 gpc5591 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[1],stage5_35[1],stage5_34[3],stage5_33[4]}
   );
   gpc606_5 gpc5592 (
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_35[6], stage4_35[7], stage4_35[8], stage4_35[9], stage4_35[10], stage4_35[11]},
      {stage5_37[1],stage5_36[2],stage5_35[2],stage5_34[4],stage5_33[5]}
   );
   gpc606_5 gpc5593 (
      {stage4_33[12], stage4_33[13], stage4_33[14], stage4_33[15], stage4_33[16], 1'b0},
      {stage4_35[12], stage4_35[13], stage4_35[14], stage4_35[15], stage4_35[16], 1'b0},
      {stage5_37[2],stage5_36[3],stage5_35[3],stage5_34[5],stage5_33[6]}
   );
   gpc615_5 gpc5594 (
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10]},
      {1'b0},
      {stage4_36[0], stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5]},
      {stage5_38[0],stage5_37[3],stage5_36[4],stage5_35[4],stage5_34[6]}
   );
   gpc606_5 gpc5595 (
      {stage4_36[6], stage4_36[7], stage4_36[8], stage4_36[9], stage4_36[10], stage4_36[11]},
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5]},
      {stage5_40[0],stage5_39[0],stage5_38[1],stage5_37[4],stage5_36[5]}
   );
   gpc606_5 gpc5596 (
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage4_39[0], stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5]},
      {stage5_41[0],stage5_40[1],stage5_39[1],stage5_38[2],stage5_37[5]}
   );
   gpc606_5 gpc5597 (
      {stage4_39[6], stage4_39[7], stage4_39[8], 1'b0, 1'b0, 1'b0},
      {stage4_41[0], stage4_41[1], stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5]},
      {stage5_43[0],stage5_42[0],stage5_41[1],stage5_40[2],stage5_39[2]}
   );
   gpc606_5 gpc5598 (
      {stage4_40[0], stage4_40[1], stage4_40[2], stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[1],stage5_42[1],stage5_41[2],stage5_40[3]}
   );
   gpc606_5 gpc5599 (
      {stage4_40[6], stage4_40[7], stage4_40[8], stage4_40[9], stage4_40[10], stage4_40[11]},
      {stage4_42[6], stage4_42[7], stage4_42[8], stage4_42[9], stage4_42[10], stage4_42[11]},
      {stage5_44[1],stage5_43[2],stage5_42[2],stage5_41[3],stage5_40[4]}
   );
   gpc606_5 gpc5600 (
      {stage4_41[6], stage4_41[7], stage4_41[8], stage4_41[9], stage4_41[10], stage4_41[11]},
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], stage4_43[5]},
      {stage5_45[0],stage5_44[2],stage5_43[3],stage5_42[3],stage5_41[4]}
   );
   gpc615_5 gpc5601 (
      {stage4_43[6], stage4_43[7], stage4_43[8], stage4_43[9], stage4_43[10]},
      {stage4_44[0]},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[0],stage5_45[1],stage5_44[3],stage5_43[4]}
   );
   gpc615_5 gpc5602 (
      {stage4_43[11], stage4_43[12], stage4_43[13], stage4_43[14], stage4_43[15]},
      {stage4_44[1]},
      {stage4_45[6], stage4_45[7], stage4_45[8], stage4_45[9], stage4_45[10], stage4_45[11]},
      {stage5_47[1],stage5_46[1],stage5_45[2],stage5_44[4],stage5_43[5]}
   );
   gpc606_5 gpc5603 (
      {stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5], stage4_44[6], stage4_44[7]},
      {stage4_46[0], stage4_46[1], stage4_46[2], stage4_46[3], stage4_46[4], stage4_46[5]},
      {stage5_48[0],stage5_47[2],stage5_46[2],stage5_45[3],stage5_44[5]}
   );
   gpc606_5 gpc5604 (
      {stage4_44[8], stage4_44[9], stage4_44[10], stage4_44[11], stage4_44[12], stage4_44[13]},
      {stage4_46[6], stage4_46[7], stage4_46[8], stage4_46[9], stage4_46[10], stage4_46[11]},
      {stage5_48[1],stage5_47[3],stage5_46[3],stage5_45[4],stage5_44[6]}
   );
   gpc615_5 gpc5605 (
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4]},
      {stage4_48[0]},
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4], stage4_49[5]},
      {stage5_51[0],stage5_50[0],stage5_49[0],stage5_48[2],stage5_47[4]}
   );
   gpc615_5 gpc5606 (
      {stage4_47[5], stage4_47[6], stage4_47[7], stage4_47[8], stage4_47[9]},
      {stage4_48[1]},
      {stage4_49[6], stage4_49[7], stage4_49[8], stage4_49[9], stage4_49[10], stage4_49[11]},
      {stage5_51[1],stage5_50[1],stage5_49[1],stage5_48[3],stage5_47[5]}
   );
   gpc615_5 gpc5607 (
      {stage4_47[10], stage4_47[11], stage4_47[12], stage4_47[13], stage4_47[14]},
      {stage4_48[2]},
      {stage4_49[12], stage4_49[13], stage4_49[14], stage4_49[15], stage4_49[16], stage4_49[17]},
      {stage5_51[2],stage5_50[2],stage5_49[2],stage5_48[4],stage5_47[6]}
   );
   gpc606_5 gpc5608 (
      {stage4_48[3], stage4_48[4], stage4_48[5], stage4_48[6], stage4_48[7], stage4_48[8]},
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5]},
      {stage5_52[0],stage5_51[3],stage5_50[3],stage5_49[3],stage5_48[5]}
   );
   gpc606_5 gpc5609 (
      {stage4_48[9], stage4_48[10], stage4_48[11], stage4_48[12], stage4_48[13], stage4_48[14]},
      {stage4_50[6], stage4_50[7], stage4_50[8], stage4_50[9], stage4_50[10], stage4_50[11]},
      {stage5_52[1],stage5_51[4],stage5_50[4],stage5_49[4],stage5_48[6]}
   );
   gpc606_5 gpc5610 (
      {stage4_49[18], stage4_49[19], stage4_49[20], stage4_49[21], stage4_49[22], stage4_49[23]},
      {stage4_51[0], stage4_51[1], stage4_51[2], stage4_51[3], stage4_51[4], stage4_51[5]},
      {stage5_53[0],stage5_52[2],stage5_51[5],stage5_50[5],stage5_49[5]}
   );
   gpc606_5 gpc5611 (
      {stage4_49[24], stage4_49[25], stage4_49[26], stage4_49[27], stage4_49[28], stage4_49[29]},
      {stage4_51[6], stage4_51[7], stage4_51[8], stage4_51[9], stage4_51[10], stage4_51[11]},
      {stage5_53[1],stage5_52[3],stage5_51[6],stage5_50[6],stage5_49[6]}
   );
   gpc606_5 gpc5612 (
      {stage4_49[30], stage4_49[31], stage4_49[32], stage4_49[33], stage4_49[34], stage4_49[35]},
      {stage4_51[12], stage4_51[13], stage4_51[14], stage4_51[15], stage4_51[16], stage4_51[17]},
      {stage5_53[2],stage5_52[4],stage5_51[7],stage5_50[7],stage5_49[7]}
   );
   gpc615_5 gpc5613 (
      {stage4_50[12], stage4_50[13], stage4_50[14], stage4_50[15], stage4_50[16]},
      {stage4_51[18]},
      {stage4_52[0], stage4_52[1], stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5]},
      {stage5_54[0],stage5_53[3],stage5_52[5],stage5_51[8],stage5_50[8]}
   );
   gpc7_3 gpc5614 (
      {stage4_52[6], stage4_52[7], stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11], stage4_52[12]},
      {stage5_54[1],stage5_53[4],stage5_52[6]}
   );
   gpc606_5 gpc5615 (
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], stage4_55[4], stage4_55[5]},
      {stage5_57[0],stage5_56[0],stage5_55[0],stage5_54[2],stage5_53[5]}
   );
   gpc207_4 gpc5616 (
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5], stage4_54[6]},
      {stage4_56[0], stage4_56[1]},
      {stage5_57[1],stage5_56[1],stage5_55[1],stage5_54[3]}
   );
   gpc207_4 gpc5617 (
      {stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10], stage4_54[11], stage4_54[12], stage4_54[13]},
      {stage4_56[2], stage4_56[3]},
      {stage5_57[2],stage5_56[2],stage5_55[2],stage5_54[4]}
   );
   gpc207_4 gpc5618 (
      {stage4_54[14], stage4_54[15], stage4_54[16], stage4_54[17], 1'b0, 1'b0, 1'b0},
      {stage4_56[4], stage4_56[5]},
      {stage5_57[3],stage5_56[3],stage5_55[3],stage5_54[5]}
   );
   gpc606_5 gpc5619 (
      {stage4_55[6], stage4_55[7], stage4_55[8], stage4_55[9], stage4_55[10], stage4_55[11]},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3], stage4_57[4], stage4_57[5]},
      {stage5_59[0],stage5_58[0],stage5_57[4],stage5_56[4],stage5_55[4]}
   );
   gpc606_5 gpc5620 (
      {stage4_56[6], stage4_56[7], stage4_56[8], stage4_56[9], stage4_56[10], stage4_56[11]},
      {stage4_58[0], stage4_58[1], stage4_58[2], stage4_58[3], stage4_58[4], stage4_58[5]},
      {stage5_60[0],stage5_59[1],stage5_58[1],stage5_57[5],stage5_56[5]}
   );
   gpc7_3 gpc5621 (
      {stage4_57[6], stage4_57[7], stage4_57[8], stage4_57[9], stage4_57[10], stage4_57[11], 1'b0},
      {stage5_59[2],stage5_58[2],stage5_57[6]}
   );
   gpc7_3 gpc5622 (
      {stage4_58[6], stage4_58[7], stage4_58[8], stage4_58[9], stage4_58[10], stage4_58[11], stage4_58[12]},
      {stage5_60[1],stage5_59[3],stage5_58[3]}
   );
   gpc7_3 gpc5623 (
      {stage4_58[13], stage4_58[14], stage4_58[15], stage4_58[16], stage4_58[17], stage4_58[18], stage4_58[19]},
      {stage5_60[2],stage5_59[4],stage5_58[4]}
   );
   gpc606_5 gpc5624 (
      {stage4_59[0], stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[0],stage5_61[0],stage5_60[3],stage5_59[5]}
   );
   gpc606_5 gpc5625 (
      {stage4_59[6], stage4_59[7], stage4_59[8], stage4_59[9], stage4_59[10], stage4_59[11]},
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], stage4_61[10], stage4_61[11]},
      {stage5_63[1],stage5_62[1],stage5_61[1],stage5_60[4],stage5_59[6]}
   );
   gpc606_5 gpc5626 (
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[2],stage5_62[2],stage5_61[2],stage5_60[5]}
   );
   gpc606_5 gpc5627 (
      {stage4_60[6], stage4_60[7], stage4_60[8], stage4_60[9], stage4_60[10], stage4_60[11]},
      {stage4_62[6], stage4_62[7], stage4_62[8], stage4_62[9], stage4_62[10], stage4_62[11]},
      {stage5_64[1],stage5_63[3],stage5_62[3],stage5_61[3],stage5_60[6]}
   );
   gpc117_4 gpc5628 (
      {stage4_63[0], stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5], stage4_63[6]},
      {stage4_64[0]},
      {stage4_65[0]},
      {stage5_66[0],stage5_65[0],stage5_64[2],stage5_63[4]}
   );
   gpc117_4 gpc5629 (
      {stage4_63[7], stage4_63[8], stage4_63[9], stage4_63[10], stage4_63[11], stage4_63[12], 1'b0},
      {stage4_64[1]},
      {stage4_65[1]},
      {stage5_66[1],stage5_65[1],stage5_64[3],stage5_63[5]}
   );
   gpc606_5 gpc5630 (
      {stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6], stage4_64[7]},
      {stage4_66[0], stage4_66[1], stage4_66[2], stage4_66[3], stage4_66[4], stage4_66[5]},
      {stage5_68[0],stage5_67[0],stage5_66[2],stage5_65[2],stage5_64[4]}
   );
   gpc606_5 gpc5631 (
      {stage4_64[8], stage4_64[9], stage4_64[10], stage4_64[11], 1'b0, 1'b0},
      {stage4_66[6], stage4_66[7], stage4_66[8], stage4_66[9], stage4_66[10], stage4_66[11]},
      {stage5_68[1],stage5_67[1],stage5_66[3],stage5_65[3],stage5_64[5]}
   );
   gpc606_5 gpc5632 (
      {stage4_65[2], stage4_65[3], stage4_65[4], stage4_65[5], stage4_65[6], stage4_65[7]},
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], stage4_67[4], stage4_67[5]},
      {stage5_69[0],stage5_68[2],stage5_67[2],stage5_66[4],stage5_65[4]}
   );
   gpc207_4 gpc5633 (
      {stage4_66[12], stage4_66[13], stage4_66[14], stage4_66[15], stage4_66[16], stage4_66[17], stage4_66[18]},
      {stage4_68[0], stage4_68[1]},
      {stage5_69[1],stage5_68[3],stage5_67[3],stage5_66[5]}
   );
   gpc1_1 gpc5634 (
      {stage4_0[11]},
      {stage5_0[2]}
   );
   gpc1_1 gpc5635 (
      {stage4_0[12]},
      {stage5_0[3]}
   );
   gpc1_1 gpc5636 (
      {stage4_0[13]},
      {stage5_0[4]}
   );
   gpc1_1 gpc5637 (
      {stage4_1[3]},
      {stage5_1[2]}
   );
   gpc1_1 gpc5638 (
      {stage4_1[4]},
      {stage5_1[3]}
   );
   gpc1_1 gpc5639 (
      {stage4_3[17]},
      {stage5_3[5]}
   );
   gpc1_1 gpc5640 (
      {stage4_3[18]},
      {stage5_3[6]}
   );
   gpc1_1 gpc5641 (
      {stage4_4[5]},
      {stage5_4[5]}
   );
   gpc1_1 gpc5642 (
      {stage4_4[6]},
      {stage5_4[6]}
   );
   gpc1_1 gpc5643 (
      {stage4_4[7]},
      {stage5_4[7]}
   );
   gpc1_1 gpc5644 (
      {stage4_4[8]},
      {stage5_4[8]}
   );
   gpc1_1 gpc5645 (
      {stage4_4[9]},
      {stage5_4[9]}
   );
   gpc1_1 gpc5646 (
      {stage4_5[16]},
      {stage5_5[4]}
   );
   gpc1_1 gpc5647 (
      {stage4_5[17]},
      {stage5_5[5]}
   );
   gpc1_1 gpc5648 (
      {stage4_5[18]},
      {stage5_5[6]}
   );
   gpc1_1 gpc5649 (
      {stage4_5[19]},
      {stage5_5[7]}
   );
   gpc1_1 gpc5650 (
      {stage4_6[8]},
      {stage5_6[4]}
   );
   gpc1_1 gpc5651 (
      {stage4_6[9]},
      {stage5_6[5]}
   );
   gpc1_1 gpc5652 (
      {stage4_7[8]},
      {stage5_7[5]}
   );
   gpc1_1 gpc5653 (
      {stage4_7[9]},
      {stage5_7[6]}
   );
   gpc1_1 gpc5654 (
      {stage4_9[3]},
      {stage5_9[5]}
   );
   gpc1_1 gpc5655 (
      {stage4_9[4]},
      {stage5_9[6]}
   );
   gpc1_1 gpc5656 (
      {stage4_9[5]},
      {stage5_9[7]}
   );
   gpc1_1 gpc5657 (
      {stage4_9[6]},
      {stage5_9[8]}
   );
   gpc1_1 gpc5658 (
      {stage4_9[7]},
      {stage5_9[9]}
   );
   gpc1_1 gpc5659 (
      {stage4_10[13]},
      {stage5_10[5]}
   );
   gpc1_1 gpc5660 (
      {stage4_11[7]},
      {stage5_11[5]}
   );
   gpc1_1 gpc5661 (
      {stage4_11[8]},
      {stage5_11[6]}
   );
   gpc1_1 gpc5662 (
      {stage4_11[9]},
      {stage5_11[7]}
   );
   gpc1_1 gpc5663 (
      {stage4_11[10]},
      {stage5_11[8]}
   );
   gpc1_1 gpc5664 (
      {stage4_11[11]},
      {stage5_11[9]}
   );
   gpc1_1 gpc5665 (
      {stage4_12[17]},
      {stage5_12[5]}
   );
   gpc1_1 gpc5666 (
      {stage4_13[13]},
      {stage5_13[5]}
   );
   gpc1_1 gpc5667 (
      {stage4_15[11]},
      {stage5_15[5]}
   );
   gpc1_1 gpc5668 (
      {stage4_17[12]},
      {stage5_17[5]}
   );
   gpc1_1 gpc5669 (
      {stage4_17[13]},
      {stage5_17[6]}
   );
   gpc1_1 gpc5670 (
      {stage4_17[14]},
      {stage5_17[7]}
   );
   gpc1_1 gpc5671 (
      {stage4_19[9]},
      {stage5_19[6]}
   );
   gpc1_1 gpc5672 (
      {stage4_19[10]},
      {stage5_19[7]}
   );
   gpc1_1 gpc5673 (
      {stage4_19[11]},
      {stage5_19[8]}
   );
   gpc1_1 gpc5674 (
      {stage4_19[12]},
      {stage5_19[9]}
   );
   gpc1_1 gpc5675 (
      {stage4_19[13]},
      {stage5_19[10]}
   );
   gpc1_1 gpc5676 (
      {stage4_21[0]},
      {stage5_21[3]}
   );
   gpc1_1 gpc5677 (
      {stage4_21[1]},
      {stage5_21[4]}
   );
   gpc1_1 gpc5678 (
      {stage4_21[2]},
      {stage5_21[5]}
   );
   gpc1_1 gpc5679 (
      {stage4_21[3]},
      {stage5_21[6]}
   );
   gpc1_1 gpc5680 (
      {stage4_21[4]},
      {stage5_21[7]}
   );
   gpc1_1 gpc5681 (
      {stage4_21[5]},
      {stage5_21[8]}
   );
   gpc1_1 gpc5682 (
      {stage4_21[6]},
      {stage5_21[9]}
   );
   gpc1_1 gpc5683 (
      {stage4_21[7]},
      {stage5_21[10]}
   );
   gpc1_1 gpc5684 (
      {stage4_21[8]},
      {stage5_21[11]}
   );
   gpc1_1 gpc5685 (
      {stage4_24[9]},
      {stage5_24[4]}
   );
   gpc1_1 gpc5686 (
      {stage4_24[10]},
      {stage5_24[5]}
   );
   gpc1_1 gpc5687 (
      {stage4_24[11]},
      {stage5_24[6]}
   );
   gpc1_1 gpc5688 (
      {stage4_29[13]},
      {stage5_29[4]}
   );
   gpc1_1 gpc5689 (
      {stage4_29[14]},
      {stage5_29[5]}
   );
   gpc1_1 gpc5690 (
      {stage4_29[15]},
      {stage5_29[6]}
   );
   gpc1_1 gpc5691 (
      {stage4_29[16]},
      {stage5_29[7]}
   );
   gpc1_1 gpc5692 (
      {stage4_31[8]},
      {stage5_31[5]}
   );
   gpc1_1 gpc5693 (
      {stage4_31[9]},
      {stage5_31[6]}
   );
   gpc1_1 gpc5694 (
      {stage4_36[12]},
      {stage5_36[6]}
   );
   gpc1_1 gpc5695 (
      {stage4_37[6]},
      {stage5_37[6]}
   );
   gpc1_1 gpc5696 (
      {stage4_37[7]},
      {stage5_37[7]}
   );
   gpc1_1 gpc5697 (
      {stage4_37[8]},
      {stage5_37[8]}
   );
   gpc1_1 gpc5698 (
      {stage4_37[9]},
      {stage5_37[9]}
   );
   gpc1_1 gpc5699 (
      {stage4_37[10]},
      {stage5_37[10]}
   );
   gpc1_1 gpc5700 (
      {stage4_37[11]},
      {stage5_37[11]}
   );
   gpc1_1 gpc5701 (
      {stage4_38[6]},
      {stage5_38[3]}
   );
   gpc1_1 gpc5702 (
      {stage4_40[12]},
      {stage5_40[5]}
   );
   gpc1_1 gpc5703 (
      {stage4_42[12]},
      {stage5_42[4]}
   );
   gpc1_1 gpc5704 (
      {stage4_42[13]},
      {stage5_42[5]}
   );
   gpc1_1 gpc5705 (
      {stage4_42[14]},
      {stage5_42[6]}
   );
   gpc1_1 gpc5706 (
      {stage4_43[16]},
      {stage5_43[6]}
   );
   gpc1_1 gpc5707 (
      {stage4_43[17]},
      {stage5_43[7]}
   );
   gpc1_1 gpc5708 (
      {stage4_43[18]},
      {stage5_43[8]}
   );
   gpc1_1 gpc5709 (
      {stage4_43[19]},
      {stage5_43[9]}
   );
   gpc1_1 gpc5710 (
      {stage4_46[12]},
      {stage5_46[4]}
   );
   gpc1_1 gpc5711 (
      {stage4_46[13]},
      {stage5_46[5]}
   );
   gpc1_1 gpc5712 (
      {stage4_46[14]},
      {stage5_46[6]}
   );
   gpc1_1 gpc5713 (
      {stage4_51[19]},
      {stage5_51[9]}
   );
   gpc1_1 gpc5714 (
      {stage4_52[13]},
      {stage5_52[7]}
   );
   gpc1_1 gpc5715 (
      {stage4_53[6]},
      {stage5_53[6]}
   );
   gpc1_1 gpc5716 (
      {stage4_53[7]},
      {stage5_53[7]}
   );
   gpc1_1 gpc5717 (
      {stage4_53[8]},
      {stage5_53[8]}
   );
   gpc1_1 gpc5718 (
      {stage4_53[9]},
      {stage5_53[9]}
   );
   gpc1_1 gpc5719 (
      {stage4_53[10]},
      {stage5_53[10]}
   );
   gpc1_1 gpc5720 (
      {stage4_53[11]},
      {stage5_53[11]}
   );
   gpc1_1 gpc5721 (
      {stage4_53[12]},
      {stage5_53[12]}
   );
   gpc1_1 gpc5722 (
      {stage4_53[13]},
      {stage5_53[13]}
   );
   gpc1_1 gpc5723 (
      {stage4_53[14]},
      {stage5_53[14]}
   );
   gpc1_1 gpc5724 (
      {stage4_55[12]},
      {stage5_55[5]}
   );
   gpc1_1 gpc5725 (
      {stage4_60[12]},
      {stage5_60[7]}
   );
   gpc1_1 gpc5726 (
      {stage4_60[13]},
      {stage5_60[8]}
   );
   gpc1_1 gpc5727 (
      {stage4_66[19]},
      {stage5_66[6]}
   );
   gpc1_1 gpc5728 (
      {stage4_66[20]},
      {stage5_66[7]}
   );
   gpc1_1 gpc5729 (
      {stage4_66[21]},
      {stage5_66[8]}
   );
   gpc1_1 gpc5730 (
      {stage4_66[22]},
      {stage5_66[9]}
   );
   gpc1_1 gpc5731 (
      {stage4_66[23]},
      {stage5_66[10]}
   );
   gpc1_1 gpc5732 (
      {stage4_67[6]},
      {stage5_67[4]}
   );
   gpc1_1 gpc5733 (
      {stage4_67[7]},
      {stage5_67[5]}
   );
   gpc1_1 gpc5734 (
      {stage4_67[8]},
      {stage5_67[6]}
   );
   gpc1_1 gpc5735 (
      {stage4_68[2]},
      {stage5_68[4]}
   );
   gpc1_1 gpc5736 (
      {stage4_69[0]},
      {stage5_69[2]}
   );
   gpc223_4 gpc5737 (
      {stage5_2[0], stage5_2[1], 1'b0},
      {stage5_3[0], stage5_3[1]},
      {stage5_4[0], stage5_4[1]},
      {stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc615_5 gpc5738 (
      {stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5], stage5_3[6]},
      {stage5_4[2]},
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5]},
      {stage6_7[0],stage6_6[0],stage6_5[1],stage6_4[1],stage6_3[1]}
   );
   gpc615_5 gpc5739 (
      {stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_5[6]},
      {stage5_6[0], stage5_6[1], stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5]},
      {stage6_8[0],stage6_7[1],stage6_6[1],stage6_5[2],stage6_4[2]}
   );
   gpc207_4 gpc5740 (
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3], stage5_7[4], stage5_7[5], stage5_7[6]},
      {stage5_9[0], stage5_9[1]},
      {stage6_10[0],stage6_9[0],stage6_8[1],stage6_7[2]}
   );
   gpc615_5 gpc5741 (
      {stage5_8[0], stage5_8[1], stage5_8[2], stage5_8[3], stage5_8[4]},
      {stage5_9[2]},
      {stage5_10[0], stage5_10[1], stage5_10[2], stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[1],stage6_8[2]}
   );
   gpc606_5 gpc5742 (
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc7_3 gpc5743 (
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], 1'b0},
      {stage6_14[1],stage6_13[1],stage6_12[2]}
   );
   gpc615_5 gpc5744 (
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4]},
      {stage5_16[0]},
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage6_19[0],stage6_18[0],stage6_17[0],stage6_16[0],stage6_15[1]}
   );
   gpc1415_5 gpc5745 (
      {stage5_16[1], stage5_16[2], stage5_16[3], stage5_16[4], stage5_16[5]},
      {stage5_17[6]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3]},
      {stage5_19[0]},
      {stage6_20[0],stage6_19[1],stage6_18[1],stage6_17[1],stage6_16[1]}
   );
   gpc615_5 gpc5746 (
      {stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage5_20[0]},
      {stage5_21[0], stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[1],stage6_19[2]}
   );
   gpc615_5 gpc5747 (
      {stage5_19[6], stage5_19[7], stage5_19[8], stage5_19[9], stage5_19[10]},
      {stage5_20[1]},
      {stage5_21[6], stage5_21[7], stage5_21[8], stage5_21[9], stage5_21[10], stage5_21[11]},
      {stage6_23[1],stage6_22[1],stage6_21[1],stage6_20[2],stage6_19[3]}
   );
   gpc615_5 gpc5748 (
      {stage5_22[0], stage5_22[1], stage5_22[2], stage5_22[3], stage5_22[4]},
      {stage5_23[0]},
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5]},
      {stage6_26[0],stage6_25[0],stage6_24[0],stage6_23[2],stage6_22[2]}
   );
   gpc207_4 gpc5749 (
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3], stage5_26[4], stage5_26[5], 1'b0},
      {stage5_28[0], stage5_28[1]},
      {stage6_29[0],stage6_28[0],stage6_27[0],stage6_26[1]}
   );
   gpc1325_5 gpc5750 (
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3], stage5_27[4]},
      {stage5_28[2], stage5_28[3]},
      {stage5_29[0], stage5_29[1], stage5_29[2]},
      {stage5_30[0]},
      {stage6_31[0],stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[1]}
   );
   gpc615_5 gpc5751 (
      {stage5_29[3], stage5_29[4], stage5_29[5], stage5_29[6], stage5_29[7]},
      {stage5_30[1]},
      {stage5_31[0], stage5_31[1], stage5_31[2], stage5_31[3], stage5_31[4], stage5_31[5]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[1],stage6_29[2]}
   );
   gpc2135_5 gpc5752 (
      {stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], 1'b0},
      {stage5_31[6], 1'b0, 1'b0},
      {stage5_32[0]},
      {stage5_33[0], stage5_33[1]},
      {stage6_34[0],stage6_33[1],stage6_32[1],stage6_31[2],stage6_30[2]}
   );
   gpc615_5 gpc5753 (
      {stage5_32[1], stage5_32[2], stage5_32[3], 1'b0, 1'b0},
      {stage5_33[2]},
      {stage5_34[0], stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5]},
      {stage6_36[0],stage6_35[0],stage6_34[1],stage6_33[2],stage6_32[2]}
   );
   gpc117_4 gpc5754 (
      {stage5_33[3], stage5_33[4], stage5_33[5], stage5_33[6], 1'b0, 1'b0, 1'b0},
      {stage5_34[6]},
      {stage5_35[0]},
      {stage6_36[1],stage6_35[1],stage6_34[2],stage6_33[3]}
   );
   gpc623_5 gpc5755 (
      {stage5_35[1], stage5_35[2], stage5_35[3]},
      {stage5_36[0], stage5_36[1]},
      {stage5_37[0], stage5_37[1], stage5_37[2], stage5_37[3], stage5_37[4], stage5_37[5]},
      {stage6_39[0],stage6_38[0],stage6_37[0],stage6_36[2],stage6_35[2]}
   );
   gpc606_5 gpc5756 (
      {stage5_36[2], stage5_36[3], stage5_36[4], stage5_36[5], stage5_36[6], 1'b0},
      {stage5_38[0], stage5_38[1], stage5_38[2], stage5_38[3], 1'b0, 1'b0},
      {stage6_40[0],stage6_39[1],stage6_38[1],stage6_37[1],stage6_36[3]}
   );
   gpc1163_5 gpc5757 (
      {stage5_39[0], stage5_39[1], stage5_39[2]},
      {stage5_40[0], stage5_40[1], stage5_40[2], stage5_40[3], stage5_40[4], stage5_40[5]},
      {stage5_41[0]},
      {stage5_42[0]},
      {stage6_43[0],stage6_42[0],stage6_41[0],stage6_40[1],stage6_39[2]}
   );
   gpc1415_5 gpc5758 (
      {stage5_41[1], stage5_41[2], stage5_41[3], stage5_41[4], 1'b0},
      {stage5_42[1]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3]},
      {stage5_44[0]},
      {stage6_45[0],stage6_44[0],stage6_43[1],stage6_42[1],stage6_41[1]}
   );
   gpc135_4 gpc5759 (
      {stage5_42[2], stage5_42[3], stage5_42[4], stage5_42[5], stage5_42[6]},
      {stage5_43[4], stage5_43[5], stage5_43[6]},
      {stage5_44[1]},
      {stage6_45[1],stage6_44[1],stage6_43[2],stage6_42[2]}
   );
   gpc606_5 gpc5760 (
      {stage5_44[2], stage5_44[3], stage5_44[4], stage5_44[5], stage5_44[6], 1'b0},
      {stage5_46[0], stage5_46[1], stage5_46[2], stage5_46[3], stage5_46[4], stage5_46[5]},
      {stage6_48[0],stage6_47[0],stage6_46[0],stage6_45[2],stage6_44[2]}
   );
   gpc2135_5 gpc5761 (
      {stage5_45[0], stage5_45[1], stage5_45[2], stage5_45[3], stage5_45[4]},
      {stage5_46[6], 1'b0, 1'b0},
      {stage5_47[0]},
      {stage5_48[0], stage5_48[1]},
      {stage6_49[0],stage6_48[1],stage6_47[1],stage6_46[1],stage6_45[3]}
   );
   gpc623_5 gpc5762 (
      {stage5_47[1], stage5_47[2], stage5_47[3]},
      {stage5_48[2], stage5_48[3]},
      {stage5_49[0], stage5_49[1], stage5_49[2], stage5_49[3], stage5_49[4], stage5_49[5]},
      {stage6_51[0],stage6_50[0],stage6_49[1],stage6_48[2],stage6_47[2]}
   );
   gpc223_4 gpc5763 (
      {stage5_48[4], stage5_48[5], stage5_48[6]},
      {stage5_49[6], stage5_49[7]},
      {stage5_50[0], stage5_50[1]},
      {stage6_51[1],stage6_50[1],stage6_49[2],stage6_48[3]}
   );
   gpc606_5 gpc5764 (
      {stage5_50[2], stage5_50[3], stage5_50[4], stage5_50[5], stage5_50[6], stage5_50[7]},
      {stage5_52[0], stage5_52[1], stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5]},
      {stage6_54[0],stage6_53[0],stage6_52[0],stage6_51[2],stage6_50[2]}
   );
   gpc615_5 gpc5765 (
      {stage5_51[0], stage5_51[1], stage5_51[2], stage5_51[3], stage5_51[4]},
      {stage5_52[6]},
      {stage5_53[0], stage5_53[1], stage5_53[2], stage5_53[3], stage5_53[4], stage5_53[5]},
      {stage6_55[0],stage6_54[1],stage6_53[1],stage6_52[1],stage6_51[3]}
   );
   gpc615_5 gpc5766 (
      {stage5_51[5], stage5_51[6], stage5_51[7], stage5_51[8], stage5_51[9]},
      {stage5_52[7]},
      {stage5_53[6], stage5_53[7], stage5_53[8], stage5_53[9], stage5_53[10], stage5_53[11]},
      {stage6_55[1],stage6_54[2],stage6_53[2],stage6_52[2],stage6_51[4]}
   );
   gpc1163_5 gpc5767 (
      {stage5_53[12], stage5_53[13], stage5_53[14]},
      {stage5_54[0], stage5_54[1], stage5_54[2], stage5_54[3], stage5_54[4], stage5_54[5]},
      {stage5_55[0]},
      {stage5_56[0]},
      {stage6_57[0],stage6_56[0],stage6_55[2],stage6_54[3],stage6_53[3]}
   );
   gpc615_5 gpc5768 (
      {stage5_55[1], stage5_55[2], stage5_55[3], stage5_55[4], stage5_55[5]},
      {stage5_56[1]},
      {stage5_57[0], stage5_57[1], stage5_57[2], stage5_57[3], stage5_57[4], stage5_57[5]},
      {stage6_59[0],stage6_58[0],stage6_57[1],stage6_56[1],stage6_55[3]}
   );
   gpc615_5 gpc5769 (
      {stage5_58[0], stage5_58[1], stage5_58[2], stage5_58[3], stage5_58[4]},
      {stage5_59[0]},
      {stage5_60[0], stage5_60[1], stage5_60[2], stage5_60[3], stage5_60[4], stage5_60[5]},
      {stage6_62[0],stage6_61[0],stage6_60[0],stage6_59[1],stage6_58[1]}
   );
   gpc3_2 gpc5770 (
      {stage5_59[1], stage5_59[2], stage5_59[3]},
      {stage6_60[1],stage6_59[2]}
   );
   gpc606_5 gpc5771 (
      {stage5_63[0], stage5_63[1], stage5_63[2], stage5_63[3], stage5_63[4], stage5_63[5]},
      {stage5_65[0], stage5_65[1], stage5_65[2], stage5_65[3], stage5_65[4], 1'b0},
      {stage6_67[0],stage6_66[0],stage6_65[0],stage6_64[0],stage6_63[0]}
   );
   gpc606_5 gpc5772 (
      {stage5_64[0], stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage5_66[0], stage5_66[1], stage5_66[2], stage5_66[3], stage5_66[4], stage5_66[5]},
      {stage6_68[0],stage6_67[1],stage6_66[1],stage6_65[1],stage6_64[1]}
   );
   gpc606_5 gpc5773 (
      {stage5_66[6], stage5_66[7], stage5_66[8], stage5_66[9], stage5_66[10], 1'b0},
      {stage5_68[0], stage5_68[1], stage5_68[2], stage5_68[3], stage5_68[4], 1'b0},
      {stage6_70[0],stage6_69[0],stage6_68[1],stage6_67[2],stage6_66[2]}
   );
   gpc606_5 gpc5774 (
      {stage5_67[0], stage5_67[1], stage5_67[2], stage5_67[3], stage5_67[4], stage5_67[5]},
      {stage5_69[0], stage5_69[1], stage5_69[2], 1'b0, 1'b0, 1'b0},
      {stage6_71[0],stage6_70[1],stage6_69[1],stage6_68[2],stage6_67[3]}
   );
   gpc1_1 gpc5775 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc5776 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc5777 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc5778 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc5779 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc5780 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc5781 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc5782 (
      {stage5_1[2]},
      {stage6_1[2]}
   );
   gpc1_1 gpc5783 (
      {stage5_1[3]},
      {stage6_1[3]}
   );
   gpc1_1 gpc5784 (
      {stage5_4[8]},
      {stage6_4[3]}
   );
   gpc1_1 gpc5785 (
      {stage5_4[9]},
      {stage6_4[4]}
   );
   gpc1_1 gpc5786 (
      {stage5_5[7]},
      {stage6_5[3]}
   );
   gpc1_1 gpc5787 (
      {stage5_9[3]},
      {stage6_9[2]}
   );
   gpc1_1 gpc5788 (
      {stage5_9[4]},
      {stage6_9[3]}
   );
   gpc1_1 gpc5789 (
      {stage5_9[5]},
      {stage6_9[4]}
   );
   gpc1_1 gpc5790 (
      {stage5_9[6]},
      {stage6_9[5]}
   );
   gpc1_1 gpc5791 (
      {stage5_9[7]},
      {stage6_9[6]}
   );
   gpc1_1 gpc5792 (
      {stage5_9[8]},
      {stage6_9[7]}
   );
   gpc1_1 gpc5793 (
      {stage5_9[9]},
      {stage6_9[8]}
   );
   gpc1_1 gpc5794 (
      {stage5_11[6]},
      {stage6_11[2]}
   );
   gpc1_1 gpc5795 (
      {stage5_11[7]},
      {stage6_11[3]}
   );
   gpc1_1 gpc5796 (
      {stage5_11[8]},
      {stage6_11[4]}
   );
   gpc1_1 gpc5797 (
      {stage5_11[9]},
      {stage6_11[5]}
   );
   gpc1_1 gpc5798 (
      {stage5_14[0]},
      {stage6_14[2]}
   );
   gpc1_1 gpc5799 (
      {stage5_14[1]},
      {stage6_14[3]}
   );
   gpc1_1 gpc5800 (
      {stage5_14[2]},
      {stage6_14[4]}
   );
   gpc1_1 gpc5801 (
      {stage5_14[3]},
      {stage6_14[5]}
   );
   gpc1_1 gpc5802 (
      {stage5_14[4]},
      {stage6_14[6]}
   );
   gpc1_1 gpc5803 (
      {stage5_15[5]},
      {stage6_15[2]}
   );
   gpc1_1 gpc5804 (
      {stage5_17[7]},
      {stage6_17[2]}
   );
   gpc1_1 gpc5805 (
      {stage5_18[4]},
      {stage6_18[2]}
   );
   gpc1_1 gpc5806 (
      {stage5_18[5]},
      {stage6_18[3]}
   );
   gpc1_1 gpc5807 (
      {stage5_20[2]},
      {stage6_20[3]}
   );
   gpc1_1 gpc5808 (
      {stage5_23[1]},
      {stage6_23[3]}
   );
   gpc1_1 gpc5809 (
      {stage5_23[2]},
      {stage6_23[4]}
   );
   gpc1_1 gpc5810 (
      {stage5_24[6]},
      {stage6_24[1]}
   );
   gpc1_1 gpc5811 (
      {stage5_25[0]},
      {stage6_25[1]}
   );
   gpc1_1 gpc5812 (
      {stage5_25[1]},
      {stage6_25[2]}
   );
   gpc1_1 gpc5813 (
      {stage5_25[2]},
      {stage6_25[3]}
   );
   gpc1_1 gpc5814 (
      {stage5_25[3]},
      {stage6_25[4]}
   );
   gpc1_1 gpc5815 (
      {stage5_25[4]},
      {stage6_25[5]}
   );
   gpc1_1 gpc5816 (
      {stage5_25[5]},
      {stage6_25[6]}
   );
   gpc1_1 gpc5817 (
      {stage5_27[5]},
      {stage6_27[2]}
   );
   gpc1_1 gpc5818 (
      {stage5_35[4]},
      {stage6_35[3]}
   );
   gpc1_1 gpc5819 (
      {stage5_37[6]},
      {stage6_37[2]}
   );
   gpc1_1 gpc5820 (
      {stage5_37[7]},
      {stage6_37[3]}
   );
   gpc1_1 gpc5821 (
      {stage5_37[8]},
      {stage6_37[4]}
   );
   gpc1_1 gpc5822 (
      {stage5_37[9]},
      {stage6_37[5]}
   );
   gpc1_1 gpc5823 (
      {stage5_37[10]},
      {stage6_37[6]}
   );
   gpc1_1 gpc5824 (
      {stage5_37[11]},
      {stage6_37[7]}
   );
   gpc1_1 gpc5825 (
      {stage5_43[7]},
      {stage6_43[3]}
   );
   gpc1_1 gpc5826 (
      {stage5_43[8]},
      {stage6_43[4]}
   );
   gpc1_1 gpc5827 (
      {stage5_43[9]},
      {stage6_43[5]}
   );
   gpc1_1 gpc5828 (
      {stage5_47[4]},
      {stage6_47[3]}
   );
   gpc1_1 gpc5829 (
      {stage5_47[5]},
      {stage6_47[4]}
   );
   gpc1_1 gpc5830 (
      {stage5_47[6]},
      {stage6_47[5]}
   );
   gpc1_1 gpc5831 (
      {stage5_50[8]},
      {stage6_50[3]}
   );
   gpc1_1 gpc5832 (
      {stage5_56[2]},
      {stage6_56[2]}
   );
   gpc1_1 gpc5833 (
      {stage5_56[3]},
      {stage6_56[3]}
   );
   gpc1_1 gpc5834 (
      {stage5_56[4]},
      {stage6_56[4]}
   );
   gpc1_1 gpc5835 (
      {stage5_56[5]},
      {stage6_56[5]}
   );
   gpc1_1 gpc5836 (
      {stage5_57[6]},
      {stage6_57[2]}
   );
   gpc1_1 gpc5837 (
      {stage5_59[4]},
      {stage6_59[3]}
   );
   gpc1_1 gpc5838 (
      {stage5_59[5]},
      {stage6_59[4]}
   );
   gpc1_1 gpc5839 (
      {stage5_59[6]},
      {stage6_59[5]}
   );
   gpc1_1 gpc5840 (
      {stage5_60[6]},
      {stage6_60[2]}
   );
   gpc1_1 gpc5841 (
      {stage5_60[7]},
      {stage6_60[3]}
   );
   gpc1_1 gpc5842 (
      {stage5_60[8]},
      {stage6_60[4]}
   );
   gpc1_1 gpc5843 (
      {stage5_61[0]},
      {stage6_61[1]}
   );
   gpc1_1 gpc5844 (
      {stage5_61[1]},
      {stage6_61[2]}
   );
   gpc1_1 gpc5845 (
      {stage5_61[2]},
      {stage6_61[3]}
   );
   gpc1_1 gpc5846 (
      {stage5_61[3]},
      {stage6_61[4]}
   );
   gpc1_1 gpc5847 (
      {stage5_62[0]},
      {stage6_62[1]}
   );
   gpc1_1 gpc5848 (
      {stage5_62[1]},
      {stage6_62[2]}
   );
   gpc1_1 gpc5849 (
      {stage5_62[2]},
      {stage6_62[3]}
   );
   gpc1_1 gpc5850 (
      {stage5_62[3]},
      {stage6_62[4]}
   );
   gpc1_1 gpc5851 (
      {stage5_67[6]},
      {stage6_67[4]}
   );
   gpc135_4 gpc5852 (
      {stage6_0[0], stage6_0[1], stage6_0[2], stage6_0[3], stage6_0[4]},
      {stage6_1[0], stage6_1[1], stage6_1[2]},
      {stage6_2[0]},
      {stage7_3[0],stage7_2[0],stage7_1[0],stage7_0[0]}
   );
   gpc1343_5 gpc5853 (
      {stage6_3[0], stage6_3[1], 1'b0},
      {stage6_4[0], stage6_4[1], stage6_4[2], stage6_4[3]},
      {stage6_5[0], stage6_5[1], stage6_5[2]},
      {stage6_6[0]},
      {stage7_7[0],stage7_6[0],stage7_5[0],stage7_4[0],stage7_3[1]}
   );
   gpc1423_5 gpc5854 (
      {stage6_7[0], stage6_7[1], stage6_7[2]},
      {stage6_8[0], stage6_8[1]},
      {stage6_9[0], stage6_9[1], stage6_9[2], stage6_9[3]},
      {stage6_10[0]},
      {stage7_11[0],stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[1]}
   );
   gpc615_5 gpc5855 (
      {stage6_9[4], stage6_9[5], stage6_9[6], stage6_9[7], stage6_9[8]},
      {stage6_10[1]},
      {stage6_11[0], stage6_11[1], stage6_11[2], stage6_11[3], stage6_11[4], stage6_11[5]},
      {stage7_13[0],stage7_12[0],stage7_11[1],stage7_10[1],stage7_9[1]}
   );
   gpc623_5 gpc5856 (
      {stage6_12[0], stage6_12[1], stage6_12[2]},
      {stage6_13[0], stage6_13[1]},
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5]},
      {stage7_16[0],stage7_15[0],stage7_14[0],stage7_13[1],stage7_12[1]}
   );
   gpc2223_5 gpc5857 (
      {stage6_15[0], stage6_15[1], stage6_15[2]},
      {stage6_16[0], stage6_16[1]},
      {stage6_17[0], stage6_17[1]},
      {stage6_18[0], stage6_18[1]},
      {stage7_19[0],stage7_18[0],stage7_17[0],stage7_16[1],stage7_15[1]}
   );
   gpc1343_5 gpc5858 (
      {stage6_18[2], stage6_18[3], 1'b0},
      {stage6_19[0], stage6_19[1], stage6_19[2], stage6_19[3]},
      {stage6_20[0], stage6_20[1], stage6_20[2]},
      {stage6_21[0]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[1],stage7_18[1]}
   );
   gpc3_2 gpc5859 (
      {stage6_22[0], stage6_22[1], stage6_22[2]},
      {stage7_23[0],stage7_22[1]}
   );
   gpc1415_5 gpc5860 (
      {stage6_23[0], stage6_23[1], stage6_23[2], stage6_23[3], stage6_23[4]},
      {stage6_24[0]},
      {stage6_25[0], stage6_25[1], stage6_25[2], stage6_25[3]},
      {stage6_26[0]},
      {stage7_27[0],stage7_26[0],stage7_25[0],stage7_24[0],stage7_23[1]}
   );
   gpc1343_5 gpc5861 (
      {stage6_25[4], stage6_25[5], stage6_25[6]},
      {stage6_26[1], 1'b0, 1'b0, 1'b0},
      {stage6_27[0], stage6_27[1], stage6_27[2]},
      {stage6_28[0]},
      {stage7_29[0],stage7_28[0],stage7_27[1],stage7_26[1],stage7_25[1]}
   );
   gpc1423_5 gpc5862 (
      {stage6_29[0], stage6_29[1], stage6_29[2]},
      {stage6_30[0], stage6_30[1]},
      {stage6_31[0], stage6_31[1], stage6_31[2], 1'b0},
      {stage6_32[0]},
      {stage7_33[0],stage7_32[0],stage7_31[0],stage7_30[0],stage7_29[1]}
   );
   gpc1343_5 gpc5863 (
      {stage6_32[1], stage6_32[2], 1'b0},
      {stage6_33[0], stage6_33[1], stage6_33[2], stage6_33[3]},
      {stage6_34[0], stage6_34[1], stage6_34[2]},
      {stage6_35[0]},
      {stage7_36[0],stage7_35[0],stage7_34[0],stage7_33[1],stage7_32[1]}
   );
   gpc1343_5 gpc5864 (
      {stage6_35[1], stage6_35[2], stage6_35[3]},
      {stage6_36[0], stage6_36[1], stage6_36[2], stage6_36[3]},
      {stage6_37[0], stage6_37[1], stage6_37[2]},
      {stage6_38[0]},
      {stage7_39[0],stage7_38[0],stage7_37[0],stage7_36[1],stage7_35[1]}
   );
   gpc1325_5 gpc5865 (
      {stage6_37[3], stage6_37[4], stage6_37[5], stage6_37[6], stage6_37[7]},
      {stage6_38[1], 1'b0},
      {stage6_39[0], stage6_39[1], stage6_39[2]},
      {stage6_40[0]},
      {stage7_41[0],stage7_40[0],stage7_39[1],stage7_38[1],stage7_37[1]}
   );
   gpc223_4 gpc5866 (
      {stage6_41[0], stage6_41[1], 1'b0},
      {stage6_42[0], stage6_42[1]},
      {stage6_43[0], stage6_43[1]},
      {stage7_44[0],stage7_43[0],stage7_42[0],stage7_41[1]}
   );
   gpc1343_5 gpc5867 (
      {stage6_42[2], 1'b0, 1'b0},
      {stage6_43[2], stage6_43[3], stage6_43[4], stage6_43[5]},
      {stage6_44[0], stage6_44[1], stage6_44[2]},
      {stage6_45[0]},
      {stage7_46[0],stage7_45[0],stage7_44[1],stage7_43[1],stage7_42[1]}
   );
   gpc623_5 gpc5868 (
      {stage6_45[1], stage6_45[2], stage6_45[3]},
      {stage6_46[0], stage6_46[1]},
      {stage6_47[0], stage6_47[1], stage6_47[2], stage6_47[3], stage6_47[4], stage6_47[5]},
      {stage7_49[0],stage7_48[0],stage7_47[0],stage7_46[1],stage7_45[1]}
   );
   gpc2135_5 gpc5869 (
      {stage6_48[0], stage6_48[1], stage6_48[2], stage6_48[3], 1'b0},
      {stage6_49[0], stage6_49[1], stage6_49[2]},
      {stage6_50[0]},
      {stage6_51[0], stage6_51[1]},
      {stage7_52[0],stage7_51[0],stage7_50[0],stage7_49[1],stage7_48[1]}
   );
   gpc1343_5 gpc5870 (
      {stage6_50[1], stage6_50[2], stage6_50[3]},
      {stage6_51[2], stage6_51[3], stage6_51[4], 1'b0},
      {stage6_52[0], stage6_52[1], stage6_52[2]},
      {stage6_53[0]},
      {stage7_54[0],stage7_53[0],stage7_52[1],stage7_51[1],stage7_50[1]}
   );
   gpc1343_5 gpc5871 (
      {stage6_53[1], stage6_53[2], stage6_53[3]},
      {stage6_54[0], stage6_54[1], stage6_54[2], stage6_54[3]},
      {stage6_55[0], stage6_55[1], stage6_55[2]},
      {stage6_56[0]},
      {stage7_57[0],stage7_56[0],stage7_55[0],stage7_54[1],stage7_53[1]}
   );
   gpc135_4 gpc5872 (
      {stage6_56[1], stage6_56[2], stage6_56[3], stage6_56[4], stage6_56[5]},
      {stage6_57[0], stage6_57[1], stage6_57[2]},
      {stage6_58[0]},
      {stage7_59[0],stage7_58[0],stage7_57[1],stage7_56[1]}
   );
   gpc1406_5 gpc5873 (
      {stage6_59[0], stage6_59[1], stage6_59[2], stage6_59[3], stage6_59[4], stage6_59[5]},
      {stage6_61[0], stage6_61[1], stage6_61[2], stage6_61[3]},
      {stage6_62[0]},
      {stage7_63[0],stage7_62[0],stage7_61[0],stage7_60[0],stage7_59[1]}
   );
   gpc1415_5 gpc5874 (
      {stage6_60[0], stage6_60[1], stage6_60[2], stage6_60[3], stage6_60[4]},
      {stage6_61[4]},
      {stage6_62[1], stage6_62[2], stage6_62[3], stage6_62[4]},
      {stage6_63[0]},
      {stage7_64[0],stage7_63[1],stage7_62[1],stage7_61[1],stage7_60[1]}
   );
   gpc23_3 gpc5875 (
      {stage6_64[0], stage6_64[1], 1'b0},
      {stage6_65[0], stage6_65[1]},
      {stage7_66[0],stage7_65[0],stage7_64[1]}
   );
   gpc1343_5 gpc5876 (
      {stage6_66[0], stage6_66[1], stage6_66[2]},
      {stage6_67[0], stage6_67[1], stage6_67[2], stage6_67[3]},
      {stage6_68[0], stage6_68[1], stage6_68[2]},
      {stage6_69[0]},
      {stage7_70[0],stage7_69[0],stage7_68[0],stage7_67[0],stage7_66[1]}
   );
   gpc2223_5 gpc5877 (
      {1'b0, 1'b0, 1'b0},
      {stage6_69[1], 1'b0},
      {stage6_70[0], stage6_70[1]},
      {stage6_71[0], 1'b0},
      {stage7_71[0],stage7_70[1],stage7_69[1],stage7_68[1]}
   );
   gpc1_1 gpc5878 (
      {stage6_1[3]},
      {stage7_1[1]}
   );
   gpc1_1 gpc5879 (
      {stage6_4[4]},
      {stage7_4[1]}
   );
   gpc1_1 gpc5880 (
      {stage6_5[3]},
      {stage7_5[1]}
   );
   gpc1_1 gpc5881 (
      {stage6_6[1]},
      {stage7_6[1]}
   );
   gpc1_1 gpc5882 (
      {stage6_8[2]},
      {stage7_8[1]}
   );
   gpc1_1 gpc5883 (
      {stage6_14[6]},
      {stage7_14[1]}
   );
   gpc1_1 gpc5884 (
      {stage6_17[2]},
      {stage7_17[1]}
   );
   gpc1_1 gpc5885 (
      {stage6_20[3]},
      {stage7_20[1]}
   );
   gpc1_1 gpc5886 (
      {stage6_21[1]},
      {stage7_21[1]}
   );
   gpc1_1 gpc5887 (
      {stage6_24[1]},
      {stage7_24[1]}
   );
   gpc1_1 gpc5888 (
      {stage6_28[1]},
      {stage7_28[1]}
   );
   gpc1_1 gpc5889 (
      {stage6_30[2]},
      {stage7_30[1]}
   );
   gpc1_1 gpc5890 (
      {stage6_40[1]},
      {stage7_40[1]}
   );
   gpc1_1 gpc5891 (
      {stage6_55[3]},
      {stage7_55[1]}
   );
   gpc1_1 gpc5892 (
      {stage6_58[1]},
      {stage7_58[1]}
   );
   gpc1_1 gpc5893 (
      {stage6_67[4]},
      {stage7_67[1]}
   );
endmodule

module testbench();
    reg [255:0] src0;
    reg [255:0] src1;
    reg [255:0] src2;
    reg [255:0] src3;
    reg [255:0] src4;
    reg [255:0] src5;
    reg [255:0] src6;
    reg [255:0] src7;
    reg [255:0] src8;
    reg [255:0] src9;
    reg [255:0] src10;
    reg [255:0] src11;
    reg [255:0] src12;
    reg [255:0] src13;
    reg [255:0] src14;
    reg [255:0] src15;
    reg [255:0] src16;
    reg [255:0] src17;
    reg [255:0] src18;
    reg [255:0] src19;
    reg [255:0] src20;
    reg [255:0] src21;
    reg [255:0] src22;
    reg [255:0] src23;
    reg [255:0] src24;
    reg [255:0] src25;
    reg [255:0] src26;
    reg [255:0] src27;
    reg [255:0] src28;
    reg [255:0] src29;
    reg [255:0] src30;
    reg [255:0] src31;
    reg [255:0] src32;
    reg [255:0] src33;
    reg [255:0] src34;
    reg [255:0] src35;
    reg [255:0] src36;
    reg [255:0] src37;
    reg [255:0] src38;
    reg [255:0] src39;
    reg [255:0] src40;
    reg [255:0] src41;
    reg [255:0] src42;
    reg [255:0] src43;
    reg [255:0] src44;
    reg [255:0] src45;
    reg [255:0] src46;
    reg [255:0] src47;
    reg [255:0] src48;
    reg [255:0] src49;
    reg [255:0] src50;
    reg [255:0] src51;
    reg [255:0] src52;
    reg [255:0] src53;
    reg [255:0] src54;
    reg [255:0] src55;
    reg [255:0] src56;
    reg [255:0] src57;
    reg [255:0] src58;
    reg [255:0] src59;
    reg [255:0] src60;
    reg [255:0] src61;
    reg [255:0] src62;
    reg [255:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [0:0] dst71;
    wire [71:0] srcsum;
    wire [71:0] dstsum;
    wire test;
    compressor_CLA256_64 compressor_CLA256_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70),
        .dst71(dst71));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127] + src16[128] + src16[129] + src16[130] + src16[131] + src16[132] + src16[133] + src16[134] + src16[135] + src16[136] + src16[137] + src16[138] + src16[139] + src16[140] + src16[141] + src16[142] + src16[143] + src16[144] + src16[145] + src16[146] + src16[147] + src16[148] + src16[149] + src16[150] + src16[151] + src16[152] + src16[153] + src16[154] + src16[155] + src16[156] + src16[157] + src16[158] + src16[159] + src16[160] + src16[161] + src16[162] + src16[163] + src16[164] + src16[165] + src16[166] + src16[167] + src16[168] + src16[169] + src16[170] + src16[171] + src16[172] + src16[173] + src16[174] + src16[175] + src16[176] + src16[177] + src16[178] + src16[179] + src16[180] + src16[181] + src16[182] + src16[183] + src16[184] + src16[185] + src16[186] + src16[187] + src16[188] + src16[189] + src16[190] + src16[191] + src16[192] + src16[193] + src16[194] + src16[195] + src16[196] + src16[197] + src16[198] + src16[199] + src16[200] + src16[201] + src16[202] + src16[203] + src16[204] + src16[205] + src16[206] + src16[207] + src16[208] + src16[209] + src16[210] + src16[211] + src16[212] + src16[213] + src16[214] + src16[215] + src16[216] + src16[217] + src16[218] + src16[219] + src16[220] + src16[221] + src16[222] + src16[223] + src16[224] + src16[225] + src16[226] + src16[227] + src16[228] + src16[229] + src16[230] + src16[231] + src16[232] + src16[233] + src16[234] + src16[235] + src16[236] + src16[237] + src16[238] + src16[239] + src16[240] + src16[241] + src16[242] + src16[243] + src16[244] + src16[245] + src16[246] + src16[247] + src16[248] + src16[249] + src16[250] + src16[251] + src16[252] + src16[253] + src16[254] + src16[255])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127] + src17[128] + src17[129] + src17[130] + src17[131] + src17[132] + src17[133] + src17[134] + src17[135] + src17[136] + src17[137] + src17[138] + src17[139] + src17[140] + src17[141] + src17[142] + src17[143] + src17[144] + src17[145] + src17[146] + src17[147] + src17[148] + src17[149] + src17[150] + src17[151] + src17[152] + src17[153] + src17[154] + src17[155] + src17[156] + src17[157] + src17[158] + src17[159] + src17[160] + src17[161] + src17[162] + src17[163] + src17[164] + src17[165] + src17[166] + src17[167] + src17[168] + src17[169] + src17[170] + src17[171] + src17[172] + src17[173] + src17[174] + src17[175] + src17[176] + src17[177] + src17[178] + src17[179] + src17[180] + src17[181] + src17[182] + src17[183] + src17[184] + src17[185] + src17[186] + src17[187] + src17[188] + src17[189] + src17[190] + src17[191] + src17[192] + src17[193] + src17[194] + src17[195] + src17[196] + src17[197] + src17[198] + src17[199] + src17[200] + src17[201] + src17[202] + src17[203] + src17[204] + src17[205] + src17[206] + src17[207] + src17[208] + src17[209] + src17[210] + src17[211] + src17[212] + src17[213] + src17[214] + src17[215] + src17[216] + src17[217] + src17[218] + src17[219] + src17[220] + src17[221] + src17[222] + src17[223] + src17[224] + src17[225] + src17[226] + src17[227] + src17[228] + src17[229] + src17[230] + src17[231] + src17[232] + src17[233] + src17[234] + src17[235] + src17[236] + src17[237] + src17[238] + src17[239] + src17[240] + src17[241] + src17[242] + src17[243] + src17[244] + src17[245] + src17[246] + src17[247] + src17[248] + src17[249] + src17[250] + src17[251] + src17[252] + src17[253] + src17[254] + src17[255])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127] + src18[128] + src18[129] + src18[130] + src18[131] + src18[132] + src18[133] + src18[134] + src18[135] + src18[136] + src18[137] + src18[138] + src18[139] + src18[140] + src18[141] + src18[142] + src18[143] + src18[144] + src18[145] + src18[146] + src18[147] + src18[148] + src18[149] + src18[150] + src18[151] + src18[152] + src18[153] + src18[154] + src18[155] + src18[156] + src18[157] + src18[158] + src18[159] + src18[160] + src18[161] + src18[162] + src18[163] + src18[164] + src18[165] + src18[166] + src18[167] + src18[168] + src18[169] + src18[170] + src18[171] + src18[172] + src18[173] + src18[174] + src18[175] + src18[176] + src18[177] + src18[178] + src18[179] + src18[180] + src18[181] + src18[182] + src18[183] + src18[184] + src18[185] + src18[186] + src18[187] + src18[188] + src18[189] + src18[190] + src18[191] + src18[192] + src18[193] + src18[194] + src18[195] + src18[196] + src18[197] + src18[198] + src18[199] + src18[200] + src18[201] + src18[202] + src18[203] + src18[204] + src18[205] + src18[206] + src18[207] + src18[208] + src18[209] + src18[210] + src18[211] + src18[212] + src18[213] + src18[214] + src18[215] + src18[216] + src18[217] + src18[218] + src18[219] + src18[220] + src18[221] + src18[222] + src18[223] + src18[224] + src18[225] + src18[226] + src18[227] + src18[228] + src18[229] + src18[230] + src18[231] + src18[232] + src18[233] + src18[234] + src18[235] + src18[236] + src18[237] + src18[238] + src18[239] + src18[240] + src18[241] + src18[242] + src18[243] + src18[244] + src18[245] + src18[246] + src18[247] + src18[248] + src18[249] + src18[250] + src18[251] + src18[252] + src18[253] + src18[254] + src18[255])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127] + src19[128] + src19[129] + src19[130] + src19[131] + src19[132] + src19[133] + src19[134] + src19[135] + src19[136] + src19[137] + src19[138] + src19[139] + src19[140] + src19[141] + src19[142] + src19[143] + src19[144] + src19[145] + src19[146] + src19[147] + src19[148] + src19[149] + src19[150] + src19[151] + src19[152] + src19[153] + src19[154] + src19[155] + src19[156] + src19[157] + src19[158] + src19[159] + src19[160] + src19[161] + src19[162] + src19[163] + src19[164] + src19[165] + src19[166] + src19[167] + src19[168] + src19[169] + src19[170] + src19[171] + src19[172] + src19[173] + src19[174] + src19[175] + src19[176] + src19[177] + src19[178] + src19[179] + src19[180] + src19[181] + src19[182] + src19[183] + src19[184] + src19[185] + src19[186] + src19[187] + src19[188] + src19[189] + src19[190] + src19[191] + src19[192] + src19[193] + src19[194] + src19[195] + src19[196] + src19[197] + src19[198] + src19[199] + src19[200] + src19[201] + src19[202] + src19[203] + src19[204] + src19[205] + src19[206] + src19[207] + src19[208] + src19[209] + src19[210] + src19[211] + src19[212] + src19[213] + src19[214] + src19[215] + src19[216] + src19[217] + src19[218] + src19[219] + src19[220] + src19[221] + src19[222] + src19[223] + src19[224] + src19[225] + src19[226] + src19[227] + src19[228] + src19[229] + src19[230] + src19[231] + src19[232] + src19[233] + src19[234] + src19[235] + src19[236] + src19[237] + src19[238] + src19[239] + src19[240] + src19[241] + src19[242] + src19[243] + src19[244] + src19[245] + src19[246] + src19[247] + src19[248] + src19[249] + src19[250] + src19[251] + src19[252] + src19[253] + src19[254] + src19[255])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127] + src20[128] + src20[129] + src20[130] + src20[131] + src20[132] + src20[133] + src20[134] + src20[135] + src20[136] + src20[137] + src20[138] + src20[139] + src20[140] + src20[141] + src20[142] + src20[143] + src20[144] + src20[145] + src20[146] + src20[147] + src20[148] + src20[149] + src20[150] + src20[151] + src20[152] + src20[153] + src20[154] + src20[155] + src20[156] + src20[157] + src20[158] + src20[159] + src20[160] + src20[161] + src20[162] + src20[163] + src20[164] + src20[165] + src20[166] + src20[167] + src20[168] + src20[169] + src20[170] + src20[171] + src20[172] + src20[173] + src20[174] + src20[175] + src20[176] + src20[177] + src20[178] + src20[179] + src20[180] + src20[181] + src20[182] + src20[183] + src20[184] + src20[185] + src20[186] + src20[187] + src20[188] + src20[189] + src20[190] + src20[191] + src20[192] + src20[193] + src20[194] + src20[195] + src20[196] + src20[197] + src20[198] + src20[199] + src20[200] + src20[201] + src20[202] + src20[203] + src20[204] + src20[205] + src20[206] + src20[207] + src20[208] + src20[209] + src20[210] + src20[211] + src20[212] + src20[213] + src20[214] + src20[215] + src20[216] + src20[217] + src20[218] + src20[219] + src20[220] + src20[221] + src20[222] + src20[223] + src20[224] + src20[225] + src20[226] + src20[227] + src20[228] + src20[229] + src20[230] + src20[231] + src20[232] + src20[233] + src20[234] + src20[235] + src20[236] + src20[237] + src20[238] + src20[239] + src20[240] + src20[241] + src20[242] + src20[243] + src20[244] + src20[245] + src20[246] + src20[247] + src20[248] + src20[249] + src20[250] + src20[251] + src20[252] + src20[253] + src20[254] + src20[255])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127] + src21[128] + src21[129] + src21[130] + src21[131] + src21[132] + src21[133] + src21[134] + src21[135] + src21[136] + src21[137] + src21[138] + src21[139] + src21[140] + src21[141] + src21[142] + src21[143] + src21[144] + src21[145] + src21[146] + src21[147] + src21[148] + src21[149] + src21[150] + src21[151] + src21[152] + src21[153] + src21[154] + src21[155] + src21[156] + src21[157] + src21[158] + src21[159] + src21[160] + src21[161] + src21[162] + src21[163] + src21[164] + src21[165] + src21[166] + src21[167] + src21[168] + src21[169] + src21[170] + src21[171] + src21[172] + src21[173] + src21[174] + src21[175] + src21[176] + src21[177] + src21[178] + src21[179] + src21[180] + src21[181] + src21[182] + src21[183] + src21[184] + src21[185] + src21[186] + src21[187] + src21[188] + src21[189] + src21[190] + src21[191] + src21[192] + src21[193] + src21[194] + src21[195] + src21[196] + src21[197] + src21[198] + src21[199] + src21[200] + src21[201] + src21[202] + src21[203] + src21[204] + src21[205] + src21[206] + src21[207] + src21[208] + src21[209] + src21[210] + src21[211] + src21[212] + src21[213] + src21[214] + src21[215] + src21[216] + src21[217] + src21[218] + src21[219] + src21[220] + src21[221] + src21[222] + src21[223] + src21[224] + src21[225] + src21[226] + src21[227] + src21[228] + src21[229] + src21[230] + src21[231] + src21[232] + src21[233] + src21[234] + src21[235] + src21[236] + src21[237] + src21[238] + src21[239] + src21[240] + src21[241] + src21[242] + src21[243] + src21[244] + src21[245] + src21[246] + src21[247] + src21[248] + src21[249] + src21[250] + src21[251] + src21[252] + src21[253] + src21[254] + src21[255])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127] + src22[128] + src22[129] + src22[130] + src22[131] + src22[132] + src22[133] + src22[134] + src22[135] + src22[136] + src22[137] + src22[138] + src22[139] + src22[140] + src22[141] + src22[142] + src22[143] + src22[144] + src22[145] + src22[146] + src22[147] + src22[148] + src22[149] + src22[150] + src22[151] + src22[152] + src22[153] + src22[154] + src22[155] + src22[156] + src22[157] + src22[158] + src22[159] + src22[160] + src22[161] + src22[162] + src22[163] + src22[164] + src22[165] + src22[166] + src22[167] + src22[168] + src22[169] + src22[170] + src22[171] + src22[172] + src22[173] + src22[174] + src22[175] + src22[176] + src22[177] + src22[178] + src22[179] + src22[180] + src22[181] + src22[182] + src22[183] + src22[184] + src22[185] + src22[186] + src22[187] + src22[188] + src22[189] + src22[190] + src22[191] + src22[192] + src22[193] + src22[194] + src22[195] + src22[196] + src22[197] + src22[198] + src22[199] + src22[200] + src22[201] + src22[202] + src22[203] + src22[204] + src22[205] + src22[206] + src22[207] + src22[208] + src22[209] + src22[210] + src22[211] + src22[212] + src22[213] + src22[214] + src22[215] + src22[216] + src22[217] + src22[218] + src22[219] + src22[220] + src22[221] + src22[222] + src22[223] + src22[224] + src22[225] + src22[226] + src22[227] + src22[228] + src22[229] + src22[230] + src22[231] + src22[232] + src22[233] + src22[234] + src22[235] + src22[236] + src22[237] + src22[238] + src22[239] + src22[240] + src22[241] + src22[242] + src22[243] + src22[244] + src22[245] + src22[246] + src22[247] + src22[248] + src22[249] + src22[250] + src22[251] + src22[252] + src22[253] + src22[254] + src22[255])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127] + src23[128] + src23[129] + src23[130] + src23[131] + src23[132] + src23[133] + src23[134] + src23[135] + src23[136] + src23[137] + src23[138] + src23[139] + src23[140] + src23[141] + src23[142] + src23[143] + src23[144] + src23[145] + src23[146] + src23[147] + src23[148] + src23[149] + src23[150] + src23[151] + src23[152] + src23[153] + src23[154] + src23[155] + src23[156] + src23[157] + src23[158] + src23[159] + src23[160] + src23[161] + src23[162] + src23[163] + src23[164] + src23[165] + src23[166] + src23[167] + src23[168] + src23[169] + src23[170] + src23[171] + src23[172] + src23[173] + src23[174] + src23[175] + src23[176] + src23[177] + src23[178] + src23[179] + src23[180] + src23[181] + src23[182] + src23[183] + src23[184] + src23[185] + src23[186] + src23[187] + src23[188] + src23[189] + src23[190] + src23[191] + src23[192] + src23[193] + src23[194] + src23[195] + src23[196] + src23[197] + src23[198] + src23[199] + src23[200] + src23[201] + src23[202] + src23[203] + src23[204] + src23[205] + src23[206] + src23[207] + src23[208] + src23[209] + src23[210] + src23[211] + src23[212] + src23[213] + src23[214] + src23[215] + src23[216] + src23[217] + src23[218] + src23[219] + src23[220] + src23[221] + src23[222] + src23[223] + src23[224] + src23[225] + src23[226] + src23[227] + src23[228] + src23[229] + src23[230] + src23[231] + src23[232] + src23[233] + src23[234] + src23[235] + src23[236] + src23[237] + src23[238] + src23[239] + src23[240] + src23[241] + src23[242] + src23[243] + src23[244] + src23[245] + src23[246] + src23[247] + src23[248] + src23[249] + src23[250] + src23[251] + src23[252] + src23[253] + src23[254] + src23[255])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127] + src24[128] + src24[129] + src24[130] + src24[131] + src24[132] + src24[133] + src24[134] + src24[135] + src24[136] + src24[137] + src24[138] + src24[139] + src24[140] + src24[141] + src24[142] + src24[143] + src24[144] + src24[145] + src24[146] + src24[147] + src24[148] + src24[149] + src24[150] + src24[151] + src24[152] + src24[153] + src24[154] + src24[155] + src24[156] + src24[157] + src24[158] + src24[159] + src24[160] + src24[161] + src24[162] + src24[163] + src24[164] + src24[165] + src24[166] + src24[167] + src24[168] + src24[169] + src24[170] + src24[171] + src24[172] + src24[173] + src24[174] + src24[175] + src24[176] + src24[177] + src24[178] + src24[179] + src24[180] + src24[181] + src24[182] + src24[183] + src24[184] + src24[185] + src24[186] + src24[187] + src24[188] + src24[189] + src24[190] + src24[191] + src24[192] + src24[193] + src24[194] + src24[195] + src24[196] + src24[197] + src24[198] + src24[199] + src24[200] + src24[201] + src24[202] + src24[203] + src24[204] + src24[205] + src24[206] + src24[207] + src24[208] + src24[209] + src24[210] + src24[211] + src24[212] + src24[213] + src24[214] + src24[215] + src24[216] + src24[217] + src24[218] + src24[219] + src24[220] + src24[221] + src24[222] + src24[223] + src24[224] + src24[225] + src24[226] + src24[227] + src24[228] + src24[229] + src24[230] + src24[231] + src24[232] + src24[233] + src24[234] + src24[235] + src24[236] + src24[237] + src24[238] + src24[239] + src24[240] + src24[241] + src24[242] + src24[243] + src24[244] + src24[245] + src24[246] + src24[247] + src24[248] + src24[249] + src24[250] + src24[251] + src24[252] + src24[253] + src24[254] + src24[255])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127] + src25[128] + src25[129] + src25[130] + src25[131] + src25[132] + src25[133] + src25[134] + src25[135] + src25[136] + src25[137] + src25[138] + src25[139] + src25[140] + src25[141] + src25[142] + src25[143] + src25[144] + src25[145] + src25[146] + src25[147] + src25[148] + src25[149] + src25[150] + src25[151] + src25[152] + src25[153] + src25[154] + src25[155] + src25[156] + src25[157] + src25[158] + src25[159] + src25[160] + src25[161] + src25[162] + src25[163] + src25[164] + src25[165] + src25[166] + src25[167] + src25[168] + src25[169] + src25[170] + src25[171] + src25[172] + src25[173] + src25[174] + src25[175] + src25[176] + src25[177] + src25[178] + src25[179] + src25[180] + src25[181] + src25[182] + src25[183] + src25[184] + src25[185] + src25[186] + src25[187] + src25[188] + src25[189] + src25[190] + src25[191] + src25[192] + src25[193] + src25[194] + src25[195] + src25[196] + src25[197] + src25[198] + src25[199] + src25[200] + src25[201] + src25[202] + src25[203] + src25[204] + src25[205] + src25[206] + src25[207] + src25[208] + src25[209] + src25[210] + src25[211] + src25[212] + src25[213] + src25[214] + src25[215] + src25[216] + src25[217] + src25[218] + src25[219] + src25[220] + src25[221] + src25[222] + src25[223] + src25[224] + src25[225] + src25[226] + src25[227] + src25[228] + src25[229] + src25[230] + src25[231] + src25[232] + src25[233] + src25[234] + src25[235] + src25[236] + src25[237] + src25[238] + src25[239] + src25[240] + src25[241] + src25[242] + src25[243] + src25[244] + src25[245] + src25[246] + src25[247] + src25[248] + src25[249] + src25[250] + src25[251] + src25[252] + src25[253] + src25[254] + src25[255])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127] + src26[128] + src26[129] + src26[130] + src26[131] + src26[132] + src26[133] + src26[134] + src26[135] + src26[136] + src26[137] + src26[138] + src26[139] + src26[140] + src26[141] + src26[142] + src26[143] + src26[144] + src26[145] + src26[146] + src26[147] + src26[148] + src26[149] + src26[150] + src26[151] + src26[152] + src26[153] + src26[154] + src26[155] + src26[156] + src26[157] + src26[158] + src26[159] + src26[160] + src26[161] + src26[162] + src26[163] + src26[164] + src26[165] + src26[166] + src26[167] + src26[168] + src26[169] + src26[170] + src26[171] + src26[172] + src26[173] + src26[174] + src26[175] + src26[176] + src26[177] + src26[178] + src26[179] + src26[180] + src26[181] + src26[182] + src26[183] + src26[184] + src26[185] + src26[186] + src26[187] + src26[188] + src26[189] + src26[190] + src26[191] + src26[192] + src26[193] + src26[194] + src26[195] + src26[196] + src26[197] + src26[198] + src26[199] + src26[200] + src26[201] + src26[202] + src26[203] + src26[204] + src26[205] + src26[206] + src26[207] + src26[208] + src26[209] + src26[210] + src26[211] + src26[212] + src26[213] + src26[214] + src26[215] + src26[216] + src26[217] + src26[218] + src26[219] + src26[220] + src26[221] + src26[222] + src26[223] + src26[224] + src26[225] + src26[226] + src26[227] + src26[228] + src26[229] + src26[230] + src26[231] + src26[232] + src26[233] + src26[234] + src26[235] + src26[236] + src26[237] + src26[238] + src26[239] + src26[240] + src26[241] + src26[242] + src26[243] + src26[244] + src26[245] + src26[246] + src26[247] + src26[248] + src26[249] + src26[250] + src26[251] + src26[252] + src26[253] + src26[254] + src26[255])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127] + src27[128] + src27[129] + src27[130] + src27[131] + src27[132] + src27[133] + src27[134] + src27[135] + src27[136] + src27[137] + src27[138] + src27[139] + src27[140] + src27[141] + src27[142] + src27[143] + src27[144] + src27[145] + src27[146] + src27[147] + src27[148] + src27[149] + src27[150] + src27[151] + src27[152] + src27[153] + src27[154] + src27[155] + src27[156] + src27[157] + src27[158] + src27[159] + src27[160] + src27[161] + src27[162] + src27[163] + src27[164] + src27[165] + src27[166] + src27[167] + src27[168] + src27[169] + src27[170] + src27[171] + src27[172] + src27[173] + src27[174] + src27[175] + src27[176] + src27[177] + src27[178] + src27[179] + src27[180] + src27[181] + src27[182] + src27[183] + src27[184] + src27[185] + src27[186] + src27[187] + src27[188] + src27[189] + src27[190] + src27[191] + src27[192] + src27[193] + src27[194] + src27[195] + src27[196] + src27[197] + src27[198] + src27[199] + src27[200] + src27[201] + src27[202] + src27[203] + src27[204] + src27[205] + src27[206] + src27[207] + src27[208] + src27[209] + src27[210] + src27[211] + src27[212] + src27[213] + src27[214] + src27[215] + src27[216] + src27[217] + src27[218] + src27[219] + src27[220] + src27[221] + src27[222] + src27[223] + src27[224] + src27[225] + src27[226] + src27[227] + src27[228] + src27[229] + src27[230] + src27[231] + src27[232] + src27[233] + src27[234] + src27[235] + src27[236] + src27[237] + src27[238] + src27[239] + src27[240] + src27[241] + src27[242] + src27[243] + src27[244] + src27[245] + src27[246] + src27[247] + src27[248] + src27[249] + src27[250] + src27[251] + src27[252] + src27[253] + src27[254] + src27[255])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127] + src28[128] + src28[129] + src28[130] + src28[131] + src28[132] + src28[133] + src28[134] + src28[135] + src28[136] + src28[137] + src28[138] + src28[139] + src28[140] + src28[141] + src28[142] + src28[143] + src28[144] + src28[145] + src28[146] + src28[147] + src28[148] + src28[149] + src28[150] + src28[151] + src28[152] + src28[153] + src28[154] + src28[155] + src28[156] + src28[157] + src28[158] + src28[159] + src28[160] + src28[161] + src28[162] + src28[163] + src28[164] + src28[165] + src28[166] + src28[167] + src28[168] + src28[169] + src28[170] + src28[171] + src28[172] + src28[173] + src28[174] + src28[175] + src28[176] + src28[177] + src28[178] + src28[179] + src28[180] + src28[181] + src28[182] + src28[183] + src28[184] + src28[185] + src28[186] + src28[187] + src28[188] + src28[189] + src28[190] + src28[191] + src28[192] + src28[193] + src28[194] + src28[195] + src28[196] + src28[197] + src28[198] + src28[199] + src28[200] + src28[201] + src28[202] + src28[203] + src28[204] + src28[205] + src28[206] + src28[207] + src28[208] + src28[209] + src28[210] + src28[211] + src28[212] + src28[213] + src28[214] + src28[215] + src28[216] + src28[217] + src28[218] + src28[219] + src28[220] + src28[221] + src28[222] + src28[223] + src28[224] + src28[225] + src28[226] + src28[227] + src28[228] + src28[229] + src28[230] + src28[231] + src28[232] + src28[233] + src28[234] + src28[235] + src28[236] + src28[237] + src28[238] + src28[239] + src28[240] + src28[241] + src28[242] + src28[243] + src28[244] + src28[245] + src28[246] + src28[247] + src28[248] + src28[249] + src28[250] + src28[251] + src28[252] + src28[253] + src28[254] + src28[255])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127] + src29[128] + src29[129] + src29[130] + src29[131] + src29[132] + src29[133] + src29[134] + src29[135] + src29[136] + src29[137] + src29[138] + src29[139] + src29[140] + src29[141] + src29[142] + src29[143] + src29[144] + src29[145] + src29[146] + src29[147] + src29[148] + src29[149] + src29[150] + src29[151] + src29[152] + src29[153] + src29[154] + src29[155] + src29[156] + src29[157] + src29[158] + src29[159] + src29[160] + src29[161] + src29[162] + src29[163] + src29[164] + src29[165] + src29[166] + src29[167] + src29[168] + src29[169] + src29[170] + src29[171] + src29[172] + src29[173] + src29[174] + src29[175] + src29[176] + src29[177] + src29[178] + src29[179] + src29[180] + src29[181] + src29[182] + src29[183] + src29[184] + src29[185] + src29[186] + src29[187] + src29[188] + src29[189] + src29[190] + src29[191] + src29[192] + src29[193] + src29[194] + src29[195] + src29[196] + src29[197] + src29[198] + src29[199] + src29[200] + src29[201] + src29[202] + src29[203] + src29[204] + src29[205] + src29[206] + src29[207] + src29[208] + src29[209] + src29[210] + src29[211] + src29[212] + src29[213] + src29[214] + src29[215] + src29[216] + src29[217] + src29[218] + src29[219] + src29[220] + src29[221] + src29[222] + src29[223] + src29[224] + src29[225] + src29[226] + src29[227] + src29[228] + src29[229] + src29[230] + src29[231] + src29[232] + src29[233] + src29[234] + src29[235] + src29[236] + src29[237] + src29[238] + src29[239] + src29[240] + src29[241] + src29[242] + src29[243] + src29[244] + src29[245] + src29[246] + src29[247] + src29[248] + src29[249] + src29[250] + src29[251] + src29[252] + src29[253] + src29[254] + src29[255])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127] + src30[128] + src30[129] + src30[130] + src30[131] + src30[132] + src30[133] + src30[134] + src30[135] + src30[136] + src30[137] + src30[138] + src30[139] + src30[140] + src30[141] + src30[142] + src30[143] + src30[144] + src30[145] + src30[146] + src30[147] + src30[148] + src30[149] + src30[150] + src30[151] + src30[152] + src30[153] + src30[154] + src30[155] + src30[156] + src30[157] + src30[158] + src30[159] + src30[160] + src30[161] + src30[162] + src30[163] + src30[164] + src30[165] + src30[166] + src30[167] + src30[168] + src30[169] + src30[170] + src30[171] + src30[172] + src30[173] + src30[174] + src30[175] + src30[176] + src30[177] + src30[178] + src30[179] + src30[180] + src30[181] + src30[182] + src30[183] + src30[184] + src30[185] + src30[186] + src30[187] + src30[188] + src30[189] + src30[190] + src30[191] + src30[192] + src30[193] + src30[194] + src30[195] + src30[196] + src30[197] + src30[198] + src30[199] + src30[200] + src30[201] + src30[202] + src30[203] + src30[204] + src30[205] + src30[206] + src30[207] + src30[208] + src30[209] + src30[210] + src30[211] + src30[212] + src30[213] + src30[214] + src30[215] + src30[216] + src30[217] + src30[218] + src30[219] + src30[220] + src30[221] + src30[222] + src30[223] + src30[224] + src30[225] + src30[226] + src30[227] + src30[228] + src30[229] + src30[230] + src30[231] + src30[232] + src30[233] + src30[234] + src30[235] + src30[236] + src30[237] + src30[238] + src30[239] + src30[240] + src30[241] + src30[242] + src30[243] + src30[244] + src30[245] + src30[246] + src30[247] + src30[248] + src30[249] + src30[250] + src30[251] + src30[252] + src30[253] + src30[254] + src30[255])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127] + src31[128] + src31[129] + src31[130] + src31[131] + src31[132] + src31[133] + src31[134] + src31[135] + src31[136] + src31[137] + src31[138] + src31[139] + src31[140] + src31[141] + src31[142] + src31[143] + src31[144] + src31[145] + src31[146] + src31[147] + src31[148] + src31[149] + src31[150] + src31[151] + src31[152] + src31[153] + src31[154] + src31[155] + src31[156] + src31[157] + src31[158] + src31[159] + src31[160] + src31[161] + src31[162] + src31[163] + src31[164] + src31[165] + src31[166] + src31[167] + src31[168] + src31[169] + src31[170] + src31[171] + src31[172] + src31[173] + src31[174] + src31[175] + src31[176] + src31[177] + src31[178] + src31[179] + src31[180] + src31[181] + src31[182] + src31[183] + src31[184] + src31[185] + src31[186] + src31[187] + src31[188] + src31[189] + src31[190] + src31[191] + src31[192] + src31[193] + src31[194] + src31[195] + src31[196] + src31[197] + src31[198] + src31[199] + src31[200] + src31[201] + src31[202] + src31[203] + src31[204] + src31[205] + src31[206] + src31[207] + src31[208] + src31[209] + src31[210] + src31[211] + src31[212] + src31[213] + src31[214] + src31[215] + src31[216] + src31[217] + src31[218] + src31[219] + src31[220] + src31[221] + src31[222] + src31[223] + src31[224] + src31[225] + src31[226] + src31[227] + src31[228] + src31[229] + src31[230] + src31[231] + src31[232] + src31[233] + src31[234] + src31[235] + src31[236] + src31[237] + src31[238] + src31[239] + src31[240] + src31[241] + src31[242] + src31[243] + src31[244] + src31[245] + src31[246] + src31[247] + src31[248] + src31[249] + src31[250] + src31[251] + src31[252] + src31[253] + src31[254] + src31[255])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127] + src32[128] + src32[129] + src32[130] + src32[131] + src32[132] + src32[133] + src32[134] + src32[135] + src32[136] + src32[137] + src32[138] + src32[139] + src32[140] + src32[141] + src32[142] + src32[143] + src32[144] + src32[145] + src32[146] + src32[147] + src32[148] + src32[149] + src32[150] + src32[151] + src32[152] + src32[153] + src32[154] + src32[155] + src32[156] + src32[157] + src32[158] + src32[159] + src32[160] + src32[161] + src32[162] + src32[163] + src32[164] + src32[165] + src32[166] + src32[167] + src32[168] + src32[169] + src32[170] + src32[171] + src32[172] + src32[173] + src32[174] + src32[175] + src32[176] + src32[177] + src32[178] + src32[179] + src32[180] + src32[181] + src32[182] + src32[183] + src32[184] + src32[185] + src32[186] + src32[187] + src32[188] + src32[189] + src32[190] + src32[191] + src32[192] + src32[193] + src32[194] + src32[195] + src32[196] + src32[197] + src32[198] + src32[199] + src32[200] + src32[201] + src32[202] + src32[203] + src32[204] + src32[205] + src32[206] + src32[207] + src32[208] + src32[209] + src32[210] + src32[211] + src32[212] + src32[213] + src32[214] + src32[215] + src32[216] + src32[217] + src32[218] + src32[219] + src32[220] + src32[221] + src32[222] + src32[223] + src32[224] + src32[225] + src32[226] + src32[227] + src32[228] + src32[229] + src32[230] + src32[231] + src32[232] + src32[233] + src32[234] + src32[235] + src32[236] + src32[237] + src32[238] + src32[239] + src32[240] + src32[241] + src32[242] + src32[243] + src32[244] + src32[245] + src32[246] + src32[247] + src32[248] + src32[249] + src32[250] + src32[251] + src32[252] + src32[253] + src32[254] + src32[255])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127] + src33[128] + src33[129] + src33[130] + src33[131] + src33[132] + src33[133] + src33[134] + src33[135] + src33[136] + src33[137] + src33[138] + src33[139] + src33[140] + src33[141] + src33[142] + src33[143] + src33[144] + src33[145] + src33[146] + src33[147] + src33[148] + src33[149] + src33[150] + src33[151] + src33[152] + src33[153] + src33[154] + src33[155] + src33[156] + src33[157] + src33[158] + src33[159] + src33[160] + src33[161] + src33[162] + src33[163] + src33[164] + src33[165] + src33[166] + src33[167] + src33[168] + src33[169] + src33[170] + src33[171] + src33[172] + src33[173] + src33[174] + src33[175] + src33[176] + src33[177] + src33[178] + src33[179] + src33[180] + src33[181] + src33[182] + src33[183] + src33[184] + src33[185] + src33[186] + src33[187] + src33[188] + src33[189] + src33[190] + src33[191] + src33[192] + src33[193] + src33[194] + src33[195] + src33[196] + src33[197] + src33[198] + src33[199] + src33[200] + src33[201] + src33[202] + src33[203] + src33[204] + src33[205] + src33[206] + src33[207] + src33[208] + src33[209] + src33[210] + src33[211] + src33[212] + src33[213] + src33[214] + src33[215] + src33[216] + src33[217] + src33[218] + src33[219] + src33[220] + src33[221] + src33[222] + src33[223] + src33[224] + src33[225] + src33[226] + src33[227] + src33[228] + src33[229] + src33[230] + src33[231] + src33[232] + src33[233] + src33[234] + src33[235] + src33[236] + src33[237] + src33[238] + src33[239] + src33[240] + src33[241] + src33[242] + src33[243] + src33[244] + src33[245] + src33[246] + src33[247] + src33[248] + src33[249] + src33[250] + src33[251] + src33[252] + src33[253] + src33[254] + src33[255])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127] + src34[128] + src34[129] + src34[130] + src34[131] + src34[132] + src34[133] + src34[134] + src34[135] + src34[136] + src34[137] + src34[138] + src34[139] + src34[140] + src34[141] + src34[142] + src34[143] + src34[144] + src34[145] + src34[146] + src34[147] + src34[148] + src34[149] + src34[150] + src34[151] + src34[152] + src34[153] + src34[154] + src34[155] + src34[156] + src34[157] + src34[158] + src34[159] + src34[160] + src34[161] + src34[162] + src34[163] + src34[164] + src34[165] + src34[166] + src34[167] + src34[168] + src34[169] + src34[170] + src34[171] + src34[172] + src34[173] + src34[174] + src34[175] + src34[176] + src34[177] + src34[178] + src34[179] + src34[180] + src34[181] + src34[182] + src34[183] + src34[184] + src34[185] + src34[186] + src34[187] + src34[188] + src34[189] + src34[190] + src34[191] + src34[192] + src34[193] + src34[194] + src34[195] + src34[196] + src34[197] + src34[198] + src34[199] + src34[200] + src34[201] + src34[202] + src34[203] + src34[204] + src34[205] + src34[206] + src34[207] + src34[208] + src34[209] + src34[210] + src34[211] + src34[212] + src34[213] + src34[214] + src34[215] + src34[216] + src34[217] + src34[218] + src34[219] + src34[220] + src34[221] + src34[222] + src34[223] + src34[224] + src34[225] + src34[226] + src34[227] + src34[228] + src34[229] + src34[230] + src34[231] + src34[232] + src34[233] + src34[234] + src34[235] + src34[236] + src34[237] + src34[238] + src34[239] + src34[240] + src34[241] + src34[242] + src34[243] + src34[244] + src34[245] + src34[246] + src34[247] + src34[248] + src34[249] + src34[250] + src34[251] + src34[252] + src34[253] + src34[254] + src34[255])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127] + src35[128] + src35[129] + src35[130] + src35[131] + src35[132] + src35[133] + src35[134] + src35[135] + src35[136] + src35[137] + src35[138] + src35[139] + src35[140] + src35[141] + src35[142] + src35[143] + src35[144] + src35[145] + src35[146] + src35[147] + src35[148] + src35[149] + src35[150] + src35[151] + src35[152] + src35[153] + src35[154] + src35[155] + src35[156] + src35[157] + src35[158] + src35[159] + src35[160] + src35[161] + src35[162] + src35[163] + src35[164] + src35[165] + src35[166] + src35[167] + src35[168] + src35[169] + src35[170] + src35[171] + src35[172] + src35[173] + src35[174] + src35[175] + src35[176] + src35[177] + src35[178] + src35[179] + src35[180] + src35[181] + src35[182] + src35[183] + src35[184] + src35[185] + src35[186] + src35[187] + src35[188] + src35[189] + src35[190] + src35[191] + src35[192] + src35[193] + src35[194] + src35[195] + src35[196] + src35[197] + src35[198] + src35[199] + src35[200] + src35[201] + src35[202] + src35[203] + src35[204] + src35[205] + src35[206] + src35[207] + src35[208] + src35[209] + src35[210] + src35[211] + src35[212] + src35[213] + src35[214] + src35[215] + src35[216] + src35[217] + src35[218] + src35[219] + src35[220] + src35[221] + src35[222] + src35[223] + src35[224] + src35[225] + src35[226] + src35[227] + src35[228] + src35[229] + src35[230] + src35[231] + src35[232] + src35[233] + src35[234] + src35[235] + src35[236] + src35[237] + src35[238] + src35[239] + src35[240] + src35[241] + src35[242] + src35[243] + src35[244] + src35[245] + src35[246] + src35[247] + src35[248] + src35[249] + src35[250] + src35[251] + src35[252] + src35[253] + src35[254] + src35[255])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127] + src36[128] + src36[129] + src36[130] + src36[131] + src36[132] + src36[133] + src36[134] + src36[135] + src36[136] + src36[137] + src36[138] + src36[139] + src36[140] + src36[141] + src36[142] + src36[143] + src36[144] + src36[145] + src36[146] + src36[147] + src36[148] + src36[149] + src36[150] + src36[151] + src36[152] + src36[153] + src36[154] + src36[155] + src36[156] + src36[157] + src36[158] + src36[159] + src36[160] + src36[161] + src36[162] + src36[163] + src36[164] + src36[165] + src36[166] + src36[167] + src36[168] + src36[169] + src36[170] + src36[171] + src36[172] + src36[173] + src36[174] + src36[175] + src36[176] + src36[177] + src36[178] + src36[179] + src36[180] + src36[181] + src36[182] + src36[183] + src36[184] + src36[185] + src36[186] + src36[187] + src36[188] + src36[189] + src36[190] + src36[191] + src36[192] + src36[193] + src36[194] + src36[195] + src36[196] + src36[197] + src36[198] + src36[199] + src36[200] + src36[201] + src36[202] + src36[203] + src36[204] + src36[205] + src36[206] + src36[207] + src36[208] + src36[209] + src36[210] + src36[211] + src36[212] + src36[213] + src36[214] + src36[215] + src36[216] + src36[217] + src36[218] + src36[219] + src36[220] + src36[221] + src36[222] + src36[223] + src36[224] + src36[225] + src36[226] + src36[227] + src36[228] + src36[229] + src36[230] + src36[231] + src36[232] + src36[233] + src36[234] + src36[235] + src36[236] + src36[237] + src36[238] + src36[239] + src36[240] + src36[241] + src36[242] + src36[243] + src36[244] + src36[245] + src36[246] + src36[247] + src36[248] + src36[249] + src36[250] + src36[251] + src36[252] + src36[253] + src36[254] + src36[255])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127] + src37[128] + src37[129] + src37[130] + src37[131] + src37[132] + src37[133] + src37[134] + src37[135] + src37[136] + src37[137] + src37[138] + src37[139] + src37[140] + src37[141] + src37[142] + src37[143] + src37[144] + src37[145] + src37[146] + src37[147] + src37[148] + src37[149] + src37[150] + src37[151] + src37[152] + src37[153] + src37[154] + src37[155] + src37[156] + src37[157] + src37[158] + src37[159] + src37[160] + src37[161] + src37[162] + src37[163] + src37[164] + src37[165] + src37[166] + src37[167] + src37[168] + src37[169] + src37[170] + src37[171] + src37[172] + src37[173] + src37[174] + src37[175] + src37[176] + src37[177] + src37[178] + src37[179] + src37[180] + src37[181] + src37[182] + src37[183] + src37[184] + src37[185] + src37[186] + src37[187] + src37[188] + src37[189] + src37[190] + src37[191] + src37[192] + src37[193] + src37[194] + src37[195] + src37[196] + src37[197] + src37[198] + src37[199] + src37[200] + src37[201] + src37[202] + src37[203] + src37[204] + src37[205] + src37[206] + src37[207] + src37[208] + src37[209] + src37[210] + src37[211] + src37[212] + src37[213] + src37[214] + src37[215] + src37[216] + src37[217] + src37[218] + src37[219] + src37[220] + src37[221] + src37[222] + src37[223] + src37[224] + src37[225] + src37[226] + src37[227] + src37[228] + src37[229] + src37[230] + src37[231] + src37[232] + src37[233] + src37[234] + src37[235] + src37[236] + src37[237] + src37[238] + src37[239] + src37[240] + src37[241] + src37[242] + src37[243] + src37[244] + src37[245] + src37[246] + src37[247] + src37[248] + src37[249] + src37[250] + src37[251] + src37[252] + src37[253] + src37[254] + src37[255])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127] + src38[128] + src38[129] + src38[130] + src38[131] + src38[132] + src38[133] + src38[134] + src38[135] + src38[136] + src38[137] + src38[138] + src38[139] + src38[140] + src38[141] + src38[142] + src38[143] + src38[144] + src38[145] + src38[146] + src38[147] + src38[148] + src38[149] + src38[150] + src38[151] + src38[152] + src38[153] + src38[154] + src38[155] + src38[156] + src38[157] + src38[158] + src38[159] + src38[160] + src38[161] + src38[162] + src38[163] + src38[164] + src38[165] + src38[166] + src38[167] + src38[168] + src38[169] + src38[170] + src38[171] + src38[172] + src38[173] + src38[174] + src38[175] + src38[176] + src38[177] + src38[178] + src38[179] + src38[180] + src38[181] + src38[182] + src38[183] + src38[184] + src38[185] + src38[186] + src38[187] + src38[188] + src38[189] + src38[190] + src38[191] + src38[192] + src38[193] + src38[194] + src38[195] + src38[196] + src38[197] + src38[198] + src38[199] + src38[200] + src38[201] + src38[202] + src38[203] + src38[204] + src38[205] + src38[206] + src38[207] + src38[208] + src38[209] + src38[210] + src38[211] + src38[212] + src38[213] + src38[214] + src38[215] + src38[216] + src38[217] + src38[218] + src38[219] + src38[220] + src38[221] + src38[222] + src38[223] + src38[224] + src38[225] + src38[226] + src38[227] + src38[228] + src38[229] + src38[230] + src38[231] + src38[232] + src38[233] + src38[234] + src38[235] + src38[236] + src38[237] + src38[238] + src38[239] + src38[240] + src38[241] + src38[242] + src38[243] + src38[244] + src38[245] + src38[246] + src38[247] + src38[248] + src38[249] + src38[250] + src38[251] + src38[252] + src38[253] + src38[254] + src38[255])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127] + src39[128] + src39[129] + src39[130] + src39[131] + src39[132] + src39[133] + src39[134] + src39[135] + src39[136] + src39[137] + src39[138] + src39[139] + src39[140] + src39[141] + src39[142] + src39[143] + src39[144] + src39[145] + src39[146] + src39[147] + src39[148] + src39[149] + src39[150] + src39[151] + src39[152] + src39[153] + src39[154] + src39[155] + src39[156] + src39[157] + src39[158] + src39[159] + src39[160] + src39[161] + src39[162] + src39[163] + src39[164] + src39[165] + src39[166] + src39[167] + src39[168] + src39[169] + src39[170] + src39[171] + src39[172] + src39[173] + src39[174] + src39[175] + src39[176] + src39[177] + src39[178] + src39[179] + src39[180] + src39[181] + src39[182] + src39[183] + src39[184] + src39[185] + src39[186] + src39[187] + src39[188] + src39[189] + src39[190] + src39[191] + src39[192] + src39[193] + src39[194] + src39[195] + src39[196] + src39[197] + src39[198] + src39[199] + src39[200] + src39[201] + src39[202] + src39[203] + src39[204] + src39[205] + src39[206] + src39[207] + src39[208] + src39[209] + src39[210] + src39[211] + src39[212] + src39[213] + src39[214] + src39[215] + src39[216] + src39[217] + src39[218] + src39[219] + src39[220] + src39[221] + src39[222] + src39[223] + src39[224] + src39[225] + src39[226] + src39[227] + src39[228] + src39[229] + src39[230] + src39[231] + src39[232] + src39[233] + src39[234] + src39[235] + src39[236] + src39[237] + src39[238] + src39[239] + src39[240] + src39[241] + src39[242] + src39[243] + src39[244] + src39[245] + src39[246] + src39[247] + src39[248] + src39[249] + src39[250] + src39[251] + src39[252] + src39[253] + src39[254] + src39[255])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127] + src40[128] + src40[129] + src40[130] + src40[131] + src40[132] + src40[133] + src40[134] + src40[135] + src40[136] + src40[137] + src40[138] + src40[139] + src40[140] + src40[141] + src40[142] + src40[143] + src40[144] + src40[145] + src40[146] + src40[147] + src40[148] + src40[149] + src40[150] + src40[151] + src40[152] + src40[153] + src40[154] + src40[155] + src40[156] + src40[157] + src40[158] + src40[159] + src40[160] + src40[161] + src40[162] + src40[163] + src40[164] + src40[165] + src40[166] + src40[167] + src40[168] + src40[169] + src40[170] + src40[171] + src40[172] + src40[173] + src40[174] + src40[175] + src40[176] + src40[177] + src40[178] + src40[179] + src40[180] + src40[181] + src40[182] + src40[183] + src40[184] + src40[185] + src40[186] + src40[187] + src40[188] + src40[189] + src40[190] + src40[191] + src40[192] + src40[193] + src40[194] + src40[195] + src40[196] + src40[197] + src40[198] + src40[199] + src40[200] + src40[201] + src40[202] + src40[203] + src40[204] + src40[205] + src40[206] + src40[207] + src40[208] + src40[209] + src40[210] + src40[211] + src40[212] + src40[213] + src40[214] + src40[215] + src40[216] + src40[217] + src40[218] + src40[219] + src40[220] + src40[221] + src40[222] + src40[223] + src40[224] + src40[225] + src40[226] + src40[227] + src40[228] + src40[229] + src40[230] + src40[231] + src40[232] + src40[233] + src40[234] + src40[235] + src40[236] + src40[237] + src40[238] + src40[239] + src40[240] + src40[241] + src40[242] + src40[243] + src40[244] + src40[245] + src40[246] + src40[247] + src40[248] + src40[249] + src40[250] + src40[251] + src40[252] + src40[253] + src40[254] + src40[255])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127] + src41[128] + src41[129] + src41[130] + src41[131] + src41[132] + src41[133] + src41[134] + src41[135] + src41[136] + src41[137] + src41[138] + src41[139] + src41[140] + src41[141] + src41[142] + src41[143] + src41[144] + src41[145] + src41[146] + src41[147] + src41[148] + src41[149] + src41[150] + src41[151] + src41[152] + src41[153] + src41[154] + src41[155] + src41[156] + src41[157] + src41[158] + src41[159] + src41[160] + src41[161] + src41[162] + src41[163] + src41[164] + src41[165] + src41[166] + src41[167] + src41[168] + src41[169] + src41[170] + src41[171] + src41[172] + src41[173] + src41[174] + src41[175] + src41[176] + src41[177] + src41[178] + src41[179] + src41[180] + src41[181] + src41[182] + src41[183] + src41[184] + src41[185] + src41[186] + src41[187] + src41[188] + src41[189] + src41[190] + src41[191] + src41[192] + src41[193] + src41[194] + src41[195] + src41[196] + src41[197] + src41[198] + src41[199] + src41[200] + src41[201] + src41[202] + src41[203] + src41[204] + src41[205] + src41[206] + src41[207] + src41[208] + src41[209] + src41[210] + src41[211] + src41[212] + src41[213] + src41[214] + src41[215] + src41[216] + src41[217] + src41[218] + src41[219] + src41[220] + src41[221] + src41[222] + src41[223] + src41[224] + src41[225] + src41[226] + src41[227] + src41[228] + src41[229] + src41[230] + src41[231] + src41[232] + src41[233] + src41[234] + src41[235] + src41[236] + src41[237] + src41[238] + src41[239] + src41[240] + src41[241] + src41[242] + src41[243] + src41[244] + src41[245] + src41[246] + src41[247] + src41[248] + src41[249] + src41[250] + src41[251] + src41[252] + src41[253] + src41[254] + src41[255])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127] + src42[128] + src42[129] + src42[130] + src42[131] + src42[132] + src42[133] + src42[134] + src42[135] + src42[136] + src42[137] + src42[138] + src42[139] + src42[140] + src42[141] + src42[142] + src42[143] + src42[144] + src42[145] + src42[146] + src42[147] + src42[148] + src42[149] + src42[150] + src42[151] + src42[152] + src42[153] + src42[154] + src42[155] + src42[156] + src42[157] + src42[158] + src42[159] + src42[160] + src42[161] + src42[162] + src42[163] + src42[164] + src42[165] + src42[166] + src42[167] + src42[168] + src42[169] + src42[170] + src42[171] + src42[172] + src42[173] + src42[174] + src42[175] + src42[176] + src42[177] + src42[178] + src42[179] + src42[180] + src42[181] + src42[182] + src42[183] + src42[184] + src42[185] + src42[186] + src42[187] + src42[188] + src42[189] + src42[190] + src42[191] + src42[192] + src42[193] + src42[194] + src42[195] + src42[196] + src42[197] + src42[198] + src42[199] + src42[200] + src42[201] + src42[202] + src42[203] + src42[204] + src42[205] + src42[206] + src42[207] + src42[208] + src42[209] + src42[210] + src42[211] + src42[212] + src42[213] + src42[214] + src42[215] + src42[216] + src42[217] + src42[218] + src42[219] + src42[220] + src42[221] + src42[222] + src42[223] + src42[224] + src42[225] + src42[226] + src42[227] + src42[228] + src42[229] + src42[230] + src42[231] + src42[232] + src42[233] + src42[234] + src42[235] + src42[236] + src42[237] + src42[238] + src42[239] + src42[240] + src42[241] + src42[242] + src42[243] + src42[244] + src42[245] + src42[246] + src42[247] + src42[248] + src42[249] + src42[250] + src42[251] + src42[252] + src42[253] + src42[254] + src42[255])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127] + src43[128] + src43[129] + src43[130] + src43[131] + src43[132] + src43[133] + src43[134] + src43[135] + src43[136] + src43[137] + src43[138] + src43[139] + src43[140] + src43[141] + src43[142] + src43[143] + src43[144] + src43[145] + src43[146] + src43[147] + src43[148] + src43[149] + src43[150] + src43[151] + src43[152] + src43[153] + src43[154] + src43[155] + src43[156] + src43[157] + src43[158] + src43[159] + src43[160] + src43[161] + src43[162] + src43[163] + src43[164] + src43[165] + src43[166] + src43[167] + src43[168] + src43[169] + src43[170] + src43[171] + src43[172] + src43[173] + src43[174] + src43[175] + src43[176] + src43[177] + src43[178] + src43[179] + src43[180] + src43[181] + src43[182] + src43[183] + src43[184] + src43[185] + src43[186] + src43[187] + src43[188] + src43[189] + src43[190] + src43[191] + src43[192] + src43[193] + src43[194] + src43[195] + src43[196] + src43[197] + src43[198] + src43[199] + src43[200] + src43[201] + src43[202] + src43[203] + src43[204] + src43[205] + src43[206] + src43[207] + src43[208] + src43[209] + src43[210] + src43[211] + src43[212] + src43[213] + src43[214] + src43[215] + src43[216] + src43[217] + src43[218] + src43[219] + src43[220] + src43[221] + src43[222] + src43[223] + src43[224] + src43[225] + src43[226] + src43[227] + src43[228] + src43[229] + src43[230] + src43[231] + src43[232] + src43[233] + src43[234] + src43[235] + src43[236] + src43[237] + src43[238] + src43[239] + src43[240] + src43[241] + src43[242] + src43[243] + src43[244] + src43[245] + src43[246] + src43[247] + src43[248] + src43[249] + src43[250] + src43[251] + src43[252] + src43[253] + src43[254] + src43[255])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127] + src44[128] + src44[129] + src44[130] + src44[131] + src44[132] + src44[133] + src44[134] + src44[135] + src44[136] + src44[137] + src44[138] + src44[139] + src44[140] + src44[141] + src44[142] + src44[143] + src44[144] + src44[145] + src44[146] + src44[147] + src44[148] + src44[149] + src44[150] + src44[151] + src44[152] + src44[153] + src44[154] + src44[155] + src44[156] + src44[157] + src44[158] + src44[159] + src44[160] + src44[161] + src44[162] + src44[163] + src44[164] + src44[165] + src44[166] + src44[167] + src44[168] + src44[169] + src44[170] + src44[171] + src44[172] + src44[173] + src44[174] + src44[175] + src44[176] + src44[177] + src44[178] + src44[179] + src44[180] + src44[181] + src44[182] + src44[183] + src44[184] + src44[185] + src44[186] + src44[187] + src44[188] + src44[189] + src44[190] + src44[191] + src44[192] + src44[193] + src44[194] + src44[195] + src44[196] + src44[197] + src44[198] + src44[199] + src44[200] + src44[201] + src44[202] + src44[203] + src44[204] + src44[205] + src44[206] + src44[207] + src44[208] + src44[209] + src44[210] + src44[211] + src44[212] + src44[213] + src44[214] + src44[215] + src44[216] + src44[217] + src44[218] + src44[219] + src44[220] + src44[221] + src44[222] + src44[223] + src44[224] + src44[225] + src44[226] + src44[227] + src44[228] + src44[229] + src44[230] + src44[231] + src44[232] + src44[233] + src44[234] + src44[235] + src44[236] + src44[237] + src44[238] + src44[239] + src44[240] + src44[241] + src44[242] + src44[243] + src44[244] + src44[245] + src44[246] + src44[247] + src44[248] + src44[249] + src44[250] + src44[251] + src44[252] + src44[253] + src44[254] + src44[255])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127] + src45[128] + src45[129] + src45[130] + src45[131] + src45[132] + src45[133] + src45[134] + src45[135] + src45[136] + src45[137] + src45[138] + src45[139] + src45[140] + src45[141] + src45[142] + src45[143] + src45[144] + src45[145] + src45[146] + src45[147] + src45[148] + src45[149] + src45[150] + src45[151] + src45[152] + src45[153] + src45[154] + src45[155] + src45[156] + src45[157] + src45[158] + src45[159] + src45[160] + src45[161] + src45[162] + src45[163] + src45[164] + src45[165] + src45[166] + src45[167] + src45[168] + src45[169] + src45[170] + src45[171] + src45[172] + src45[173] + src45[174] + src45[175] + src45[176] + src45[177] + src45[178] + src45[179] + src45[180] + src45[181] + src45[182] + src45[183] + src45[184] + src45[185] + src45[186] + src45[187] + src45[188] + src45[189] + src45[190] + src45[191] + src45[192] + src45[193] + src45[194] + src45[195] + src45[196] + src45[197] + src45[198] + src45[199] + src45[200] + src45[201] + src45[202] + src45[203] + src45[204] + src45[205] + src45[206] + src45[207] + src45[208] + src45[209] + src45[210] + src45[211] + src45[212] + src45[213] + src45[214] + src45[215] + src45[216] + src45[217] + src45[218] + src45[219] + src45[220] + src45[221] + src45[222] + src45[223] + src45[224] + src45[225] + src45[226] + src45[227] + src45[228] + src45[229] + src45[230] + src45[231] + src45[232] + src45[233] + src45[234] + src45[235] + src45[236] + src45[237] + src45[238] + src45[239] + src45[240] + src45[241] + src45[242] + src45[243] + src45[244] + src45[245] + src45[246] + src45[247] + src45[248] + src45[249] + src45[250] + src45[251] + src45[252] + src45[253] + src45[254] + src45[255])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127] + src46[128] + src46[129] + src46[130] + src46[131] + src46[132] + src46[133] + src46[134] + src46[135] + src46[136] + src46[137] + src46[138] + src46[139] + src46[140] + src46[141] + src46[142] + src46[143] + src46[144] + src46[145] + src46[146] + src46[147] + src46[148] + src46[149] + src46[150] + src46[151] + src46[152] + src46[153] + src46[154] + src46[155] + src46[156] + src46[157] + src46[158] + src46[159] + src46[160] + src46[161] + src46[162] + src46[163] + src46[164] + src46[165] + src46[166] + src46[167] + src46[168] + src46[169] + src46[170] + src46[171] + src46[172] + src46[173] + src46[174] + src46[175] + src46[176] + src46[177] + src46[178] + src46[179] + src46[180] + src46[181] + src46[182] + src46[183] + src46[184] + src46[185] + src46[186] + src46[187] + src46[188] + src46[189] + src46[190] + src46[191] + src46[192] + src46[193] + src46[194] + src46[195] + src46[196] + src46[197] + src46[198] + src46[199] + src46[200] + src46[201] + src46[202] + src46[203] + src46[204] + src46[205] + src46[206] + src46[207] + src46[208] + src46[209] + src46[210] + src46[211] + src46[212] + src46[213] + src46[214] + src46[215] + src46[216] + src46[217] + src46[218] + src46[219] + src46[220] + src46[221] + src46[222] + src46[223] + src46[224] + src46[225] + src46[226] + src46[227] + src46[228] + src46[229] + src46[230] + src46[231] + src46[232] + src46[233] + src46[234] + src46[235] + src46[236] + src46[237] + src46[238] + src46[239] + src46[240] + src46[241] + src46[242] + src46[243] + src46[244] + src46[245] + src46[246] + src46[247] + src46[248] + src46[249] + src46[250] + src46[251] + src46[252] + src46[253] + src46[254] + src46[255])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127] + src47[128] + src47[129] + src47[130] + src47[131] + src47[132] + src47[133] + src47[134] + src47[135] + src47[136] + src47[137] + src47[138] + src47[139] + src47[140] + src47[141] + src47[142] + src47[143] + src47[144] + src47[145] + src47[146] + src47[147] + src47[148] + src47[149] + src47[150] + src47[151] + src47[152] + src47[153] + src47[154] + src47[155] + src47[156] + src47[157] + src47[158] + src47[159] + src47[160] + src47[161] + src47[162] + src47[163] + src47[164] + src47[165] + src47[166] + src47[167] + src47[168] + src47[169] + src47[170] + src47[171] + src47[172] + src47[173] + src47[174] + src47[175] + src47[176] + src47[177] + src47[178] + src47[179] + src47[180] + src47[181] + src47[182] + src47[183] + src47[184] + src47[185] + src47[186] + src47[187] + src47[188] + src47[189] + src47[190] + src47[191] + src47[192] + src47[193] + src47[194] + src47[195] + src47[196] + src47[197] + src47[198] + src47[199] + src47[200] + src47[201] + src47[202] + src47[203] + src47[204] + src47[205] + src47[206] + src47[207] + src47[208] + src47[209] + src47[210] + src47[211] + src47[212] + src47[213] + src47[214] + src47[215] + src47[216] + src47[217] + src47[218] + src47[219] + src47[220] + src47[221] + src47[222] + src47[223] + src47[224] + src47[225] + src47[226] + src47[227] + src47[228] + src47[229] + src47[230] + src47[231] + src47[232] + src47[233] + src47[234] + src47[235] + src47[236] + src47[237] + src47[238] + src47[239] + src47[240] + src47[241] + src47[242] + src47[243] + src47[244] + src47[245] + src47[246] + src47[247] + src47[248] + src47[249] + src47[250] + src47[251] + src47[252] + src47[253] + src47[254] + src47[255])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127] + src48[128] + src48[129] + src48[130] + src48[131] + src48[132] + src48[133] + src48[134] + src48[135] + src48[136] + src48[137] + src48[138] + src48[139] + src48[140] + src48[141] + src48[142] + src48[143] + src48[144] + src48[145] + src48[146] + src48[147] + src48[148] + src48[149] + src48[150] + src48[151] + src48[152] + src48[153] + src48[154] + src48[155] + src48[156] + src48[157] + src48[158] + src48[159] + src48[160] + src48[161] + src48[162] + src48[163] + src48[164] + src48[165] + src48[166] + src48[167] + src48[168] + src48[169] + src48[170] + src48[171] + src48[172] + src48[173] + src48[174] + src48[175] + src48[176] + src48[177] + src48[178] + src48[179] + src48[180] + src48[181] + src48[182] + src48[183] + src48[184] + src48[185] + src48[186] + src48[187] + src48[188] + src48[189] + src48[190] + src48[191] + src48[192] + src48[193] + src48[194] + src48[195] + src48[196] + src48[197] + src48[198] + src48[199] + src48[200] + src48[201] + src48[202] + src48[203] + src48[204] + src48[205] + src48[206] + src48[207] + src48[208] + src48[209] + src48[210] + src48[211] + src48[212] + src48[213] + src48[214] + src48[215] + src48[216] + src48[217] + src48[218] + src48[219] + src48[220] + src48[221] + src48[222] + src48[223] + src48[224] + src48[225] + src48[226] + src48[227] + src48[228] + src48[229] + src48[230] + src48[231] + src48[232] + src48[233] + src48[234] + src48[235] + src48[236] + src48[237] + src48[238] + src48[239] + src48[240] + src48[241] + src48[242] + src48[243] + src48[244] + src48[245] + src48[246] + src48[247] + src48[248] + src48[249] + src48[250] + src48[251] + src48[252] + src48[253] + src48[254] + src48[255])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127] + src49[128] + src49[129] + src49[130] + src49[131] + src49[132] + src49[133] + src49[134] + src49[135] + src49[136] + src49[137] + src49[138] + src49[139] + src49[140] + src49[141] + src49[142] + src49[143] + src49[144] + src49[145] + src49[146] + src49[147] + src49[148] + src49[149] + src49[150] + src49[151] + src49[152] + src49[153] + src49[154] + src49[155] + src49[156] + src49[157] + src49[158] + src49[159] + src49[160] + src49[161] + src49[162] + src49[163] + src49[164] + src49[165] + src49[166] + src49[167] + src49[168] + src49[169] + src49[170] + src49[171] + src49[172] + src49[173] + src49[174] + src49[175] + src49[176] + src49[177] + src49[178] + src49[179] + src49[180] + src49[181] + src49[182] + src49[183] + src49[184] + src49[185] + src49[186] + src49[187] + src49[188] + src49[189] + src49[190] + src49[191] + src49[192] + src49[193] + src49[194] + src49[195] + src49[196] + src49[197] + src49[198] + src49[199] + src49[200] + src49[201] + src49[202] + src49[203] + src49[204] + src49[205] + src49[206] + src49[207] + src49[208] + src49[209] + src49[210] + src49[211] + src49[212] + src49[213] + src49[214] + src49[215] + src49[216] + src49[217] + src49[218] + src49[219] + src49[220] + src49[221] + src49[222] + src49[223] + src49[224] + src49[225] + src49[226] + src49[227] + src49[228] + src49[229] + src49[230] + src49[231] + src49[232] + src49[233] + src49[234] + src49[235] + src49[236] + src49[237] + src49[238] + src49[239] + src49[240] + src49[241] + src49[242] + src49[243] + src49[244] + src49[245] + src49[246] + src49[247] + src49[248] + src49[249] + src49[250] + src49[251] + src49[252] + src49[253] + src49[254] + src49[255])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127] + src50[128] + src50[129] + src50[130] + src50[131] + src50[132] + src50[133] + src50[134] + src50[135] + src50[136] + src50[137] + src50[138] + src50[139] + src50[140] + src50[141] + src50[142] + src50[143] + src50[144] + src50[145] + src50[146] + src50[147] + src50[148] + src50[149] + src50[150] + src50[151] + src50[152] + src50[153] + src50[154] + src50[155] + src50[156] + src50[157] + src50[158] + src50[159] + src50[160] + src50[161] + src50[162] + src50[163] + src50[164] + src50[165] + src50[166] + src50[167] + src50[168] + src50[169] + src50[170] + src50[171] + src50[172] + src50[173] + src50[174] + src50[175] + src50[176] + src50[177] + src50[178] + src50[179] + src50[180] + src50[181] + src50[182] + src50[183] + src50[184] + src50[185] + src50[186] + src50[187] + src50[188] + src50[189] + src50[190] + src50[191] + src50[192] + src50[193] + src50[194] + src50[195] + src50[196] + src50[197] + src50[198] + src50[199] + src50[200] + src50[201] + src50[202] + src50[203] + src50[204] + src50[205] + src50[206] + src50[207] + src50[208] + src50[209] + src50[210] + src50[211] + src50[212] + src50[213] + src50[214] + src50[215] + src50[216] + src50[217] + src50[218] + src50[219] + src50[220] + src50[221] + src50[222] + src50[223] + src50[224] + src50[225] + src50[226] + src50[227] + src50[228] + src50[229] + src50[230] + src50[231] + src50[232] + src50[233] + src50[234] + src50[235] + src50[236] + src50[237] + src50[238] + src50[239] + src50[240] + src50[241] + src50[242] + src50[243] + src50[244] + src50[245] + src50[246] + src50[247] + src50[248] + src50[249] + src50[250] + src50[251] + src50[252] + src50[253] + src50[254] + src50[255])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127] + src51[128] + src51[129] + src51[130] + src51[131] + src51[132] + src51[133] + src51[134] + src51[135] + src51[136] + src51[137] + src51[138] + src51[139] + src51[140] + src51[141] + src51[142] + src51[143] + src51[144] + src51[145] + src51[146] + src51[147] + src51[148] + src51[149] + src51[150] + src51[151] + src51[152] + src51[153] + src51[154] + src51[155] + src51[156] + src51[157] + src51[158] + src51[159] + src51[160] + src51[161] + src51[162] + src51[163] + src51[164] + src51[165] + src51[166] + src51[167] + src51[168] + src51[169] + src51[170] + src51[171] + src51[172] + src51[173] + src51[174] + src51[175] + src51[176] + src51[177] + src51[178] + src51[179] + src51[180] + src51[181] + src51[182] + src51[183] + src51[184] + src51[185] + src51[186] + src51[187] + src51[188] + src51[189] + src51[190] + src51[191] + src51[192] + src51[193] + src51[194] + src51[195] + src51[196] + src51[197] + src51[198] + src51[199] + src51[200] + src51[201] + src51[202] + src51[203] + src51[204] + src51[205] + src51[206] + src51[207] + src51[208] + src51[209] + src51[210] + src51[211] + src51[212] + src51[213] + src51[214] + src51[215] + src51[216] + src51[217] + src51[218] + src51[219] + src51[220] + src51[221] + src51[222] + src51[223] + src51[224] + src51[225] + src51[226] + src51[227] + src51[228] + src51[229] + src51[230] + src51[231] + src51[232] + src51[233] + src51[234] + src51[235] + src51[236] + src51[237] + src51[238] + src51[239] + src51[240] + src51[241] + src51[242] + src51[243] + src51[244] + src51[245] + src51[246] + src51[247] + src51[248] + src51[249] + src51[250] + src51[251] + src51[252] + src51[253] + src51[254] + src51[255])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127] + src52[128] + src52[129] + src52[130] + src52[131] + src52[132] + src52[133] + src52[134] + src52[135] + src52[136] + src52[137] + src52[138] + src52[139] + src52[140] + src52[141] + src52[142] + src52[143] + src52[144] + src52[145] + src52[146] + src52[147] + src52[148] + src52[149] + src52[150] + src52[151] + src52[152] + src52[153] + src52[154] + src52[155] + src52[156] + src52[157] + src52[158] + src52[159] + src52[160] + src52[161] + src52[162] + src52[163] + src52[164] + src52[165] + src52[166] + src52[167] + src52[168] + src52[169] + src52[170] + src52[171] + src52[172] + src52[173] + src52[174] + src52[175] + src52[176] + src52[177] + src52[178] + src52[179] + src52[180] + src52[181] + src52[182] + src52[183] + src52[184] + src52[185] + src52[186] + src52[187] + src52[188] + src52[189] + src52[190] + src52[191] + src52[192] + src52[193] + src52[194] + src52[195] + src52[196] + src52[197] + src52[198] + src52[199] + src52[200] + src52[201] + src52[202] + src52[203] + src52[204] + src52[205] + src52[206] + src52[207] + src52[208] + src52[209] + src52[210] + src52[211] + src52[212] + src52[213] + src52[214] + src52[215] + src52[216] + src52[217] + src52[218] + src52[219] + src52[220] + src52[221] + src52[222] + src52[223] + src52[224] + src52[225] + src52[226] + src52[227] + src52[228] + src52[229] + src52[230] + src52[231] + src52[232] + src52[233] + src52[234] + src52[235] + src52[236] + src52[237] + src52[238] + src52[239] + src52[240] + src52[241] + src52[242] + src52[243] + src52[244] + src52[245] + src52[246] + src52[247] + src52[248] + src52[249] + src52[250] + src52[251] + src52[252] + src52[253] + src52[254] + src52[255])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127] + src53[128] + src53[129] + src53[130] + src53[131] + src53[132] + src53[133] + src53[134] + src53[135] + src53[136] + src53[137] + src53[138] + src53[139] + src53[140] + src53[141] + src53[142] + src53[143] + src53[144] + src53[145] + src53[146] + src53[147] + src53[148] + src53[149] + src53[150] + src53[151] + src53[152] + src53[153] + src53[154] + src53[155] + src53[156] + src53[157] + src53[158] + src53[159] + src53[160] + src53[161] + src53[162] + src53[163] + src53[164] + src53[165] + src53[166] + src53[167] + src53[168] + src53[169] + src53[170] + src53[171] + src53[172] + src53[173] + src53[174] + src53[175] + src53[176] + src53[177] + src53[178] + src53[179] + src53[180] + src53[181] + src53[182] + src53[183] + src53[184] + src53[185] + src53[186] + src53[187] + src53[188] + src53[189] + src53[190] + src53[191] + src53[192] + src53[193] + src53[194] + src53[195] + src53[196] + src53[197] + src53[198] + src53[199] + src53[200] + src53[201] + src53[202] + src53[203] + src53[204] + src53[205] + src53[206] + src53[207] + src53[208] + src53[209] + src53[210] + src53[211] + src53[212] + src53[213] + src53[214] + src53[215] + src53[216] + src53[217] + src53[218] + src53[219] + src53[220] + src53[221] + src53[222] + src53[223] + src53[224] + src53[225] + src53[226] + src53[227] + src53[228] + src53[229] + src53[230] + src53[231] + src53[232] + src53[233] + src53[234] + src53[235] + src53[236] + src53[237] + src53[238] + src53[239] + src53[240] + src53[241] + src53[242] + src53[243] + src53[244] + src53[245] + src53[246] + src53[247] + src53[248] + src53[249] + src53[250] + src53[251] + src53[252] + src53[253] + src53[254] + src53[255])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127] + src54[128] + src54[129] + src54[130] + src54[131] + src54[132] + src54[133] + src54[134] + src54[135] + src54[136] + src54[137] + src54[138] + src54[139] + src54[140] + src54[141] + src54[142] + src54[143] + src54[144] + src54[145] + src54[146] + src54[147] + src54[148] + src54[149] + src54[150] + src54[151] + src54[152] + src54[153] + src54[154] + src54[155] + src54[156] + src54[157] + src54[158] + src54[159] + src54[160] + src54[161] + src54[162] + src54[163] + src54[164] + src54[165] + src54[166] + src54[167] + src54[168] + src54[169] + src54[170] + src54[171] + src54[172] + src54[173] + src54[174] + src54[175] + src54[176] + src54[177] + src54[178] + src54[179] + src54[180] + src54[181] + src54[182] + src54[183] + src54[184] + src54[185] + src54[186] + src54[187] + src54[188] + src54[189] + src54[190] + src54[191] + src54[192] + src54[193] + src54[194] + src54[195] + src54[196] + src54[197] + src54[198] + src54[199] + src54[200] + src54[201] + src54[202] + src54[203] + src54[204] + src54[205] + src54[206] + src54[207] + src54[208] + src54[209] + src54[210] + src54[211] + src54[212] + src54[213] + src54[214] + src54[215] + src54[216] + src54[217] + src54[218] + src54[219] + src54[220] + src54[221] + src54[222] + src54[223] + src54[224] + src54[225] + src54[226] + src54[227] + src54[228] + src54[229] + src54[230] + src54[231] + src54[232] + src54[233] + src54[234] + src54[235] + src54[236] + src54[237] + src54[238] + src54[239] + src54[240] + src54[241] + src54[242] + src54[243] + src54[244] + src54[245] + src54[246] + src54[247] + src54[248] + src54[249] + src54[250] + src54[251] + src54[252] + src54[253] + src54[254] + src54[255])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127] + src55[128] + src55[129] + src55[130] + src55[131] + src55[132] + src55[133] + src55[134] + src55[135] + src55[136] + src55[137] + src55[138] + src55[139] + src55[140] + src55[141] + src55[142] + src55[143] + src55[144] + src55[145] + src55[146] + src55[147] + src55[148] + src55[149] + src55[150] + src55[151] + src55[152] + src55[153] + src55[154] + src55[155] + src55[156] + src55[157] + src55[158] + src55[159] + src55[160] + src55[161] + src55[162] + src55[163] + src55[164] + src55[165] + src55[166] + src55[167] + src55[168] + src55[169] + src55[170] + src55[171] + src55[172] + src55[173] + src55[174] + src55[175] + src55[176] + src55[177] + src55[178] + src55[179] + src55[180] + src55[181] + src55[182] + src55[183] + src55[184] + src55[185] + src55[186] + src55[187] + src55[188] + src55[189] + src55[190] + src55[191] + src55[192] + src55[193] + src55[194] + src55[195] + src55[196] + src55[197] + src55[198] + src55[199] + src55[200] + src55[201] + src55[202] + src55[203] + src55[204] + src55[205] + src55[206] + src55[207] + src55[208] + src55[209] + src55[210] + src55[211] + src55[212] + src55[213] + src55[214] + src55[215] + src55[216] + src55[217] + src55[218] + src55[219] + src55[220] + src55[221] + src55[222] + src55[223] + src55[224] + src55[225] + src55[226] + src55[227] + src55[228] + src55[229] + src55[230] + src55[231] + src55[232] + src55[233] + src55[234] + src55[235] + src55[236] + src55[237] + src55[238] + src55[239] + src55[240] + src55[241] + src55[242] + src55[243] + src55[244] + src55[245] + src55[246] + src55[247] + src55[248] + src55[249] + src55[250] + src55[251] + src55[252] + src55[253] + src55[254] + src55[255])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127] + src56[128] + src56[129] + src56[130] + src56[131] + src56[132] + src56[133] + src56[134] + src56[135] + src56[136] + src56[137] + src56[138] + src56[139] + src56[140] + src56[141] + src56[142] + src56[143] + src56[144] + src56[145] + src56[146] + src56[147] + src56[148] + src56[149] + src56[150] + src56[151] + src56[152] + src56[153] + src56[154] + src56[155] + src56[156] + src56[157] + src56[158] + src56[159] + src56[160] + src56[161] + src56[162] + src56[163] + src56[164] + src56[165] + src56[166] + src56[167] + src56[168] + src56[169] + src56[170] + src56[171] + src56[172] + src56[173] + src56[174] + src56[175] + src56[176] + src56[177] + src56[178] + src56[179] + src56[180] + src56[181] + src56[182] + src56[183] + src56[184] + src56[185] + src56[186] + src56[187] + src56[188] + src56[189] + src56[190] + src56[191] + src56[192] + src56[193] + src56[194] + src56[195] + src56[196] + src56[197] + src56[198] + src56[199] + src56[200] + src56[201] + src56[202] + src56[203] + src56[204] + src56[205] + src56[206] + src56[207] + src56[208] + src56[209] + src56[210] + src56[211] + src56[212] + src56[213] + src56[214] + src56[215] + src56[216] + src56[217] + src56[218] + src56[219] + src56[220] + src56[221] + src56[222] + src56[223] + src56[224] + src56[225] + src56[226] + src56[227] + src56[228] + src56[229] + src56[230] + src56[231] + src56[232] + src56[233] + src56[234] + src56[235] + src56[236] + src56[237] + src56[238] + src56[239] + src56[240] + src56[241] + src56[242] + src56[243] + src56[244] + src56[245] + src56[246] + src56[247] + src56[248] + src56[249] + src56[250] + src56[251] + src56[252] + src56[253] + src56[254] + src56[255])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127] + src57[128] + src57[129] + src57[130] + src57[131] + src57[132] + src57[133] + src57[134] + src57[135] + src57[136] + src57[137] + src57[138] + src57[139] + src57[140] + src57[141] + src57[142] + src57[143] + src57[144] + src57[145] + src57[146] + src57[147] + src57[148] + src57[149] + src57[150] + src57[151] + src57[152] + src57[153] + src57[154] + src57[155] + src57[156] + src57[157] + src57[158] + src57[159] + src57[160] + src57[161] + src57[162] + src57[163] + src57[164] + src57[165] + src57[166] + src57[167] + src57[168] + src57[169] + src57[170] + src57[171] + src57[172] + src57[173] + src57[174] + src57[175] + src57[176] + src57[177] + src57[178] + src57[179] + src57[180] + src57[181] + src57[182] + src57[183] + src57[184] + src57[185] + src57[186] + src57[187] + src57[188] + src57[189] + src57[190] + src57[191] + src57[192] + src57[193] + src57[194] + src57[195] + src57[196] + src57[197] + src57[198] + src57[199] + src57[200] + src57[201] + src57[202] + src57[203] + src57[204] + src57[205] + src57[206] + src57[207] + src57[208] + src57[209] + src57[210] + src57[211] + src57[212] + src57[213] + src57[214] + src57[215] + src57[216] + src57[217] + src57[218] + src57[219] + src57[220] + src57[221] + src57[222] + src57[223] + src57[224] + src57[225] + src57[226] + src57[227] + src57[228] + src57[229] + src57[230] + src57[231] + src57[232] + src57[233] + src57[234] + src57[235] + src57[236] + src57[237] + src57[238] + src57[239] + src57[240] + src57[241] + src57[242] + src57[243] + src57[244] + src57[245] + src57[246] + src57[247] + src57[248] + src57[249] + src57[250] + src57[251] + src57[252] + src57[253] + src57[254] + src57[255])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127] + src58[128] + src58[129] + src58[130] + src58[131] + src58[132] + src58[133] + src58[134] + src58[135] + src58[136] + src58[137] + src58[138] + src58[139] + src58[140] + src58[141] + src58[142] + src58[143] + src58[144] + src58[145] + src58[146] + src58[147] + src58[148] + src58[149] + src58[150] + src58[151] + src58[152] + src58[153] + src58[154] + src58[155] + src58[156] + src58[157] + src58[158] + src58[159] + src58[160] + src58[161] + src58[162] + src58[163] + src58[164] + src58[165] + src58[166] + src58[167] + src58[168] + src58[169] + src58[170] + src58[171] + src58[172] + src58[173] + src58[174] + src58[175] + src58[176] + src58[177] + src58[178] + src58[179] + src58[180] + src58[181] + src58[182] + src58[183] + src58[184] + src58[185] + src58[186] + src58[187] + src58[188] + src58[189] + src58[190] + src58[191] + src58[192] + src58[193] + src58[194] + src58[195] + src58[196] + src58[197] + src58[198] + src58[199] + src58[200] + src58[201] + src58[202] + src58[203] + src58[204] + src58[205] + src58[206] + src58[207] + src58[208] + src58[209] + src58[210] + src58[211] + src58[212] + src58[213] + src58[214] + src58[215] + src58[216] + src58[217] + src58[218] + src58[219] + src58[220] + src58[221] + src58[222] + src58[223] + src58[224] + src58[225] + src58[226] + src58[227] + src58[228] + src58[229] + src58[230] + src58[231] + src58[232] + src58[233] + src58[234] + src58[235] + src58[236] + src58[237] + src58[238] + src58[239] + src58[240] + src58[241] + src58[242] + src58[243] + src58[244] + src58[245] + src58[246] + src58[247] + src58[248] + src58[249] + src58[250] + src58[251] + src58[252] + src58[253] + src58[254] + src58[255])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127] + src59[128] + src59[129] + src59[130] + src59[131] + src59[132] + src59[133] + src59[134] + src59[135] + src59[136] + src59[137] + src59[138] + src59[139] + src59[140] + src59[141] + src59[142] + src59[143] + src59[144] + src59[145] + src59[146] + src59[147] + src59[148] + src59[149] + src59[150] + src59[151] + src59[152] + src59[153] + src59[154] + src59[155] + src59[156] + src59[157] + src59[158] + src59[159] + src59[160] + src59[161] + src59[162] + src59[163] + src59[164] + src59[165] + src59[166] + src59[167] + src59[168] + src59[169] + src59[170] + src59[171] + src59[172] + src59[173] + src59[174] + src59[175] + src59[176] + src59[177] + src59[178] + src59[179] + src59[180] + src59[181] + src59[182] + src59[183] + src59[184] + src59[185] + src59[186] + src59[187] + src59[188] + src59[189] + src59[190] + src59[191] + src59[192] + src59[193] + src59[194] + src59[195] + src59[196] + src59[197] + src59[198] + src59[199] + src59[200] + src59[201] + src59[202] + src59[203] + src59[204] + src59[205] + src59[206] + src59[207] + src59[208] + src59[209] + src59[210] + src59[211] + src59[212] + src59[213] + src59[214] + src59[215] + src59[216] + src59[217] + src59[218] + src59[219] + src59[220] + src59[221] + src59[222] + src59[223] + src59[224] + src59[225] + src59[226] + src59[227] + src59[228] + src59[229] + src59[230] + src59[231] + src59[232] + src59[233] + src59[234] + src59[235] + src59[236] + src59[237] + src59[238] + src59[239] + src59[240] + src59[241] + src59[242] + src59[243] + src59[244] + src59[245] + src59[246] + src59[247] + src59[248] + src59[249] + src59[250] + src59[251] + src59[252] + src59[253] + src59[254] + src59[255])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127] + src60[128] + src60[129] + src60[130] + src60[131] + src60[132] + src60[133] + src60[134] + src60[135] + src60[136] + src60[137] + src60[138] + src60[139] + src60[140] + src60[141] + src60[142] + src60[143] + src60[144] + src60[145] + src60[146] + src60[147] + src60[148] + src60[149] + src60[150] + src60[151] + src60[152] + src60[153] + src60[154] + src60[155] + src60[156] + src60[157] + src60[158] + src60[159] + src60[160] + src60[161] + src60[162] + src60[163] + src60[164] + src60[165] + src60[166] + src60[167] + src60[168] + src60[169] + src60[170] + src60[171] + src60[172] + src60[173] + src60[174] + src60[175] + src60[176] + src60[177] + src60[178] + src60[179] + src60[180] + src60[181] + src60[182] + src60[183] + src60[184] + src60[185] + src60[186] + src60[187] + src60[188] + src60[189] + src60[190] + src60[191] + src60[192] + src60[193] + src60[194] + src60[195] + src60[196] + src60[197] + src60[198] + src60[199] + src60[200] + src60[201] + src60[202] + src60[203] + src60[204] + src60[205] + src60[206] + src60[207] + src60[208] + src60[209] + src60[210] + src60[211] + src60[212] + src60[213] + src60[214] + src60[215] + src60[216] + src60[217] + src60[218] + src60[219] + src60[220] + src60[221] + src60[222] + src60[223] + src60[224] + src60[225] + src60[226] + src60[227] + src60[228] + src60[229] + src60[230] + src60[231] + src60[232] + src60[233] + src60[234] + src60[235] + src60[236] + src60[237] + src60[238] + src60[239] + src60[240] + src60[241] + src60[242] + src60[243] + src60[244] + src60[245] + src60[246] + src60[247] + src60[248] + src60[249] + src60[250] + src60[251] + src60[252] + src60[253] + src60[254] + src60[255])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127] + src61[128] + src61[129] + src61[130] + src61[131] + src61[132] + src61[133] + src61[134] + src61[135] + src61[136] + src61[137] + src61[138] + src61[139] + src61[140] + src61[141] + src61[142] + src61[143] + src61[144] + src61[145] + src61[146] + src61[147] + src61[148] + src61[149] + src61[150] + src61[151] + src61[152] + src61[153] + src61[154] + src61[155] + src61[156] + src61[157] + src61[158] + src61[159] + src61[160] + src61[161] + src61[162] + src61[163] + src61[164] + src61[165] + src61[166] + src61[167] + src61[168] + src61[169] + src61[170] + src61[171] + src61[172] + src61[173] + src61[174] + src61[175] + src61[176] + src61[177] + src61[178] + src61[179] + src61[180] + src61[181] + src61[182] + src61[183] + src61[184] + src61[185] + src61[186] + src61[187] + src61[188] + src61[189] + src61[190] + src61[191] + src61[192] + src61[193] + src61[194] + src61[195] + src61[196] + src61[197] + src61[198] + src61[199] + src61[200] + src61[201] + src61[202] + src61[203] + src61[204] + src61[205] + src61[206] + src61[207] + src61[208] + src61[209] + src61[210] + src61[211] + src61[212] + src61[213] + src61[214] + src61[215] + src61[216] + src61[217] + src61[218] + src61[219] + src61[220] + src61[221] + src61[222] + src61[223] + src61[224] + src61[225] + src61[226] + src61[227] + src61[228] + src61[229] + src61[230] + src61[231] + src61[232] + src61[233] + src61[234] + src61[235] + src61[236] + src61[237] + src61[238] + src61[239] + src61[240] + src61[241] + src61[242] + src61[243] + src61[244] + src61[245] + src61[246] + src61[247] + src61[248] + src61[249] + src61[250] + src61[251] + src61[252] + src61[253] + src61[254] + src61[255])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127] + src62[128] + src62[129] + src62[130] + src62[131] + src62[132] + src62[133] + src62[134] + src62[135] + src62[136] + src62[137] + src62[138] + src62[139] + src62[140] + src62[141] + src62[142] + src62[143] + src62[144] + src62[145] + src62[146] + src62[147] + src62[148] + src62[149] + src62[150] + src62[151] + src62[152] + src62[153] + src62[154] + src62[155] + src62[156] + src62[157] + src62[158] + src62[159] + src62[160] + src62[161] + src62[162] + src62[163] + src62[164] + src62[165] + src62[166] + src62[167] + src62[168] + src62[169] + src62[170] + src62[171] + src62[172] + src62[173] + src62[174] + src62[175] + src62[176] + src62[177] + src62[178] + src62[179] + src62[180] + src62[181] + src62[182] + src62[183] + src62[184] + src62[185] + src62[186] + src62[187] + src62[188] + src62[189] + src62[190] + src62[191] + src62[192] + src62[193] + src62[194] + src62[195] + src62[196] + src62[197] + src62[198] + src62[199] + src62[200] + src62[201] + src62[202] + src62[203] + src62[204] + src62[205] + src62[206] + src62[207] + src62[208] + src62[209] + src62[210] + src62[211] + src62[212] + src62[213] + src62[214] + src62[215] + src62[216] + src62[217] + src62[218] + src62[219] + src62[220] + src62[221] + src62[222] + src62[223] + src62[224] + src62[225] + src62[226] + src62[227] + src62[228] + src62[229] + src62[230] + src62[231] + src62[232] + src62[233] + src62[234] + src62[235] + src62[236] + src62[237] + src62[238] + src62[239] + src62[240] + src62[241] + src62[242] + src62[243] + src62[244] + src62[245] + src62[246] + src62[247] + src62[248] + src62[249] + src62[250] + src62[251] + src62[252] + src62[253] + src62[254] + src62[255])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127] + src63[128] + src63[129] + src63[130] + src63[131] + src63[132] + src63[133] + src63[134] + src63[135] + src63[136] + src63[137] + src63[138] + src63[139] + src63[140] + src63[141] + src63[142] + src63[143] + src63[144] + src63[145] + src63[146] + src63[147] + src63[148] + src63[149] + src63[150] + src63[151] + src63[152] + src63[153] + src63[154] + src63[155] + src63[156] + src63[157] + src63[158] + src63[159] + src63[160] + src63[161] + src63[162] + src63[163] + src63[164] + src63[165] + src63[166] + src63[167] + src63[168] + src63[169] + src63[170] + src63[171] + src63[172] + src63[173] + src63[174] + src63[175] + src63[176] + src63[177] + src63[178] + src63[179] + src63[180] + src63[181] + src63[182] + src63[183] + src63[184] + src63[185] + src63[186] + src63[187] + src63[188] + src63[189] + src63[190] + src63[191] + src63[192] + src63[193] + src63[194] + src63[195] + src63[196] + src63[197] + src63[198] + src63[199] + src63[200] + src63[201] + src63[202] + src63[203] + src63[204] + src63[205] + src63[206] + src63[207] + src63[208] + src63[209] + src63[210] + src63[211] + src63[212] + src63[213] + src63[214] + src63[215] + src63[216] + src63[217] + src63[218] + src63[219] + src63[220] + src63[221] + src63[222] + src63[223] + src63[224] + src63[225] + src63[226] + src63[227] + src63[228] + src63[229] + src63[230] + src63[231] + src63[232] + src63[233] + src63[234] + src63[235] + src63[236] + src63[237] + src63[238] + src63[239] + src63[240] + src63[241] + src63[242] + src63[243] + src63[244] + src63[245] + src63[246] + src63[247] + src63[248] + src63[249] + src63[250] + src63[251] + src63[252] + src63[253] + src63[254] + src63[255])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70) + ((dst71[0])<<71);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he09f35413664c4236c77a820d5851eb33ab4cb9ac4409d6a4ea393a9acc6f1eb5fa3e9a6860090284a1e31afb4506419c5ada3459624020a54827ba850f0d89d930306ee07550c0c2b8fe15b2099adc9a698e539dd18ba94735caaaec22c594d532bb31f8e1be9d7dc400cd173a9db83a587c05341f1a1cb91be2a39723de1337295dbd34168efb3740e49b14b47378c26b9059eb57ac332d9055022c8fd3b8f659fccc489a514492c2074e1a08163a29de88533a84fd469ee6cbdee1905adf50e40099ca1663a0664ad11730b906719bd053816aa2128bbd8727f4934c8d0d779c52ce8f0ca1cac71c33f8f0ec27fa4f4da8185b94ad433693311fc16a8cd3eb7f0a249b3a50a2798a4fc7ed1ab181647e05989ddd7205ed2efaf0c5c36d7ce9d1ef424a10af4c4eee86ebcd5b4a3eac33551664ffcc9709ebdb55e81af12f5d02bfea21b0176dba2afea882b84b69736b3e9b839dbba86e6d7abd372a556efee59cdcb80cea8888c4bc62f915bac96cc795fdd3506fece0a46d09f58d17a58f9214e57b2c0699105bef91d315eac93129d079df1db410088dabb97e5dd68c5aa57aa5ea1da1647d303d9540779259be2ffe7feec166db0b8c55b36823cee5ce73b9bcafb5205c7964492a994c6f366de3676809b22bbd28c2a84dd38c867c4e3d1d8a478dcad94f047bcb4fd1572bfaf0039edde44e6b73efcd5f192a55fb55c9013e9afca38cb3dc3fdc90e299a9a7f0dd349ee9b795e2fc49620dee8657d4ca990166fd8c7a4aa022e210f52b34aadb79599268ad816af3d2f085df9c5ff8ad160d56f5437c2fe996a78eb74239f3bacd46562b4e969800394bf6383199195b174653509fa21965432420cd67a793bae052b73ca8ca0b49e778e54aa1649d17dd2a2a06387e91b49077f589b8ae71e87ab7a862a326db58c812fa7531412ef4d954bb37573dcf0a73517de3e671bd60f4671b88332d486afc58e8623d60eb91981cb78d494a9a66f35378c027fde2a461a1abbe9b69aa5ec3faabe51e7e55dd137be95a140d3483f06ec7a2cdaeb31cd705a9fe1ec112f4336e982e6eb3c7e0ddb7544304467df367a842737bc118f129447788556d83744178ccff1bc9d7be9617397fc2ba38eebc29fd9ea012d4e4045e6041c1c18537461a156a072d98e5ce4748f91aaa4e616a32bedb789fe45e9cd19bf224064e9b4706d158abf60132c814934137cc0636cfd983e5614f24aad9f27ece9fb513ed2a6bb2acd48776bd5a34e11dab7f98cb1bbaf373577eeed3f8a64ec6c02fbddb5a8b9aa42c555bb0bfb856fb62d710920ba30c15e78c6f5477aafe7266688f1c4286077a4017a4142bd379ac5e3be77c8a63db2c921e3d1d70697c797335658bb0005fce7d4e4091f195259b35ca76daf41eaf35fa0725da2c552713527bfaeb3373abde4502f61e6262eee0fe09de08e65e8739358b4afeb7cdfac3449864621ad2855e12e9894c3919576077f446cfa68219cb465a1c399948e78720867be9292a9ccf55e467ba524dc6f57ae969b5643fd4cdfcefc76a31136b585fb90672d5af54f22530408bebfe6f5a0e12412663e2739b8628a3312f8ccbc837c89c7fa88a2f59976f342b8724abb691a3636c008307d8d415b4a498ac15071a1804ba05e8835412d369812d28d446fd5df908cfa1755ec09a2b2fc1cea07637d9bb317e32e0338a20b7a1d2af8a22f107df0605697e8194d4164ea15da2d64f30004c9e282be5aeb35790b3d68520b0b02ff50164d8e5c1ba35573dfa3805ed3bcb0d2d380b6dab7ef11f516c90b60ed11f9b583ce53abac90c6f3f5c8c51dec394a49fff2c69aa2e8a64a08ea10a4f986fe26b5b4f4f851d8ea3c5f6f2cbb4cb923db95c01efa8275757921184b2e4891c58fd1b7911c0735998287b58dea9164ea40a2c071729a3c8e46f5d3a889ad1c0be89689840ad06441fcf6e74d67306996588671bf646b514c54d119f9cb0ad50bcea8a9612167fe14ed44d8f3f708ec85e8ca8884ff2bc927755255e7ab85d1d0b76db9e5d0aaa8f440baaa5862324437591ae54bfbeef9ed3bbd50eed4a24a7f6ad606a40e53ea26cc32825841a57ade1f5caa561fd62b6f58327c2aac85e37e2f08034eced66c4361ddc6b6ca7a45cd9a7381ef3c90e5d0be1cb3732f0538772139ed02211178386da538a45fad1a2e6a0861bb989f642638547e51db6c5b260150240bac4d29cc08e33bfa9bbf184761bc6e3dc6952e9800fc4403748cf88f1ca3e1fc6a7d75f626a26a3fd6bca435f7547cde9ab2a6784114fe60221d5a68f0b5384116ec4e71cd015729425ee7645583e5f420e9b6f5798183d3ed9b81cc6fda43628a814ae05569934908705817132c95f4e16fe3a83deb33357b5ed02531df7d5d09f908fbc32ff1815af5eee0a643cdb7f1270bd85773cf56e0f4e1b37f544b88d245dc42d10c01103e0d35e1cb45f4bb964150ae421c00d39eb125f823b64351f097118d7181da7308a8c300e63474bd2de2de0f3cd5349236037203826219423fa8a6a59b72845bba9367e647500a142c8cb96b5c43fc28f33d28a05fc063a6f70567b79c638d445ab9ba3fde4721c8296ed6768858625e49ab5a55919aadb0068813f401c2f01fcfced44927973f828ed8f9940566fa00ed9504dd8b5d6dc2c124cd52d87d47e0a7e0a0e3569deea80515219bffbe2d5f5d68355e9de4f3c45f1643e841c90afdc5a94f0dd7ed7bbe94ace7c066dcb82b17b5867c6982ff5b198367e62f39f1fd29967dd06cd6327da1950df2fc7d989dd3461080b1a81495391fa0be19ac842a1f62482a8f1d1fab1baac67ce039afd54b37c61d71f41c417d05c8f1584f4fc530327190e58a814550638c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hed43e86d3a374c1d4b1694ae539ec01b489cfa8093a4989d9c134f10d24a4b8ab184031ddd7e213628f9ce7c893cbdb2bf6ce3f02965c4f2ff9314e65156cb47452df82955ea5d2ec8aa9e6b0eebb58e8e132667d33f89e2f761d4186def9573980d32907d10a80363efcff87f9e775e8cb6f598707acd4954d8f5497bc321cff1e908a1afe0b2f72cb5fd472449057840a704a2e6c823736c0e0059793ad1c6a4eb7661ee0ada1bcebcaeb7b75ebd32632644bdd0b9b8d97178b3f6d9ea477c4a12d8d2343400d0040794e1c90114c00d33a56d776551aa70f75a327875243044b297c052b883e9d2c077eb2094caaed5692b0f06040404fba60c96bbc0caac3699353712ad071cbad724a5d160e542fd94074972b5c77963857c1f221fe11c166a37934c403042f51b926058d51cfb931631e7930659602e16e31e9c01f64b011b292e42165e15ff902edcfeffc92e2d70462459ae07eb90ba4815586f31b84df968bab41c13bb49aa3102fa8cc19922851c1e819793495ce1647259745489407ff6acd0b12d4c708f76be517a8845694b8768f32f44a4f0d524993596d09dafce3374ec981690df6edea81cfbf15574830f6fe9636c211ad5c099d477a27faaac8870f8a582b274c1caa5bd9474eac2c6c3cbe4884437d1b91245ec9c094851787b27376e2efc8de00d034ec670b75ba82a4f9cc1441d8cf38d31236a9adc8b69ac7b4180434009bc1ff220f4a3d4e7e4b2ec913754689173d66b0576b10a935f8e9bcdb5882d84f6ac6943c9ebd1610a725a7f27a46750043c8751c8cff46ffc0dd6f39c8dd19a9308914fbd22fd5fbad6de47421112f096ea2ee132c89c61366527cbd30e97b426c7f0a87e4c2ee9ce1b2c9ea2a6eb6f8dc7fcb9dc09672db01341b50c479320a40e2e421608b0561173b2747df2a4bad7db1c84ea4295ecdb093e0a7d9644325fedb2e176f7923a6e3aa50ff43f9e70137582755ba03d07333f6cca396f1de354974a5af2e2a748b5fa707c3c97d8af8f45a4e83430127fa2896017d8572643d3cc48c04a931c0e0b890e6b72f5f8ad42534d4db925f7cd4d59867e2858f1e63a43904bd97571176ada1c30bd49dbb087c2c27afb88dbe400434439605ba5e9f50f8df54cbd22adc3ccd8a0710eb1f2eba7e4b7f5bd8a882796b2eb3702d91ca63a865c63a8728be6858a1339d71f5441df51a4cf84b5c8141668525199bc6a5637cdb2f9d1dc51744079e18b46e9a317b515441184b4386453d7f4d9cd780515a6cdc43e044ebcba4138b19dfc8d13d28acd7c7897260de0d6964968132728ed7ef20f29405e7f1f976c3b15bf239588508b9f2f82a4b61c60c2827aef4e75f31519a6d25869e2cb34fa3523b1ae92cce0037794e77736a8f9204baf66ff174ecd5ca31bdd9c40fbce3e699619c0a0a1b7ddea859201a21125adcd44fb28a2aa5323959be5ed6d3f0766447c8134083cbdd670502f159f5bb9784dec3061ac72079479af8069da9a9314c14a80dc81da3e182bf7fe53662046761e1f803c1f4464839c62068f26ab0af4523d5bc311d71f150a8963ccd69364c22181fe6e27da5f0129afcfc27a28e599058f200161b46c46f968aff8be191c59587bd368be9db5141dd582bb35a6cc902f1556cd0b53a2f87f1dd101533fdb4c9623b845bb3d3c401e3d8f49f24b1c378a2a1d3d8ef085780cf63e07e461419ea3e44284d446c7854832cb8cb8a1ae7c454a1477a9eed56129e92acab8751d7ff1c20d695bdcdc4a8a69d4b5aa7a6abc417e856dc408364d7b88a2ab668ed1ed7b8010b2f0d582272f417136383d49e32a286453dd8f12416c9c9b8fcd6eb5c256f726864bb66c2cc0cf0572ffabb9c4703688206729ebfac950cfeace1cafdf292294aa5a0785f9f421ad267e4814da85612c5950db3ce46251de84d7841edffc097fe83376f1a7a8bdd98577c5f947c2b7f50e3998d09910855ea1fc2e1903bf63f8d043ed103a3077769608ec044e259479078978e86b9f752a25feff423424476f38af240c8ca6d10e26c003b1c4f2569cc65df3503ba952c15cc856d6a6d806f4e3e0f50c474155be503b54f679731e723db793647c90ddfea8e11f29d24eedc2cadcbcfc21457a19178f9740394da5a81f78b4aeb59ead794ffe238bc436e9ae9b6439e7622c9557dda0a0c5e554eb53b58692d40a0141bb43dd1e904e12b5ed46c9f89d4110453620c6b05847c828555ca9857ade01a5e70642b7d5ac2b99a549305bb928dcd57b6c4491fd617ab43665e55893770db11d565507aee60374bb9aaa97bda5d69730b6395182a46c8dd28fe134aa8c8f26e5c410663b68cbf0f6641454e3be3b3b7bc5b80d763ded2db3988be0a283cedb23e88e187cc53d5faad75dd8630a0dc4beb78e9d29fdc8eb5757264d4a2d90ab1d9d7501fb15497a36e365edbaa4603103a584a35daf6dc6ebb7ef4b768204e92b6ee524bfd83b151cfdc64cac37405bc62e2d830ef221f2c71563eca3f1525cee335b2eb0693f63da09248050f804f8651e759c66027c6cb1c527387890b335ca2e9be15114d7cee4f7df6467797a19c09c54eb81ca633dac369772a867b3b7ae183a56fa6b1d02762534436eae76659238772d547a02564f83977e4b0bbc40b0b4a9d781102ff8222ad383c09e53d8ccf1fa697889d72eb51a7a0886a92d1eebc538501210f5312c2279fc8c2fc79a3c8e08b03b7e55210d7ea746ea842cba9eddc2bf16a9a25db928e034bbd7d924c3ab23afca4ee82ff3de87152b7795014812070df3f35d4fc6e323c5e368c108e42401ebb035e5f5433cfc539d581f7c19f5079e2f2dcac803e1382ab1cf1869725097b1b404b994e21a40ac96e0a8785f8c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6d7c0852ca04ec0efeef8cc20a01402e08392b100ffda593e03b79ad0f708dc094b963402e08d5fdd29e81f24f2cd9e2c6dba6af47e80bfcb0d7da559cdfb1d1bf9f7b86882297b8188c10ea1b0d28a24fe0449bde34656f00ca91ae7f8aa04583332b0afed9f4c0b18bc6020483304257e806f4116585db3e179f81cd11000ef3258eabf4a7e2daa69328d98a4560f0dcaabfebcf7452a6a4a252e47a3f96368af9e023ab05990508acca9e0997ef81c78ab84855d7d752e7c3204b02a8969d4c72dd4232eda5214e3b334d60868fe5fb63b24e13d15885f284af4acdb9da4aff8575f5f456b8240c0b528707e64be1a8119fdd23726ac7e393cdb069eb94857be1ce4dc0170052858f764dfdf12c20d84959a8cf91a4fdcdd084ad21bce7be7bd4b77d8b3a287843808ffa737159b62566e8e1b700ab301b81c4e75afbaaecc4420412d92a805c27e660869f791e1303ac4348946aace5fc2eac10ad521cba1a19ea68ea303d6516ec6e16e37e2d9905db859c9d25798e6ade450b5611aac53aa634cf277fb888b3f6769c009d6a16aaefefcdbf698c812cacd1d019eb905ac13bdb6f535123d294adb4f523e7efa48834c9e804365824e671d9b90b477ae3a0f8147e3a49563a24275d00a9b7b0f24180aecfbc6a0374aeca38800d8ace49296c89135c61878853fadff1a99474251ef998a21f53962e5d297c4a9ea6a0a51f735b2e4abbeba171b5eeccdd299088a5fb61b189eb8b0a3ae00f7781b16c7bbd109cd66db9c20ba8df8dbe2e473324b91d28157edd737aab4ed3b78a33a340039a36c7ac00bf083cf308e3ff64483db8473acaab4ea9b80086d35a68960a284b11e40fb1166717112d9ddac9895a15e3f2817e17fd7a4b107554e866edff00dd5acb8933e34577cbfcf4a093e32fca3d41c933914b649f7f20d93c78551aae7d3d84652d7c45b11bb58217cf7018a6f4572261140f6eae7b1707777e74575d8f7be6f4c02b6527d63f7b9f9ad3d6b9f0bff8d1bed0433df73cef3a60926810e55846a05b46dc562288f307106062e0f794da1e157700a1f10d85b303417032305d372d6bf013af3c5335a7ed00c314df3f363ae96e1b796ed33d38b59314dd8891f60fdf7f513694dbd9a9d6432f278991b8d7093d7cec2e3524e78852406b13cc9dcfa53aab2b3a88eeed0b36a9fb1d5e59e1edf84de7995bd98095c126d09d217b213ac1e7a326871c5950e0e3e413401da39f7adc6457081632201b34dad3eb11244dea5eb5ec71429bd38c2a47c82460fc21eca93f9345d90f8cc37103219ab83b1e90297875f50ecfb5096519bab7799d9ccf9042e37de32fd9d949113c75a950086045c234fe27d79550464bd90c0b0e9689714610844ccf755d0a80d53d2a184da44ec48425465f0cf64303ece5b8335c7fea523fe90caec79ba5c7e11979d19af7b1afd0d49a9fc3f43d9afa095c0580e9b3e5004b1bbfcf0fef8ed377a42ef3e42ea4ee9dec148336b03bbfa0a251e639aa3450dca5048595323f8f4d6a8fb841596c38d8c08e153786af028e788bd203b40a566bf7acb0c106f5c45eef180212ac50e9e82db87362906447c27bea82906ef1a902a62099ab0764507d30b48ab6a57bed908bc91e4a0de9a61f294f4e11f9c2b5edfe4be4875a387fcb9b07b394081afa47975c0f63cfb2f463c1995623bf9ab3d25b0a614a59df05f9f4aad631484447d0d534fb42e0af10a37b199209caed1f8062666247b67102e3e722bddeac5791a50cbab37a4e7a4124a984ac91cad1f9fe57d7c4569fbde13e5ac244ede577e66aafde8e85329da25220041bcd606a6bb89ec3cb6ecb482253683282938b58e09d32e4666a185454e3957d174c6f0969797751ca35417fd9be7ebeb37cccf00bc381f15765d2748a774a82ccad155daad7487e121867304ef4ccdde8c4e9526dbdcc7a95230a19cd863367a867c1f4785d78aa55880846603bcd208eee793fc23142caf405ee2ff0b0178512f3d6374572cbd6f529a7544fdc1f89d7b6d1edd585b9b0be2eff5ab56152c2f506ae6c213eed402e25955c42538211baa08c67d87fffbfc9ab448d9446a4424cc044f3ac14c98a6657d1d0955c1b285d7b1b66fa43d0431006c75eb63239ab4197e59104ec4f12ed2470ed66c28a8304d079f5e5230035a5e9c9ab2bb9212c082d98034bbceff41ec3f28c0d9492ab4186c01b9df4d1e349266ddb696edf352974eecbc51131a4ce937555db2dda268bcd584968ca9a521a1d1384e76ba723d44d42b08ed8e6da7faccd0264fe46a360d8cf628a55e3ff0fd48d8cb5c30af804a52d289cd8cd1a35f3507f19cad80edbe5ffc8fc1c3d6ca0ac91b151fc4a24a37cc5d5e477bd145e4f9b4fe4be48b4360c4d818d249b7279f54b345a8e7590f52ebce2d1515e45676967ca0c755cfcae6a0df4d985d3d479b6928e3a0cb9dafe7f3ac3cd8a9048dcb35707679ea2b55742175188a5bb63e7fdee5721a47c8e6462d738dc9b595d8288bc265b90e42269308eac8e254a3c945bfcaa2535aa7b0d2072b4c81dbbaecf77e934f977685015f8ba5853397147f9c7bfeaea04c92433654018d7e825bcd3a6d00182de3ae1b52113264bc1a4dbc85beb6ff523d89743a8ce0d01d2f8b277c74b95f55337c759a28a962a9d5bfcb83617ff5ce9cb323068760e1df21be1b1331d4a3428d4460cec9bb497369005b6aeb32cf5c70b3ffc812775a97c2fbd5e6b1de9e898912bbcd7077ca2a0e203604ed2b281191eacb5ac54d0f35638623a044d263a63e556efa99aeef7034825eee028bdd177e869594bbd013ad0242bb62ce93254cd336b6ccab0dd9b193eaf651832b0930ba25040e7fcf5cd37efc7d3fef9f9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h451946169411ff8763cd4204a490c395c98f432ef7e85db7580b2b6bd3f7ac67b56db4b3ccd0e61ca82be4fd8591794e0ecd88010f5b2459443620653c12407304a4e956625686993278faa8df53c7eba7ca4f153772047c13846dfbdc041fa0561f1a333ae95c3a35534489e55df205fe204a291c30d4c2851febf4f743510c5704981fdc56132e725b7be2207cbfc8a8316d125432f819228edee948a70d2fae0a0aedd2fb1494d23554af9c8ead247cf2759ab5b420e3b3924068a5c203426da97d0f99ae34c4962cf1fac9c5ca9043130fee203b4eca103c5d35b83e37beaab7c31f41ba49c6cb706ccd341e259d01a9146e85e928d61d9f48823d030f271c755e0419024c5b70a783fdc40a9ef29bc07c39b075dfd3f9bd0c63349093b9cbe6ab8e4005c7c5cf67373ba3e90d54261c0dfa630b60b967dd4794d56f97a0aaf81645c198af1e5aa9522f6d96d4c0f54200770e25510e9e7278d6c6b3d5dd824e531818c51943b79b426344c8ead02e2d62eb9e7ccab072d77ff61b28c6d0c850ca420ea55dabfec2927115b1a777899fa4a5a4e5728b25a3a58af544a2837b33a142dbbd09b3327bc6c1a3fcc0aab87d5cb5c7aec9bdff354493cc0f12e37c9bf0ea3396c7800a506c35eaa3df6176ba6913fed6e870655aca07178a82c100944d14c310918ac3187e50f7a881aedccbf8ab76badab64009c4cf4c8cd7b5ff6b975d53e3b3d301942b8a9158ba37723cb506c95c70fa16979faf7a08b06875ef2166e12459382d1f7fdee1245f8ec7666c5e956e913f62cc8c46d9b43679e8e69e393aff7b7c2d7749200acd71a2925bf8647adc64cd8d834f5a82afb28e3d47d9cb7ab61858ef30a0b1fe3c09af70d45add7e1b8c3dce0de46b0e6d9b5bea901d9cc385bd9741dfaa8daafb5171eb1fbe3343159ccc6a3186324d25cbf19c124747266452bbabdb594c2d7cc0dd8c84334b7701adb08147dd63b129f36bc0c5db24646001b3f3111afa8bcec6231272dd7854d0847cf6c953a15320d331459bb26bb343c90f64e3e9e8734368e10d20e13bc825b84701da0998979c0ae127358189e95ad128fe043c6fafc15820ec9421e45aaf50dff680e53cf84f9541a305916a079452426bb8246315fae540ae437916ce904714af66caff6ba6675638b602ca824c69048322773afb12f7be31bed68a255692761c242f67470d9f39f8bd7ec4b89ab16ddb501bb2925d8cd6372027889b31bcb35e8ed93dbab6e5d860e019402f8e8a3749ab319cd17cf4271016aab226f97b28749d93c30d834abe8cdaf6ec34f59eb9be5670c6754b323a73aa82ed360b1e0bf5bea79b81064f7ddc2880eacbaf02159fd86badcc8c362377ec5a073727030ff78e3523244509ca9791e85d0dc7313bcdc279a12db03e37f54654c44b39ccb6150342caa6cd4fd2b5cf8156fc5123f33b6328fc309111e83177a54bd6111f1f96bd95c673598450207721f5ab3aae7e616490505a17af0cad244755c5ecacff84ec81b7c0e6839a637bcc4cd44ab84545bc728b6cbf9d21e3e1515868e56ecfb162842b5609a73f87e534a65412a510384800add1da60512e302b8a685e84385c06143698cd251ec0f76e7764ba79333aacc4c3e3609c198cd14192bfafd71740cf8264778b402493f50029f49040793102ed84decd71de28787aa8e4fba8ca30df85740f289ccbf083be1cc08838641c798f35ef51a464f1e45892abf710d2345737236b93b6b0687607ddfb1201b45a97e001dd4c4fc7e38927d197e500ec4a301f67816d2b5ca362df88d9811d2d297ade150fbf6fb3529ebabd425deb4fac240905b62e04578feee409c4460a32aa7f541f8689ea1f648d8998138e9206ffcef185bf292f780c66d38ba64b6f5c456e96ed34d9c93d30a9af0e4be945226e0846bca7c4934c06388aecab5dd397c366b3752757ed7655bd52fd38a94cf1f31ca234bfaa1df651ab397dcdc03f1723895156db16ac47fbad855f688897da9109de9c4c5838c2027209b7e186675f8fdebfb7c8f298df390ebdb4eda8d087e2af40c14e7e36c793ea671896ff5f9915311695e8c5a24654d70433405cd5ccd0065fabfee78d6eb7acaf15055968ec207f319a2712dad13c46b8a76ae04c58c8c4dfd596f068381d3fad01e16856196a4fc9cd45c596d95f910ea667848187993f8dba7e4d739ddb1a48c135e6fbe7d5c8727371388eb75c5d3e3b4ae450e7a812351bae93e031300c3a82a8697bff74e37f1211aabb12bec314517bace30c2ef291436a53d4dad0130a04dd95476582a5fb766b79332d81d5aa27670525f0bbdbf33766d7448e20b0e4064d7c64fb52f7fe858b9e09efd04fdb280190ec1e6cdd54b6fca87f891557fd8fd40ed0e5320be262b92aa23b82bc13e36ffccba5ed71b01c111423156f52146e048ba853407aaf52c01c09ab02c7d8b16981d5a16e22be07c27f447ada7c16c9140479b79875bebc34168a0dd425e9ece6f0a4d42471981f94457269c8a04fbc9e4a8e4342782f661ee4c6f5d0ded8de963fbcba2fe17800670172cc68ab03a8b0cdba9e278d8b9d87b537fc9a4c7569fde9d7f59abbdca4f8256653d1b0d0da544825bf93f215aacac5258ddfa355ccc3ab8e1dd08a7b79ff88c091bff8ab31d1a9cde10547cc95660375cc5ae57ee48e4623cb5c05bc93303d08f54fa5adbbd83fe83e7a5252708ce54f04254d5500a51b66bcd1f7650fbdff394ce5f5ff4d6347e4a836ccdb85ea059c351d1f6cd0fc6b061e8dd79c85ec563ec327af4e093e5ea6cb84049acf289ef32873eeb5bcc4b23275ecd5179a0fe4400f1a0c2cfe7087b0e9d12700a66a0b0374d5205c530f588afd44ca3be65a8e433a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1bea4475212f0616c14c682b6e21a9e382c8143fe9091792fc74e45f46732a2e1bd580cf67551253cdf73e04cf90619bbecadcb5cf1b458c4bb12beaa952e864527bf706ff7a87575e346fdb47090e4c07afb061c44fbcdefdefe7ed00d5a2780f68b8d4378cf9018183406e1ff6e52310600d202d4d35e11c1d007241c54589c852a86c83de57d637fe87c2878ffe88077024af2cbe080afe6ee956fea91ae7e0a619349b3c3000b5e2f3bf75293c850b1aad613218862d9bdf9a442db945cd9fd90f5f01b4153399b78a62510e190a463c24323df9fdfc99bb2c32b54ea75ba134512575afbeee5ab46b8a7a4edc8a0a95212c634a60587019c4d024097e603ed8dac981de26cad91e2ab0b5f27a37243db05dacef35b40e1fc13ef1a028d793097d5ff57d8623635fc14e609d975ca29302bfa21041dfeb55f6e1d9c5c971b625e574dd528ba648e665dd65a5e73570e00adc1d02288e213d956fb862cd7527f866f9c9cc841d6135d273e410a19b58ce86cdc757f6a80717f707bd104d2c9b5dda7245b1c81baa869c03d421e0e57540f4f45f6a12e379a8102e0a075fb666b0211168316f338833840e7046a5201d2529fd3a38f0ffdd8f73194d2eca9b145faf67956feab60eb901cb1edf6fa5b675add40dffd6feafa0329bae3fb595ab87f7d1e927763120193d919b9fa88ebec901ebb51958fa499a6b40fddc301ffa646fb9c1f34ddcba35dde3ec5fed9f99de99e993f79fe10f7adc03f5ad3bf7469e238444079bad79232f2a59eaf72797c22f3211dc225b90afeaa4a5d056ef15b24804aff121695e2751019bb172e4d5d961646da11219aa3d88320009ad0262190968c6e634fe60662ca1c8766fdb1776423c7c9c7c874286b284f5c884c90d2eb2f7287bd7e801792b9f3eaa55cd1772a7cadef767ea13759295f3628253dd7c73bbf5b19ea5dba9a585edf470941a90ee7004769e58bad118716574bf833e6cb648df4f6d6e4e20a6a8e88fe5ca1690df58875e4b61706cbbd3fe27ad461a51f0e0e482f04a234934929304c4f0ca19225bdebc105cf716d66ce0eda2bcd1f401e610723119c96c2432cff758202efaf67cc293d7458fffae4144c8fae9fbda5214977c52be527602efbac16c2239d4a2efd74856325d1cd22e5899e9077487f4a87c2e7fc9074fe1bfccef6281b9f49c6c2e46e410f79d7531c66c1934c0e05485027c4fd502701aaeefd942183be01ad4a9506e6cd7c5fa7fe4f00ef5e9c4558a8a3eb9622cf2673a84d60e8d308428fa232c5a22882e169ae4b4bf352fdc29bc221a63643c085cb570a38dd835a44061cbde9ac7718f970f897f439dcc643e807b6bd20229addd0d214b28614726706f76139ee789ebf36829a05adb76366c696ddef1e1f0c22073052aae10593c31dc28618d7d752bcd4b1f4fa90b2c9e238d1961dbf76303870568a6fb1593003db8701c545a0a91728f759790219702c260875eb2f992fd3dbb3c5c51dbd453f56135825df4e7dec8f5f45b03a2e41ef4a7acf88f8b1f230d75b932f2be3e1a9fa042e328d3e2cbd79c3d745c87d8c3a4b85eb48c5010d9b459b1f793472562f8c331281565a406e0a3e81ca63d07f95db8f024c12c15ab8a605c833ebc8ffc666fd4f681280b3ac83158ad719646b23d7efd96b9f97fd4caf0a99c499e5ac2d4cc9d20c395b73c1b4362ee6302547facb18a850374dcbb7091f9caee158ba76fe5c6a2c9327d3ed90c6342b571ddef417fd6d8d9ecefe9b16be5b5010497eff50c7156a9fc3630975e946e975d1461b65765eff35a13367479c6fdf75fde1bfc66979827f44f3f8d080acd7b54c18bf94adfbdc31536120dd7facc3b3d2e9d66a76d6be612a37edf5e5b38c7001fed8309215dd6312d50c6cac4beac4528805b1b55ed503df53f7aab16d8569cb0ff4dc69215c0156f2a6f40c12847efd4d05668f048380c03b86438179afb755ad76c49b44207773137acefc7b802137da11fa5688b5e8edcb4b866dee223dbae41bd5340ee25d4e57d49f9e160bd81595f56d9a5fec0cd85403d2ca49af3335edcf86ad1475211cb13c36ca18374839269e77bb9785bbb4b09d2bfddcfc1e1c46ddcedbdb84b077034aec242488fcfee4af77ebf40938c2b23155faf61a3a915e880207580edef3dd482c444f5b6ee6d1f28e519fbca7cc437b42b7e7ecdc7c427bc07a1cca902a368ae055bb7d1e687dfa590ae195c05e6f239529f1e0760a9d2e7178eb69779603828f92b29c7fa1884b86ea08efc16e2857471c6c36f2ac40e546e5ec355e2626d14a35e8b0eb35a304d864e3225a125aa3f5da2325125e92046f5f7882c85d07b69f78d9f7f970a1034ab20889f80182bf6823c30adda5fbf01371ca5965d1100a2ad5a5eb2a59c2b7bd18b4ad6ceb9b2189607296d5b105c4944a9b4bd254a90cfd738858c5d1f40f43dc9a21e6e28f31e79f77e33cb9500e43ee0962585aa030347c0751e9eb15752be8707eb21cab67d343cdb827110302f17728fa2631ea01c73638ed097f31081e43dd6516bad576ce70a923c0fdf795f01c936659236baa09900a40021b876f00fec46a9591fb5e7f7470811a8baa3c0683bf598bcce0976f3aaeb6d587ea269bee8c272da900135708a2b1fc152d39d16a9906288997a60c8306fc1447eeb98b7b3d68ff80df1ffc4cce35122deae00dc12bf3f832bffe96db338050a64a51b81f27c28bc7aaf09dff9ce3261751f4835f616fb56195447a26b404ba59d7322fc46c867c507f008a404e18495330325d940f4d87eaead00dbc66982f9e07ee8238e92cde82a2ab589a15b408d66c289d554a46e4c499ad0ff5ab4caf707410991e8ccd0b8dc388eeadee80b02;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4fa1721d5d4bbfc84d9a31728c51b581b7912430bc2f2c3cf5e8b8b8d93342533e82e72085be04cf41d7fc4e955db20f97be18a4924f9164a77a51c87902f2908b70b06eff25dc60834889e582dd68a2ea5202a3734aca4704ffbf717b4ff3123a838b7a2bf32033a21547765ec1bfb871c9caf297f82920c3ae185825d1afd4b38021e302b279f85649e236789ccd136590c69e3ed215f3b9e0b5ed84957a7b93d3e42b3be63754d7d03380a8ca938a4f27e5676dbaadd52caf53e8bb24910e54693f407fd7e3cae4f46a904da692a76c061c222deb3b375e23a0517b7a4ef3399d1274302973592c2b3df70a2c3a53e269a8f83004103af608d7104543054e2486c1b968e2a22e673e5585aaf4627e13108fc113d1f918c7cf6d76b5048d6bce1706cb8c5b48ab90033d8b0182b2c86fcbca44109a16f3ba140df89ba53e0d85cbe0585f5df57634bdb65ecb0e1591d5a904e42ac5871c310c84179845eebc568dc0bd11ae68055b0113505e90a1c87f31005a4d48ee121a91190ac20bdb21fe7de8a3732e4faf0788995c67e018b2f138d434a9998b9e1fdf597a175ea0cf45486cc2ebf78bb3023b33fbf8e4c6009ec3ee071edd0d437c61a6240f59bc73b41a63eabbd536206535540b0f0a788c7531a3c5e8b926c5975423bdaef898acf4972588f4c599b0e5e56ffa56f2e63b6db3f5a734ea84f10a69fea9c7af17c141d6bc651ad70fdc9929ab08af214bfb8ec6e342cf2a8232b3b7c1e9f9d1014f2465047421a1e60eb2af01366e5ef42ee1245fd5b6638b0da765e048aefc349b15eb36627da021245d78ad04c1e684745337cb997d013e5a95283aa9be9c580e511fe10f64a00573b923d743f88dfd08dbe524f7eeea169b294b5c1aa6a4e8c2696d73823b6a7b7c89c6d0e70a4b002be4f5a23a238bc35829f952717dc1310ab9ff2aeb5a006a9b68648569deb03902214e53ccb0ab98a092f042ff391edecb8dd409eecdcbc7e3003fb1d5054086977c68a0cb46c71c3369c8b32acc341de1fd3c1eb17cdd658b1c03416e675c707ee46c76f8dca4be85041797ff392a8fc1811b38d0ed2ac3b1eb72d52cfb38d65701146aa216d995e21c4f98063e62862f27985df5a97038366d41c6399c804cbf3ab2070a4a855ae17cc17db7915037afda2ddf6d434dfe1cdee31ef4f11339fd08808829d01a98873ba6e35681d0f012c344fc8be7f5d20c2d9849ac944d92e920e0aa8c5b6ff4169956d0009c20fc3a2c6ac6c3a9c99bf96450feb53fb2d0a4955295269513ce683f7d27fc0643657ffb9e8d5972ea691c54c31ee68604b978afd010905c358ce702cff89eb9d7cc3512324e0f129f0a94b43cc3482ef139543cc9b32fe1f52493211943ca8331b8cc51ed09aa5950471c8b1b578943a1af9cbb8f772b7015976e6f595f88e9902cd59ea82e9a7b22d6d38fa14a17c6930f69ac2c2952d89d6a7e6c43482e34b484da201ab845abc7caa4df5394729cc83bf32a5770f123322a86f268f64131a8cc984df52fec2633ffb616d536eb000c87422d75e77f6069ab201acbc14e4f90d167a9750ee331e03a63d9ccfbb590983658c75a11001bbc2b6005f4b8011e5bf2ca79cc7ffcb84f85eb0754fe60415887a55c0dc9fada4672f250e4fce418289f9fb693b2b586882d5996d3480c143913a42989b978a189029a73a6473d2f65544f3eab946ec0358e5e839777386f4d3224af6805f84abc229a3da653f96b07183bba8943a16d2448351b9c65fa8832890443945da64d91cd4c762ee8177351c1b2c24c481a33b2b4c61d87a532964c3d12a048eca66ecee2c02080dcc28cb9f72b3b0a6b671e112441b8e7bca136e1e1c3c5aa9db385e9f8589288abbe0cb5cb03a1cd32b90a076de2247a4dee942438eb901aa23ee0a11e534b01a871ae9ba2ac3df3bd021d7a079b315e8e71eb2c3c6e44bbf2a360536f726215a673d7c2bf2048b0fa561f3e4831bcee5109ee2dde64a988e36a5c3dd8c1b08d4b35a1695a9a41531d75815a414856b746ae78fb6a13370dc73cd28a8d84bee94581780892366e876b50769f833f84fd84e905412f4109060a2896cda33cf9052d5be3aaac5575ef01ff8831b81a5f9571227380ac34485f4ca7a6b51e3ff3542aa0a690f6281770e3d20bcf89c1025719fdcdedb7ea36671f2c9f4bdb94a8a5a2c38154e60534dc9474b0153599b2f5737be06982997cde3e41879557d1307ac747ba5394fcd3b6137ac70abec587d9942d7d1d398dc23453c8ce983ddf0179904baec0c62d1631f9c01b1ae9567bfa4f58cce9bf327eb69b8feca45fae319dd6c93caf4b0aae56cf851a54391830afea8efc2bc893a5eba01d10018beecd571e66ccb4b7d560d5d9929290897e51f5c507f878eca5375b012c30b0be0eb39a25d48848eabc7d45f365507c566a3fecdbdd5c6b8715e20c4ba623a289c3b5d120d430214612aa6c5d6a3d217f074a58c7794687d61194e82bf843702bcb4148b41ccba271fc8070a1964a95c739ce27461f7ada3da65383694524f21064616f31a04f2a75be663931dea6e6908ebd7b6ddb963f998a6041d9ea409f22043a95955def3acf261690ecdc712555836e212b0e291c92666813baf7b06f976b9994ed37011591c0b30c749386e8fb10884ae40dd6c51f05aef948072ce4709e3ba827e05658dd8d15364dc3551fd0defb36e56c86073b8f7ac89ee355d85e2755375de91aba416a3f31306d27f0363ba0a61725e42c817f9eec182771b5e1f9e98bf99e800412c202becd4267595932fe27b455971406165222cf835fdae7ccf59dc3a19391c25e5fc8f6a86923f9ac049725276c8fb48efafca0c1e4aba6a2bf4a0154a13c8b7f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8943a562c224f293866329a7f26dabc8fb6b2fa875fc2f2a5ce8a90b4ba76c6ef42ec904152afa351e90079cd55b638d76e2aa21c1f08e0b27676290ccbd6a5a640b514b73850e23b62e78ac16db2a927fdb11b84010dfbd7dc67c630158103710833f692f17e90a24206cb3e776744df357647e24cb5d91ef807d84871445a4cb24c701bbbec2cf125dfb10d189218d169b854fc3bde788f139d99db4d5247fd71ec14b44fc54428a2ee2f35689bfe49798eca1a3a6fcd24ecefdbf9497b27bdcbbe6c594b1d6e77c6e062b417c7eddac8cf652fc73aea40f2f989a12918bcd8f0c5db7fe83c926ad9450f134c0512feca11268e1708d05bdf0db160463c0c2ea331db86b63e7bf91b61ce7d28a2099ef9a08ceb29ce8ef4e0f92e4215235770d6d6d2479b26b9657bd787e4abb9e32cffacc83db489dfe55430b1fb9b92d53c23315babae811d0d16616ce6d58353141b2d0fe2f5a301628309c1db587638fda86b6024e397236e25cc18d5fdffb546f53541cebcdadaf43821bf74b4b3cc7a27293a4ab555bbe3073bdfd84e57cfa56ac95e7efc07e62a2a0ba5cccc1f501b07c3b8e91412d04e0b63811cade50a3e1355be6ea1ff8e4b39cfdd001af303606ceb17bc0ebbc13116983f61355b432b5623b48440b81a19907837e72bc16efd3e9cb5b4ee0b84c0a3a11fcedec6448f2e55e22dce82bb8ffc506bf8cba1016e89385fc98749b17d06138c043cecc308d009789bdc07824fc657fa13815098ad3eb5961c402abcec2e98896e5fc5a21ab07e25d1d3de8236b5d998e9d0ca428e2ad633f671617af144224e304412bc93d0944cbff6e568967ddc18085980c17b465b4d8e6f0b06b21959f63b41228fc7497f892381d9ac5b827547bc26e9014d3ac1d9ba5a8c11bab3d6a64d9a65180e4bd010f761e2ab048de616e0d3a6f3fb40b461cd976905230dba84c5f120f5d65d739237d76787a75ddf6afa050cfb2cbe12325d5eab8ac8256e75bee1c05aceb90054f4c893a894361369532fa6744a0ff52e9c2bbeb5ce01c88ee0834d3dc057821cf26e211a7e312ebca4dbe08c2e910129a2bb0c6c03349a510c9adea616c56934710dc25ab8e221e130954340fcfdd33ed78f347bcc45aeba24778358a25658928d15ec5da76bb11afbd8516b2891a7e78694aa73860a750ebff0c01707bf72aaa850ba4cece2a34ffc93a6790e81df323e2457a8fd9beecc36b3fd88aed1299af91bf8cc8f94102eefbd31e00434c07f194693f2790732e6cf770e6a856db7ee86a527db2ded991a99f84d7b3497cf8c8cfa320ca43e2986031ae2a24b986e7394a35c364ab54655db2918e98f532ed60620233560837f7d9d2f1351ab14c9e13bc73de396cf77ae3fc4d0784adfb9119bb4ea232b61b166840f4c8a2d5eb1588009f471bf6f8d29336fff77be302caea23d4afdf2c0afd4db83a3516e3d6880215e55a94110d6b269099db5f063ceaf502cbd634c47dcd8abf61cb25dfaa59c63fd8769d0ffa7438d3d4d5c7dcd269a7de3e7cbd323d1405403b5680cba888b1138d85c9b73df12d1bab1f8ed16b630fc4eb86dc65c1764619032663456e8f17d6c8b3f77e626b998ffce62d09c5962ef0b74b5309f4f717a0ca43d87c487cbb529fdca0e739d2c51eadaa7afd92fa7e54da7832eb95cd4278364592564e00fc44c5fcb1fc8592891dc149af2387b32d493e5bd6bfad6d62c340b25c9fe5d0b55f616be91e5b7e70db01f046484b3d7326a7851330e5ee1e6e4f45e5fa54b4994ae4074e8cbcd1822ad394c47070faa4660a1cfe591997901f588dc1852bc5d2672fa873978290ea144752808d1f4f65c1b2a359194715618ff7e063d741800ccd7ce6a59f5455b3779408e3694fac57d21ea068d012966f860716e22d2fd4053d1aa5d77ed51864e62713510f2c2da84c77f19cb647daf8f7b9002cb0419c331aaddcca7d2652fc2580dde66c02ea159c3653e40b9cccb4d021814c0524b8479acc02a11ed6eca8d4ddd38b4acfec95f82a1099a5106aa45a201daf962ef4884a3053107941aed5aa329b96616d6ae814546153c68ebc6dfdd81bd18efdca0bfdfbbe5f89023b2ba9b27e52f5df98396ab728ea097e20697974890534d37f65d17111b93c27ea020b2d91a666f1018fd0e71642c900840e1056cbe54b4f537ca510d21246409ab1f1c020c8603a9c4a29a7775fb79cfeb4426eccad6d6ceb72aaf75a30e488822a20b9c93c9099c242f3d31ed8635f4294e76bc04d0512a3d20a09ba54a6d6a3478a2b3247ba3f1dd7fad20b63cd208062f13a10cd436d240ed22bf89b786f7d6899f84c7d83b9462e392965ef53b0fa624d8c2a25d94f9aea119eb61c32621e1457988d8f1518115ab9a7a4dcf4b213101dde099d3bace47e4642a6dc93f2b93fd89282f1cdcbd9665d043b2aed1b14afc0de85db2d37664c857934af9bc3805f9fd26c9a9eea0c688b12979fe30965594dbafca15562ec173a48c6c1611ab4f4a29948eb2e752639f26cd23be787eb7757658f4b14a40f8325dfc42f202725967f3eebeb25a9eba94b32befeab1c5eaa906534a338b2867813421661abd7ea02cd90f87d64141cb80b0403ac36510f06c3e506ae36abbcf26bda2930a19eeef78a1017bc9fd6d71d53251999f0e17a124945890d581f1beda6cae1202929d2895aea3de3cc2d501a947e946bdca6ff9f7340128cfe2eff78ddcbf1635382e313bfa6357a238bff966a649db351f30e3db6289e8264792a3f60bf105bc2e2c82f25731817f3c1e4eafbad3b5dd6ac1f71dae20dffa19b7bca03b290a2580b9970842bce1acbfd8f1085e5e72328c09a453883f45f3e2314a3f35548a87e7a1ae2d46ea3fe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h797e1ca55d2dc815f3c40b4ae7297bfdc1b26e07bd43d2e83b9b8a3077887ead8fbe88019afb772021a0bead9d0e605d51bcf22da817682e9c6a0344986defbc7e426ca97f2158fa429112872672d170bfd3b8964303e4701f82a7cdf113de2151dc20e6f0b88eb245b72602196b33a86121f3922a079fea75e9ebce89aa135c66d773a33d8088ff8709e63527acc773b72f410674f02839ec17b538bfe6bb9768eb09b0fb3b1c7b407950899d865fe45b1401a72b9c5aa0652b7ec6e632511fdbf72fe538d63240c6a868f717126bbbff3ceed8a2b6a1c621a6eb3146b2d655b56631e0b50dfbae98de834c059fa4c64267a538e72a247d09fc61c77264bd8a987c0db0b573c1963587c20a6f58a8793e930b5787eebaa6beda6217edc8481b924aa2e1f993d80ce952fd4b30948f76e938aaf044d3b5c21bfd2812fb819a018d50ed3173beb8e5dbbd9f0b4ade49bd5dd2342735937955aa4d43de5e8535cad360f26ccdb060bb37abd2f351365d4fdc9c91fbbd401c9526c3af0dd368a8f696a27a7a99bac4201ceedb51fb401aa9ec42e97dabee238d9f9d5e7d0c0f08eb4e539738d2446fff90ac38c0e79641e695381773039466271cef74230591fe54ef9846d1baea0113af930e55f2981a101065d90bec707674db5cf9f5594a71e90589cd241e5e496bb6c4383d004b6254070199f3c78ed6359f86d7f364b7d52fb98fd419873ed97fbed5dd6bb76aaf62b7a76ad3f3602a1bd3ae7282e609175926d56017a0bdd1379fa58dc042eb95c9eb2a7457c712533426253fb212ed2a36c397104977c7db103e5122c13b503c9259032f1e2d4d49b5a2c488203dea10be2a858d53f21cdc45b788e607bff2afd71733c3deb8efdc26a05566ece80bc3ffece00edb268153e9d363604adad188ea971dd9f100a919e8ec4056288a2e4e02c9d204022100acf689310c04b9a1d98624fbf872d7805523f36055625cc0c09a12d04891add5e51d53d7db8140b74fc59e20bc2bb23eebe5c6b864a0a1c630834b41acfe921f26e600d37585a9311b6eb113a83d054deb6b05c06c25b37ffff1d5cd9249d32ef53426ed9af06802fd7cb6ff71457b192a9d091fe5d50bc1c161c6ac27ce531ff101470d6b6216b5aaaae3a74e647a6cd5cf055a5c383ae8fcdecbc542a465ae7fdd4512790cd5223c9076476274edc7c735c51ded31b47a94a084d72b7650fd504f5b4e37179a9ac9babeea54ef05f60023e708426a3908150bf3004308d35a7c34955b7551af4af93aa5f88e07b03b73d169716376e81fceba0b3feb8dcf396d59c745920fd157f5add338a539774e1c8661f6a2d03c6dbc608430f537c1f374e6cdf4015276e3a3a6d0f82690424eb95c952ae3a3a342d897fa36b49c8a0ac88b397147da7fc2a73d98db56ad94bce04d65b150791a763851023b2483a7e51e03489058edeb4de529e5e952d990702b2125720d38e37dcd6270f6a8142e36b57de08fcc64edfd2c475ee95ff73049d02585b948c028bf974eb6bed65df2bde438d9f37147aba5470169b7a2d6b7e7e95556e033bf2ada7334a8ddc8e8e76d9bdaaaff4e5433855db4e016e49044939119b5d5fa13f37192892692c956964d16c9a71ed2876d0b64489f1ad15f87c5e67d12ed51360779174afbb2926409efcd864d79696b62e33cad6c9f617b515d8eea38071c2bcb36e2472dd5932bebf2d550c2b868c90b20e4aad85d03c27942965b37a2ecbd1db35517fea0725546802844fade691292086d72e3c9b1c13a9e807a607a489515a136a7f066ddbf694540943dc97f912a65f30b0d89fc4c72233634f90f1c0f50fb52b27299d300b7b3fb9d07847c86b944014ee7a3e8a0aa0e4eb32e7e025afe6449f217356624f9a604c4ab1add2c27d8125747b6933e47e2a211d22c672ac5da755cf8ff43ed54e63a34b825e6e8f398066fc4e8136f4a25778e4752b283daf11b8ae71f29bf8664346eedbd47d967987111d35b1078d5f5a6b57594ffb6eca626b0fc69c08a20bfd22fd0918b2d2243a45d50fc74ac643c829c93ceffb046dcbb5d723717f2ca2ca849a03fe81cae5fc0a442a4cf631228584aae4dd7896078beee6949c471ea750afe4a2bfbf812004d804e7e70a1f97709ccaa5e607f6b1a27dec8ddfa5d2d8caec5ab32420ddbf4497d1888b53bacfc54247d8f1d6d5b79462d59ca583e4fe2172d2380ec7c9806c6863dc1ab3d0f09f36079054bdc3f4c0484ef46368a0c7c3483ad958eada3617ebdd767edd84f40234bce318a5b80354cd2a826755f7b33e71f5e62caa9c6bf1ac453d0417409e651c56ccf5d9329803c0ae23e6ff1543e0b2d9388b44514951ccbc3b143bcc0bd0f8213bc56566b19e7381fa053f51e4b9fefd1e0b0f880fd26600049f25eec2d7b13943860d430b4a2734594688a6953033c0e68738c038200a3ef618e56e42e0e1f8daa750c1c0918c509834ba6349bd25545e6c95264fe0979d1f54accbb8464fd66690715bb5a4552f0c8b9232db5df2ba3f225c807648beb0fd90017c6c26efcd884b77ef09627e0ec7f52f838821c649583559ca1e6c3daaf94d41e8081ac0fd46bd0ab68bb082d39e0e14c25ae4317ab114ccfe48b53ca2fe5d1e93dcff5df7c40833a895863110c7f2172864c2f3409ff31f8a46d668dfe690bcd16e5baace4ae47265eeceb999eff8e8ee5d9ad6ba2dc86fc0e0d2bc5df181c319bcd0cea5ea93ebabd7d739b1c62c6ffa69c61506d384623dcadf777e932a323d21696ace5e853e8bb0caf5c0e4815405b54f21398b9a5b42ed2b74a2385b5c9c742037b570ad5d74e5ee18b7ddd156a7921041133b2880cc6502bd2a72c7cdf104333d963166fc2ba233a3d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h48020f64c4d337976ed187eb19484269100a40df2d0e16f14d9920838e01cd74d2c32a8d41494cfe2a0201bf79d61d3cb8424c12869569d478bc22d9f5795e7759b0a52d6cd5e8d3ba2fe118f21d8a106d3a4924db9c8b9cf20fb23af8e24abe91b5966d756ce23331574db6388d0ef48d86671836de90a6f53fd2139b7604c00159f2fcf2a4cf69093ee0486cfa3f246019d8bfe9c99ed037042a24662e5989bc6b806ef5978fa5a04ad04464904c49d322cf147c435220cc06474ec99afeda60cbb97635339d84db024cbc3fed3435a65c9d57c572e0eb3296e185d286e8b1e8981c5299d8f6cb4a4aec5cc0e57b3750739cb7287d8514f714a63f1ce0ded6ea0934e0b8fede11dac51d97c1e07dab8ffc011f80911d772439e8aee6004b959cc2737c8ae834c5632bea8fdb8a6322cd35137059864f035858e67afb8926a30a39b24505d695952c37564b075ae5d0fe5437b34de92fb7f0a6cd10c52c7b32d4d6c669946ac12fc3515036ad8c2a304ca150e239c7fce1b964cd21db08dadb54ad83adfe3bec0a2c8ff78ff7af5eb42e2586db0c5201dc1bee93a6826e0db88c59c6daf0d02e32533dd01e74cedc42068aa972be9a1fbb09e6702eb1c55bc872b33bb07546c877cec4f2352eedd243f29b1d2eac533f3d1c2004be4cde64c3e908cbc20295c43451b7f9074c03b119f6b79adf4f9e2ba1709bc63a8d6e68d84949306e22cfa6e330cc61ba7693f412f8c3e990208e53263174feba7d7a22b18493f0755b347c895ce2c5937f962b2f2920d1cb8d0bd9c646dc55e821a27c9bd5956fd0e6d91978554401df0492bd9f7532caf3bd19b3aae2bac6969053d12528491b5e1d6894c601c81b244b451b0c1fa75710b58e275c0d63620146ceeaa5bdb2b8ae26efb6d59cbf9b0809b2f9df4faf4304a7e36be4e519edd68924ae25843bcc63f72168e1475ec3a2a39dcb1a54ec5b838516835df32f2324e76a448cafa65bab3c2a92869529b7d740367b463812b961efef2851cd8f88382155796a983f7198a47d75384fb0a5b6cd211968ba7859f81821f42ee48bd650c05766cbc72c32f91647b2dcbfcd4e9de5d645dabb8c54aff2cc03fedcdf08e7a35ae7b73e2a503ddaf5a095c071ce7baa66f846abdfff5862711ae9ea844fc509496352cb1a52412087cbcecb658a4d93b1cc0b12da49b8c043f1cfe5127c1891b58e045f78ebea17f296bd2baf017905ba2756e1a7303033a96ceafe6c4f67bf2873cb3cb8f37bba32e964a935efe8127e313e87b2419ea452e610ac9f3088bf67b59c34a8fb0ae5dda09b562b85ca9b1f17ebec87cdd9cd221a9d93c1e88e011109803afe3324f842e23f49e4a2724b87dd29b4e3ed16cd81c807f904d88e221d960283b5f0ca5d0876e631adb6059e7d5ba2a89183a826c84149ad7a464c4d6eaa76ad57083d3a8216bb42c4ea9de688a99c70f979f80cd38d2c761e17e436b1fbb61cb77e6585dd1af4e9e1e289dc9a1913bc46367a72c38ed62449c9d75f6a05fd704239f55163879edf402722a9df300fdf36d3f2b385c1e5f6af9b015f092dcb387515055ff8dc0ceba01a9976ae4143adea188a02f12d8032afed372e7ed159ef73e3e97e4ff886b758d499d548b62463deeb8cae31dab15c30a5eb8aa0baf2c960d8ff24f438c547e758d94ac72dfaee62c8579ae0026a61822199097f01b3255e8024b7faf6a7b219cddbd5411338040fe0bd062a16988018f93f515aa5158c553166cca085a5456b2087030ab19edd09a3b69589a2bb5d55402c1f8a2471deee7368c20e69fd8a01fe33fcdbde871be16007486063deb40285cd26a97595987d543b107e77f0723ede8e483fd1313cadf93b331ba8bf2d33a14c8c9cea1575ffcaa50f83ec14376cfa04eb15480d05d8a9b4956eab3ba435394dbcff8774e07e7d42f9e0123244ab49b8b1ea29efbe0f1c0c9845ba13167fd844b3402fcddfb993542542c6770b543cbc74396b240c8d080e5f2fe9d6058e6e184260f7ef0718804c9a71f4acff96072d83968a808c7400ba234fbb30203969807a6cd5127061abba2fda266dd68c7b61544a8e6d56cece52e55f4bd635145683a3d71f270b6ed803e93c396612eb4e1c5eeec88c6a54ebde21036142cac05815009e4e7489e33a92968304d6e51ad4c253055e54180a0f9ce32e8595cc2cf47a46928e16951ba9aeb09bfd62c05e772d731ac3682139d46f7dfafced0f1b117b2bfc3bbb5b46bc6afd249ee53e014ac166aa0e92683ab0a13433162143c363dfe5b076e05f272e2f0d96c732d6bec6569fef4ea321fcfa12aaf3eaa232499c0ceb5408a077c5589d7fcc8de669f68cbd5fef955c8f8b09233040b4d1143bb23e85934edba52c7db769433f63b59653886dc99466f57febc3e9896af2b81599281b9e649384537b9992812cd4b316caa29048b9599d362c85c89793e27d204b8de0d900c0d7a0b937633a3ecc741b0f312176744fa8263b0eb7a0a8293a582a9f562e5aa1eac3fdb6b60de5db35b36f75812489bec540f54d04972d34c999c698cb60849654949fb1d4807b2643815e58fe86a8117c77792da62da6ebf268ae390418de87d253d50c25a0e17c23dd0739efa222182c7d0c2b36ef298c19474bebce52606143ad177e99587b4e62f73fdcba239b06e062c6794a00e66fe0077c752ae31cf0736a930726e7856bb7a9488736cde6f36629b92d960827d11fc4ea2e4b9d66a1cf8df1eb78060b073687e5db04e782fc73fd4804e0b8f2473cf881fa103a6015704e3fbc133c6d5cb4ea35dc8250cd4c30f7103eb65cc1d038dffa55758208361ac2613d2b4844fd58a6a224407b8b8150a7be2b09de1420a165b6d28db89299;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h88bed55d7e4708093885bf9a06c734d8acebcadd6cda487c1be778ce138351107748ee8fec940434a58869c19e50fb8d535a28f45589aa20d301c9dddc118c37170f14d8dab030b8ca57e3a09defeb80a65ca798e84f917b2b32f58ef05f83c4f4e676bfc719115139746dc42247320e65b5b5c4f0856351580983078213ded82d774cbda640279c4b5426754252ee2dbc27e776e64bdd4a5a6bd7282344648c94f4be381004ca268212cdce2455c89d2ed4e52ec0bcf88a14d61f5d46c0b0c08d880474c430d4e82405a7338c64aa776e591376fe97067f86a65de051f9698b5bea546cba056e6b9433d7e59b6ca2b3ad49442b76540249bc01379f0ac869ffd9870bdc7f23e4074858802fd92df311493535b74521bded1cbef2ceaf1c18c342e51b87427220fcbb7fd90a7976154be9068db6de809fc11a366f30c2f17ed41cd93df4b4dd903586c6a1dcc9c18a01c243dda40c0a14231e58b8c820f13c66095662e1ff458e9ab81c7ac434402e523e9662c2695ad2968757ee890bc0018ee3e9421c4805dff27ddbf8d9108054c3720f33961aa14c43bc30217d6e8d8bf359a1127792ec9d72e434ec0b4c0209b4f17b10a746ac04c9a9983a739fb0241889ee76247034ae4645f6bb27b4aca7d971ccafb09d28271189b5dbb63dcda3030487c22a2e081611446deda1d93e86bc2f97a386a52b3288aef2d887d33bc75cdf2ae87bed87e8924ced1bc19c301a7934c59250caedc26e34a90d63745d9fe823f0ffc580e2825b15eaae22004fe999e804059f121965f9d217e60b35847a6e637b36a1a6b893d9d07d370f9e64f40be01a068751632f1abfaaf423e0d09fab04f6782df05b681c5fd2415f7c94cf99868ebc502f4afa46729d5a56fefff46eb930312c0b4a24c3c1748358ee4d9ad7250e4efa42c3d0b691d5f2e3de7ae6fa380e4c12556f86df6b4a032cfe4de53d7021be9a3318bf24d5231095b2c7709f67d0aaacaea478d07384f18d984e6dac6046cfd91e9b548ea80d1064ca7f026097ea24b47139e8da2091e002642d7eca9cfd40efa5d2945bb1c6c18ca656a933c6520bd78d679bbd5c32d63cbd0a5eadf656a367439372d3ef7bf39047d05d97dadfbcbd26bd10412e6e2964de6c2094218c2ac1e83412b5bc8bc0d243b38df9c4ab35bc1cfed6e3e65284d94e9c833921b9bf88b5b6b5c03635ee3ee3b824f77534463af01663ca9a24a2f3b7e08f4c81c9a1aaf57489423ab14ed3492bb564d84a373f4bc696919962f337658e511c2d51ffc155bab763a41e36195a1c832da693ec6d360c56ba6086304233948f345c65bd59408de29b0c841496c0ee5dd86428f454570e044a2accfbca1556134c180c70a5c72ef87e360a0f01702df239315e366df7ea2fcb71337a7c7d05f0e796aaa3ae42dd45642ca6262ef05ec55e92c955c712784b9b9504bfcbea02c3fcf574e8f290bd533b0f26de50232d4eafa04857405ea23a1f08ac5d717cc3c462a1e10602ad654650fa7d277f3661dcf9c4c43c361c0787613799ee382bfa85d01e6c6c761714222c8700fd5b397ade949962f1d6a671e1d307ec0f1ad94b0082b9b5a82077b74140fb10aace5ac68c6b45a51602f9f4da5acf8962f806265a9eb448d9c8062a9da235932a0c7a11713c554ccf43201b7c7495db95794fd2e8759e57594e0cc60ac53a037acf10bf65702429f88d82d0f10ad9d97da0b637ebcc55fe5d368b3f0aab6a41b4fcb4cc2869055b4c4a3bd061d6693b64af6de8b2ed22116c2e889b91051f352b2604436eb0c53f6e37935d22f80305270fb63f395061c60845fa18245c45fffb952bfd1171fe1c1a363cfcc1237a2b9cc59d429deb041596dfcbf86df69568bf08fe2e7906ac4c7c533d9cdec154bb0d2b27ec1537df06dfd78dde1097503d2de065279e66b33afc4b037d85a393053f8433b5ae7a14bcc1c8f2db6e9fb0529e2521385a19395a131e7314b8a693ab31f95b6ce21fd2d99bc40f0ace58cbf54495aa8a411a5957aa9001b2a5b529e543492340f87c585a206aae2c9fa12055661dff35fefa074e9d15906678bfea24f7214064c375724f64df538e16dc66c54b696bfe78d3bab45ecb3a5caba6c85be43fb83d154538ededecaaaac0e45ed7553571fd986fa3057e1761e8a0d34b68243c2560b26ae2277f53e0c00512d7f7861a28a059c1d421f8895052d66f08cbb3da0c8769c3bbbb542d11b74682102aa265881b05ea430996f3ef21843326621c1adc61ba9996fb416e32308ec4469e9abbef74b81ea99c8d20ca582e3415297c02798262a7c3a8f755ba60486fe123d9f98080ed03c90d55720d3ca898faa5fb300f461b66a041f822ce92b5c4712a5dfb2a64d3f23ffcd1fa5be2b26ecee7beb87dce836bace3f7841547b82556732a0731d48acbc37176b81c0dd906837ca0715005f50d608d057b5085e8301ca87ad7570aac67478f4f94edbb29461e206eab7b686fcfc038235074dd17a92a3f3457e250d65370b4582c77edab4762c77420ccb3cae46e8e63d97305a1bfd116a670e22729d8b03e222fc0a2c29822dcc4746e6893fe3a07e466d1c60f40683b9219ed9c8676bc4f4ffd05fed01e16d7144a50b0dadf7018fc4f190d4b820b7a20a9daebe9a07e93dde867fdfce6082b9b3174919b4949f48e3681cc5f5f04b231c5543a3fe060eb2695e41b66538faae2185865169b3261de2962b27bf17f0b10b1b7e50278c3a7625e9df6bd0aa4e9b6554d549e80e075bf3fd0a3f3b5e0886f2e48dc1e52c829e475d80f4f8a3ce45607055d227f8a4e74feb8c376d9467cf39dcebc8d3a1fa74db872543268e79537385213568d4ffac41b889b144fcec1c3c7dd5fd649;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6121285e0fd85e116ecfc6df3c3165af1b87608ce30f609d71b3eb8a4939df93c05d6fbf777aca4ba6a8d5aa175257da9a4d04b9f5249324440d0cf595bea3040337fc7cb73fa0ef99e5281354a9febb1370172183b7b879756fa86a244eb85863bd6f1ace4afc3ca26adacea81852f9f661a2792c3af270c3c7acf3187a67d6235823a253cf2d84662511ada7139818c1ebb66b125219e78553df76f67a7f855f811be416f81991389d42fe123d061780cdbf2077f3ea87112f29ae410a5f82f4a4b816643d0890c0595713535bf91dcd4e3f68228d1a8af63e69213eabada8710e50466a696684be70c7ca61283f121ba00df19d0c38d8d53f1f19248f26ed4aafd03bf29e8f46e4ea32afbb58db564cc287faa227d5f2b49e2eb2a2a702355f15ffec0c559713931fe1705d88226598c6f30dc774bfd0d59f302597cc43734d7546e9e486093cfb77783de4927349f45d6a28da2158be2be257eb076c7feb2ae7d7a5a36205ecd1df45a23b33aa4c3109580253ec9111a9cc568dc035af5581a5810b1be20557bb40818981d1a97a1f6de91bd96ad56196de53dee01bd439c3afc443d34e58a695a489a86fb6cbba84c0efeff141455401ef5b5a1f5ba7f0f3febbcda00f7c55c896aae2833018d73f270a22689a4023c956b5dfd0b024036d491bd952f48d9f9e0ea35812c84129e1504bfb9b7440873bc5344391268a519d51dd1a17229e6e0879698c8c71f58baf133cb13628f9e84b0d75427469a6188cb71c01e22adfba887652d776afa99dbb2d5a4701fe1e75bed3f930d85066d73b08b44aaac4857220da59576c4dd87ddede7a9e55664e14b3ec2e67effb0c88db5ba461d9402000f01f47fa3205a66dc256f58cef110fc452d425d0b4c6021f08184099b60dd21d06122f03d7acfbb296297951d3fb4b2731c1f531998cd04643e0b0603e970032e2d6650bcfd180fec2a2ebee4ae2d271e21df51cf54863624e6ebaff78a4e5fb1823429404dc0d4165538ce653eb16a4bcea610acb7c3d53bab8db90120f78c250ff1c7c83c7266d49322a783a2e3f6b7f79adc9fbea178a0105183126da7b8a4e84f8f7585ac1e1f7741c6d34702512311320dbc81680ad9190c75e02d3c08886060a4a2c30874fa825ace6428ff1caac50a147f4d3f91061361bfc8c48b1b05bd855571135db9611c9e4cd324a47abc993dc6b4f05a76a05c15078648d2d6e45ea5ae46920cb3b4a398de1a4df09203c8570b760585aa58c9e89fcbf08ad0820288b220d67cb4cc2a2c4fca4f5ebbeb8c4f83eae9a0c66e70f1864968a0e2cf46611605f46351dfbba2343ae9483a989afef25dba213560c77e9c9553ce4483ed974bc7ba2f7040ef1c69ca979d2e5cdbe6dc780ef5e72aab0d1c229a0dde0ecb2b2048c6e31c3c0bef677d8b6d3a57e910eaa48328c416d48a320cab2d4e1dca44ed776052b7bcdd3850dbfd05866f130ed6b624e8e43e82c2a31566b21f12d01847ad259d07fb34af3bbd27800cfd5574801844348df35236a241431ef99e82a680082de1ab067dcb9c0cf54d629ca6ae81912c53048d81570c7820d1bb161ac8ea368a198e6117a9cbb896c1a0c6a0e9519786db1340bfe0cfa49e418af31c4d787979b20d8ae2e3ffd98b9f55eec994e133cac611e99f7b319fa3526fcde72fc948d486f881310c03499b467b4d5860a65a962d7be525279392ec5c91bc749b54ca401570a307c55d17513a30c182d7c5d6af86119a75526d42088f38144ff269d97a90d517557fbd9af529f84131655321e448a27c883dd8d1eed97dded199c42f86e14815b8cbe86b777f006f123a8a8a0683c7516ee5e060ecc02e011d4781535e944cba48c6f1a1571f9e646d16a8d81beb00da2a42df7281fe5ca3994d18c097ccddb2973c41dd52ac45bc7e4869bda7f2003059a429c7d7cb2960f43b6f022169748f33552f324d73f4afcc83b7553c14bae39ba7d9c45ddeee503fbaef3ac76974847a7e47ef08da1d79756bbc65a51051d281fd129b6f58da60ffe442e85521ff9bedde657091f631059ce871ddf28fc5e51379414f32fa84d78d565968580ecab89de541949bb86f57ced4fde870e012f684fb5a94798e5249cb8eed283c94d8015c7a9134365000d9a240237c3c15b8d3c8e820ad2628e40b1e100db618b7b4445157e2beab4a620160f13ea123f0972f2e54d770bcc9704a42e949abea130f4ffe2688a1da650906e15a821897ee62964fb769f4c69f9ae75b731027086ffc0e68e6ed56a36702d774f4a76f1c345cfa03f621a75821dbdb454b1c4c7f90f744329b757786f7f50831e80e25a26d77a225504f5a1ac31d16ba19f2bf15a7a88a4d74b2fb4c97f672a7fd837d860128a085c2c302af1e70eb795c736329b21aa5a6e55c3643cd14a1e82f4f22595fdf3993cd62d08afc7e4e0f198008359789b4f548beeba464bc5c8c2473c1ea5d03837b8d978146a3b46e87fb7590c634aacaa9f27e441c005767669aee7424aaa5324b078a67c440aa325b6245a9944d52382ae8067618935a30e771f92ad64724fc0a71885f32f4e060fcd45c382e51160b8777a8d29624f231e4a6fa99c23c647a80b56858aa89457e1479cbbcae2ad34257a31fb5efe3211bfcf79a71b67f8f951cea7aa97b4f07c27ac75ef71cd916016438bc4029246aebf3b3bbab05a02d6901790db79a6dc105544d989b47822683ad2b0eb6947c9055442f170dbcb8e5f894cb03e0d847f6033cb63b4036a8d8c119add522502a7c9f04be62394cf390e11bb2853c2e33c8eb972f67d4fe0f5d44774e8098e5a3a3efc20511bc019b2c2e28acc47ab02f2679be74411acb83896bf65655f5439f00fcd6cec68b68f15b2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4452f595d29e403636e4f25af67824c9fec5f5f95ffb8093c61d3ea363a74cd099dc40bf12a419100057888264c1cd52880b390f7ee936b92e440d494c549f8a19a17d69c4ff611d3daee5d3f003a87b6f7c343a5f7f5b502825cd691e14d42cff603cd32c83e2013e4ffe315a1e19fd377c88d1dd91890addf520a4f93e5208b492e46fe6f23f302add22a9f6f4931807669c5b523a271310b73822d875738b2395a19dad793412f7dad2be062a0090d0adf5a459bade395fad7b58fac683f90603022b65f69d684867aecd6c67b50c05e8285dc5cdff0255ea1fb3aa87af3332069600086bfd81d71a911e3bb104cf65541a887a3de1e618de2dc49c7df09640725cb2917f539b9fccfc678f965012dd88f807b7bb97ee8f83368e8db5d56da8b83c549ce679ca6ea7c36d5f08e7ec8304a90aba9d3a07d9abaf95d70e685dbd1cfa226e9150e2abf9fea795d44a97c03821a2c82a44068e8159cf57cac29ee4d837e2dce9ff17c45f4751e1b0512f74a1e7739867c14fd50a1b5083c3b06ceb79b74bcd22432ce09f774432165b33576122aaaf82f937cc86660c2279ba887903e81a573daed46b93df5030fea123032e1305e130108fc5c6b01a581889c1fbef44381426f1e2b42534312866bf5b6db04c5eee6a711ff20180d3566d80d3f7113562a68bf1501e04cc2da5dd989042eef7e182023644d8a8617ca0abd996cc5d7455b3a7671eb3000e77909760a9eec48bf8fd9096d58992367c1005df3d04eb3a40809796a30d88911ff8a57044e5736e92b303a533de0b5d9db64985bf73f9241096eb428cbdc1b133024895969a1a86e25f1e2351c49449628bb37623017800840f5c51717fd9aa1647a2c8c32ef6f199da6ad6e2f3f7c08ab86165512524bb6aba6ff821d2df28318bb04a65a56b362a93c33d3ce525aa791ce24522dc5775e11794bad71b49f939c991d3ad0c974973749aa6091d1eb92849a72a39bdfde49c28bffd8869cfeef9d802f7ca31c2a45f92a4a9d847def61ac01d0f3fd6961156219b34f6c37981bc74b80c0327721a0f4f9d41890ff4c2917a469883612a84e6a1804cdcf3fa33774dadd3af87860294053d3196a8dfc73dbf2d2270cd4a0bcfed2f2296943a3ab07555ec3c5d577701830072b30a2b8026b8846e679aafd381064a65499edaa21dfeb455dca39524018c184ef2960836648cd4f154174f3e2cbb72d2c95d7faa0e03ce617480d94fa0e9484a5a250f275aa0f2839185a461d2a0cd2a786a79823b713183ca178ad60df3726dabdf2bac4f2cfa87bd8e96bb0b3ad8df2a6ca118bcd54b6a2f61881011b1a2d38beb0f613f9236d15504dae4f37c974da0b9e03d5d4fda0d0ff88535ad79b5a5c9776e20d20d2317fc325eb4c013c18af3c524fbf1258ff0461fd4c1768537820e5e6c8b73da827e51c78dc7c4a3f03e0e4b90f031401466fa0ffd55797db661f1f9fa83babce82c61d3e7b8ee50e842e1e4d4f3e672da13729fbf78dc444260c9f00457c80fe83f82b5d54f804ee5fd51b6007f92ea274ef09416616b16646d01df6d786c928a79a7bcdee2ab2a111672d5033b137f8d9db84e59cc8dd152776321bc5f958ab8aebeae0a059f6a65465a10cfcf0f0739df90e8d46c7c82ad3d0e129ba2fdfe2627300dc6efdfca2a7a1816b83d33fa831bca284a5fb2ecf17e2b0afa9700924084abb21b3e7fe002f966cdf1804d3ad1f5ac74c74a7ee3d546ba7502e73a824c155114e8b15dcd2a399461163d394024e1e5bc59e5df9597479b6e27ac44f6547200a1241bf0857d756a42c95945096170dcfaec06c13dcc0e1a098a8890d55afc51cb9ce6d81f81951b17152b500ce3d4087a4715c313e2cddc86874f947b9fb30e45586e0cfd4f96a02f916f484ba3349795ade81696b3dbf7eb16c4e2b4418c069092ccc812d94e0c1fcae0dfab280c0fdecd6abfd7a0beb079e955a09346c15a4d554dc6a36156181dde06e8e9a13b1904627657da5ad714c6fd6fcbdbb8169ed36faa6af399c6c3c5184dee761702ac69cb411bc5257d4b83b31b90ea482dfa2474ae7cf2ee04570d8c7a9f07982404444a4dbe0469e135ada7f247edf2f2a56f978e3a45fda3a34d7f2046cf796f4dd0715bb065d770b15115022a7284ffc48b0e2f8abc44cdf861a24b397d3658c56c127a66143c918a75be0b828d6eaefb903f63449c2ac8f813fe025478c2493e2d7fcda0d2167838114d8a382dc6048c31f15aa31d66e224180cb9e556510ec45ebe41e5c529047b95d4b0d791ed9deae1efbba5d0015ba5acc55f7f9d17d3bf7c69d7a87faccaed012a24af07af0e4188508852751adf0c005dbcffd73ab1bd06fce7a877687f2b3512ce54c3ad0438eb3b337a53bffb24bca4cd09f00f360fd4082174014f1324f62ce679984115f099a0b6ace4880236364b48deb69bd904ceaf9173479c32c3a5c11e675d0815bf84550ecbb5fe2daa99f6fc066aa3ccd68e96ec9f8de83fe9445de2188f0f5f94c3501e7f17be125ca2a48b24b769814e87d4645d6a9e6a76341c0f7d648b6796b0980e20960621f7c9485e21094b6e692abc644166ad321a48780bc306dd63235c3afe731e6755a67349dadf4d60e4f1bf7e3bdd9b18a3ea568767468c7102d92aaa48a5b026bdb0202a10f7edb511670911dae6a6d1542f2739e169effc7a99ed6bc91b5dbbc90b6edfbb866aa14ac0f5d81301c5634fe0fde5d1ed915ed514d7be98b228ed5764bbac4a3c07f0903650f32005a9a0fba4a195faeae1b178c4b682792c317a3fb9b5b23ea43a5adfb25086c2b8dd0868f483d24f41a0fb7656c233910d59e7a33fd82b47f620c27169eb2fe580f5d42ca29a22836d5c4f12f7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4a100f1522c69d051f0fe13bdef7fe87c8abe03ef2ccea763c9bbec86bd5ac49fabcebf7d3f9cb20437d788428e890d8085de426f2e21295525c8c6d1de9b6395f7a617b8a87264a1e885d842f88f9b60db23a513c7db545617cc36bc1ace3097702837f26bad974e6d201b1ca4e61f9a2d6127c2b6f755e669077c7de64175603770892ad0587101d48995fe26a0c0037f140d836eae5c405bb7e1c0b4e466707c381988753d71a00ceffc552f5d9981d4e69db646ccb9437ff0357444e493e51617cab900d208525d6ac8340d34798bcce3471c17428e6dd2ea12b3ceacb496c0b4952932a0bf6a1c3ebd4c0e5f9fee5da1aad338c0deca3fc40f390a6fccb3cd5057617c4d6a49cd0ca43d2b3bfa27b226d9ae7480f4788b8b15be56f88cc87ab2fa70546e7170917a767d270ced8ee91f2ef80f149f3b041e0875a175481daa7afc27633bd75312d817f04a2914b3ea58b5349184015e960067411d441945e2e86becc6dae83182daf6c0895a6076be3b77bb76c5e4bbb5c28bc52dae876c5ee92947db89cd6392fc03f200441c6a97a76f508dc1e41d91f6c786e17297ef3cc8e475d49b1a26db64f6aa0aa4871231a9bf0e0bbec6410633ba4df952b05a9b5f0b28250dbbc19756314a82a385bd82408d1c156af39af5234e3e1c0983d02af139a83d98229febf2dcf813ec785ac081f9c3e3b5d53119897d06eb38b2575bd4b333dcbc5b29148b8a505d7eb762612c6838ce0e8fd4bf8475f50738f510785016fc436a6795fc51e0f6fb9a81fb9391dcc9ae120714eee806f0d7d7e26940ac466efd2b061c04fa0ac5fc59bd7aba3f6ded6d66f2c0113a2c9f12102c02ca03c5a161cc28b7051ebaa2b1a57a5ebacf968d52d8a69fce53feffb9c6fa5b111a219d49dee420a644b48fd7366281d35a25bb6664aaba1b71fdad5c8881370357a01aa8e37b7ab7a6befe697010e265c2939499568b8467e2478905cc4a7edf4789b5955ea638d45fb421563aac977b4506d4fd668cc2e32128cc5fd85bb337732715045cbc271723fbff151b08f86662356e7839f2bcb320a549c2f991e5dad420e853246920b5fda3034d3d1ceeacc73b917a9b168db3c2d4b9d6f2fd9f1c12bd273fb4caec425d01dab409c93eb7868158ad8946ab0c95a2aaac2aaef002bf4aeb6347af9fb79899eb4c3d0a096ce822682e7c0fd3bc5880365e9a253f85f33ea3138d6d6acfbfb7b9c7b971e848379933eae4fbeb8d0edbebb975e34095e3e3f02c44d798f8baa42c1a6bcad85691cf191e29c73410a64eabf54fdc5ede36e86a6c49cc91f30dea62130e59b24f5f6f84121923e0a0079b3fd20100a347b508167b6ebf766e7c789b4855362a86a1c4ce278be4d12a91ffe075260cc93761b7d4e8126138d42deb0c809d40df114c14e972c71bc242c02b1c2e5d8bcca256e321b8840652d4d09b9bac06db7771ef1dabc3bfaa5616d376c982e85cf0459dc7feb16eac5cfa9fbd8413c1a8441a2c4f046de3328de8467608e992a5c11c0af05c32512ad864905f3d11094588ec65918252b17aa603c920f731e2cbf757e37100fd67fc3f6d32862893f6c2ee71e6bcd69e5fe272f6740d866d5b5ba452f1b9b8f3c722a9596c9df10c3181d0d911986fb3a84f6e9a7e9e4f1bdf38b4019510fd2d763192f204ed33c9b4265a2aa1099a2b9dd1a877826af3440ee0070064ed8ca3d1a22aad50791d8230fbd8f8c40c525ef845f57d3b887659c635ea500d32b1602e9a4361b3c0c6ae810cf168e459af266876c9b47ace501a2a8930e220ea1ef878029020c46c57c091134816292a682cdd31e211817b08a2efc764ce6db4d205e7d824d4d6233ddc0ede05e621fe4720d558adfedddf14845ee57352704aebf3b6e432c5874ce36bd8e07cfca21aac937216cd74f45a81923393f3f854bfb3856cd5d97144102ded4bbfdde9f8c14da03e9b9884c877c7ba58fcda78e2db56598a10e4d731ae032e37a7021c0cbf179df81154860271bf03fa4c553a7456b2c983be7ce350457334b1f7b6cb1edfaae4cfb4e61e779a6166362dfe80de4888ddbd83f9022751ec80ed8a7d0f18ed54420126d54854a5dedd432ecc6ed5e5b65c9210e9dbb353fe13495f670698c2777d17959541fc452d9fb9d8080ce10487a166da491f538461771642c447e6db89cb12f8689142748d5863da06753df4800f8095d572e033afa1d736a6143db99bca6600cbb2d20d3f8aa468c94665537ff96a45dda63b4db736c77757a9a521238ebf5fcd2cd1e1cf2bdbadededae021d69be9099a4909c09695a13e8e43d4edbe97cac8216922958a222dc1edbda9230e10077bb611b27f5701c50176f4e4f33b008f7d350b7a4d954d592e2303e84581bf67c8237be42013d72221ba62013113f9084eddf5a5f28d5f3cdbd2f8882d13c1834b7b9cd7d9a4f13a3cad386730f725b398ebf9722fa81e7e39cbfef009c20060290ed74e73a2693beb5b18289abae2d0ea68e93b9a9ce97f24e29bf8e973d852e205d6a172177511791cd2e83f706e5b3c0db1548d2fabbc49b3d4c7537dbf3cc0a809e06541f3a229b127d376b0902f90e3479fe5138e1fec06c6950d47255518a7423302c7b8b3c6cd083f781415a35c8b498e89760414cd4503e7fa5592c08906558f9f36cc8d850598d37b812f4a233ade47135f84b39bbca54e4eb5166d750639b8cdc37c9f3c07baa630385397cd98b1f2b48ae25844bd14e91c08020bcf7b95e7fd3da73f06da5b456c4a139dee081d317037284ca69b3c968fc8f5bea498e25fc82af92742630cee72789246d1328f1fb7615245dbf2a0ac0b5c779092926bd302866cabdf71fb32ff5238060f1d58e81393a94229;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha9a489c4636202134bd10758778d2beb4f6f09d019cc9025c76379e35e5cc6c6ff78acf4afd50a98bbdc3e457763b15a2414d91c19cfa6f9932c62956ad62551301b10751bd8c86699a0e0fa0a572e0eb5b3ff919444151ec1ebe588b295d6580a92e500785ab06a9084a7e94a4af555fed97f7aceb0812a7765601ff13a11911fd3c405b91e70ceda340ce9225da8a2d88c4d037236fbada6fe960c31f529983809c17e044e64b242bbb5b25d229e38a9b0e2d5cb7ef027cb1242655d448e3e1f1f40e157950415727080f790e2c92cecbc28108fcb1bbedc4550e1e416217d31e29633d4a16fdc5ad8d4e99550b1c924ff252cfa184167b6dc59d03679f733e7612f25aa2491adb8da409330717b38db5b4e79112d8f69f19cc747ff8a6863ddd3bbd0b5cc51c495cb122579c0f2a8fd8ecffc49ef50c842d5f63bbb09a3f2206da9e4a638f9114e553818f22b587a30964a157a5712338ce9c6c9cce0dc655c01bf7352647fe2af327adbd46c291afe9490f104bd1d9f65c3c59eddc23a51af4cf43359e557e6682afff07ad13ce822215ae470707ac691085d25731b0a65d56138f18f858adc63840d607f26a6eb6671b683f3ef69d042b6b41771856f37dead61dded463781b9a6a53dd75de330066e2981490a1dcb33bd82aebfc164f187d7f45b7f8d6cc891f639d7797317be432775ddd173ba257853420db257ae64f5842bad634a239ede39fac254e2820d13cc7ebb4798c31303a09be217752c3798d2d2249e320b741e9eaed99c25ceb39cef2b47a483f7bb9179ae968a32df1f08669cf96e529120ad867460e7ca33af062446af0f97cdc32a1b11e90fcad1564a30bd9b7a401445825f4b831f5d5548f425407fba538d9fae6ef8413eaed1f1485a251de29c955f05e43d70e7028acd949d57377ec2d9c5a44e3ca649af5171c01dd2f90d139a449f78715b8740d1db4201424f02510c9ae55fff803a214a1aa0946c2b0b7664e80692c7c263349a066e5d2e889ed2462d01b0a16819daad2c6aa30411b977e522cf3dd49915399a1f6c7a8646f3371e62948af924c384673bad298659a442547089955c3b7926dc5a92f650f7b44a481d59788636374b2b9c0dbdd44abdd0923fd47a32494a2e1accc349b4a26a26565dd1200464f4031ed68a122c32f47270b9876d4c96bd2cf568d1a450ecac3941089679229a42c433bb0728c04b1a5a6a9478341f038cd6b2f6e19cb819c96c3d04d82d76b881719430038dbfe414b02c76392e112fc346c0e9ea6fd7b4851efb49ca7314c6f5d93bd0a4f4b07de7b6b4bf81ad4618f393114afcc3903bca6e06046cc14a419fc9a0cbf9298588352bca5b5db16226194d197c76195e345d4c1a775b32972ffc2d2199907b24b924813f91948dbc7ba4e55442f90e85cd6da9ac701ad9ff5352800a1d5b4c03f0e63949ad5565f91a94ca3a833794c8f53427434dab34445b6623da8e21e8bf463f05c6ea1dc9b79302695131a16878f658ca90de7767708622601235747ce370d6f12125c623ddb98fb62f6203cc6f64fa1bcca30472cb09f5b73da93ee8179d28fe72cf177ffdb519351adb9a9906e378e4920bb0315e68a5571e2c0d9a9ea4cdc6b591db23dc619b63f3199c64bdc7fc58cf69208f463c8cac6794f9aa84a30977a3d1223f9d07d9820d960649d48430fa5b726696db9540dbf2040d33f158e8ca33a5a6bd2941553e273c5c49f52551a9f87f70cb4f5d6eb0985442bf4aaf98cd63d837fd886fc77e7a4c6914f3e4914784b57eb27f11bb4eac1a99b6f450bcb09659c0e6661b26411cce29471f746fecdc9e64f51fea78bb3c5ae19c1d944553b54bea2acceeb7d8237391dc1dd2f88a1fa8c7b3b5c1c24858ea3ad2148a0a2b1a123677a225a020cdc67b830efab24e094974dd5f2256e974c13a492f182a08076a3f9828414c1c179daac8d866a967a19b499cd43d7ef29867d861bb8662ec22f30699f252a3529f1dbc22f8e0a2114ba0ec83cf689678f1cbf8411b9f152df6165ad384b3c124d00570576af65294040c5a09eb6840db4b7e742c02b90e067dd3bc0f13c018074f54f9f4ff926fe4d7d2be4efc38489f6c6aeaf16ef14a6cecfcf0451211814da5c91822e47de40d49ff19e0e68e7208bdd49dbeda3c69be49f3fcdff68f8afc0f6a0a6b875d6de7e50fc52da9736e07dee8049e75959056d3ce4517886527826babff1426f411053a94714c973e61187db6512ecb68b8e2645808ee01059d2cec3b3d087ed63e44181ea8d8cbb387aeeaa731e505b97731a0bb7ac500fe07b56743fe219358c46be029419545ac23f026a362cf518e83633adbca6b033a5c1d34c9d2a1cb6182cbeeede940c155cedcc32fe458e73387cf8f08bbb18e2345d88e00eea4a855708a7bb5607a6eb8a01bfe2e5dffaf17d065020f3d854d934309f83d748f5e18c1f15bb3ba6ecc8fccd4ea43954ac297280244250fbef7041562282892343db7eee1dc43a1cb246cef7c6433c7b432f8d1f14c458272ee5091f677d99c16ab2301347a889b5f3f6397cf73276afa45af6e910ce3c695ca03ee99b00595401f7530e63aebe35f0f587ac563b8c5611990240c2382231aebb0ef2a847e722a15a2ee6cabf12f89be190955e513a31460914bc5b9b2b42cef1b9fb43b16257fd0fa8b49f7bfccb717009e651ee490c2c4e4f7c98014ca6c62988c69b1ce5b8632e5817ea9f1185d7755effab8ec783dee1cb16ec03f7503c8cc991c197718bc2235b58312089c1e6a041933a7444daf06e8a02b002c0eaf02f8eafbacd4b91c3066ae09e58e3300d350c2d123ed8903ff235307ee3f639fea482c48ee59ee7d5b7ddc2b9f0daec21dc18799809;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9c7415a5d9546400e3c4c4e297ba62c37e22fef04371470d32cb3d36912290f33e5c5c8ee04e15222b970f2035ef993f625de3c9a1b7ea04a47556f145143a4e9cbd8e03bc550ed096a70ff4c455fa972b575c61ddae512425ecfeadc722856ffa04054091deee61f625a4755fb624df77f6d2a2d243d7b8223db0e085b3c8a048c323d81fc5e735e530f4dc0897d49354c5adb60e19b02379b65e5015257a8373d4ea5550ed471b6916385bba2caadaa480aa2c0dbbf790540f12ee6ae48a95452d0b7becbe6f26c37cec94c85f7448c89df7c6f981205d6f06ecd6a3ffd55e4109a7e7600401bb5eaa005b95173357cd8bdfebc570c33b6e548228ffe2aee024c8bb0f15fdebd7b7e6c014c77d46a9a6a209e27a122209e89e8f71df3c5bc1c35b5e48d8307700b8a9abf99cce8c144020392fca2b25d36c47687ac717e7bb6803ff9867f6f0480b19a2c0cf44a4934d6eee817427fa5791ff9b86dfcb290ee1c33b53e516c74b994d01e290e13cf3523e1c26c0a7364d62c4fa519102e7f14a5df910e39449252ffa6981111e15ff0de9e2ac7e621e4c40114b875065a4bee018fdf207fa3d572ccb26957b415e71433f3ba90d119379e14da2eb31189d406aa82e589d20e2dc7f3e53fa175f7b598afac9b9ea703bfe9518a78e99a0b7fcd51ae76e478c39040ffbd7261f108945e4fc098724597e6ba9ea3eeb7a6816f8b618157cc84111a1dabb0039fb64ee6014b0e8b773d67f2b81b8d9fbbc6b55567a64f4f20353420902169a2e02eeb81eeda3e1ffa7f406c07f2e9825c07ae8b11437c562dddf0bcbba163a6e0f1ae0d3cb0cf53c12d9701de1ea5caea80992e9b7afcf901d564efd29f3c2013561d18f81a19ee66dfd52a33abe4b79d2c124e8531eff3e74368f1f9c75fef6706ee5f57954cdb56e1ea77540f538c4eb65cc0b87f4e282a6c2924d20293fff2b3ab13604ace3bad41cb7d3ce9a668d5048033464921909d175019994b9c4e394e7d2f157bb27916d4ead6ae3a6d53587bed11ccf67892902efa14ebddcb9d9729c616e21ad3fdc6aded1f99e8c03e8fcd75e84bc5b30026205b662600164fc074814b5f1bd554a3bab15f3b620a1c4fae2afd6ceed623f45ca575ed446f5699e08a1274ecd4c68990ae47e00e3b8b05bd46e1db986a905de99490c1bce576e4e1b116f4ab9e67c8e02bda33bdc5f6f3b88504d53d69baa085e55747e142df4865668b2195a89a42954a0477ed6d960e07e5865884b5dd6075c2255860699b79b7a09f47f70e905c5fc52a8b5d86ee3a95343d4c1f5c082855faf1b08fff89428402ec6e4007c25d907c3fb1bde5a6404c564dcf799d805474291c376faf4289c25dcb0f69848775d3edd04f607a1cb3beed06f634e9acc6a1f780493c3678b8caafdd359f030360ea09e6249b158513eb1a542ee4bf7a01143dda23f8f3b7ff7b71bc9b0217acf66fb893f87c2731e9bad89c45bbe85d05c8403f47b9391347da91f9f404f0cd0d86c040bf34199f5b1f70815f4fea1630b97b19e1714b7901df9db77496d0ca1cd913288ee5e7785b898e41b8b5921e8077ce3a0a04f6772065fc4c19d5b1dc47765386f28c0f3a35871b2baae3c8376e91f443059f2e9d59e7732b36c6ebf4c17fb6dbef423d95d8a516ac0fba90fd0ec070a3f49b40ea65e2a2e5b6883c4b3a592eeea64740867f4590b656f3b557bf95c06196f2e7268965e0d9c19a3c6c42488456417a4c3917dba45a3af6d1be2c7bec1ecd542a5864d2702f979ca27b3238694bf0a6ff586bc8ed96e7a45184637eef0af49a6c11044b91210063a662958a1f7c03f13252d3012a742686f8044f21a88f28e34aa95b10f1bd9a80b41f64c63e1cbe694f90d3f393cd19c901f26ef0b3a3a03605ac60ca027b91e1215ab8999d77c31e38ca1a23e77bfac5960fcb0750b21123e821d9ca21a5927e312d32ba2c823133bbbf7b4828e0fdd4e22bfbe167370b9d33a424064811811307ef1657967691c698da1116f2d518c407cb0a89f73ffb18388bcbcc13c1a0791e82f1cc4023dde4ce8abe05ffefc620308401d920c225133e376ecc9e325a0eb7164286d56c8521f989321de36bad391fe2d6fbbb7da3a92153fe05743341f45c39a5baf700687b250b44aaac456c541026e063dbc5ad0ac298af6c12d6fabb5f3c507db167816f0e5f05620da91c8cbeaab2f7bebfbccd64cab57b055902e53bcbc61b23516f051ccb6c21827356829728b4d8ab494ff3b7021ffe24f0cbeff2f3f4f33dc016194f7e32a9f1b90aab55aabda6236446f021af49dc9ea99e90cff2ae3ffc5dbc59f11e7abdc9fa74fe7f066dfbd50e61f8feffea78df6eac0d9a02893002056980c17909a23d75308f02d84f7f0f8fd159f9f91fa07f947eff6c59f6341a95ae9b09cb8b60c0a6f954dcdcd175c22d64ded5d4dc7daccc657ff1efb91b00c78049af4fb8ecf79904a61f2fac8ee9151590d49c0d71c1e4682ca0d7e21fdb52a21de507a6819e7435e5d666a3ae3bff26859a5566adf458e56082fb9c21dc2264ae0db8c356d2413eb1d395b425b838e4f84532c93f0af4caf87b351ddea4dc54a3b606a71a0d4d5dd7dedc7f092cb7ab03a5dd1cb8f30d6e8787f4b521b7796f8cf04ea639ccbd0f4e9014b92518587607c2fe9b94da28d590c7809e472bdc7767d4c70fd281621a27f6a2d6a2746a881540b08ea70954e451e5c6da48a09725979c6bc34f59ee1f8871756dc8c792bb280ab73e028b48b55860040e055b3c8f42c999f1ebcd9ff1bd46c38258a4492c41113594259f74c59e7f3fa46eebe35014dbb21b1189554f9b2f3b2ec2afa3fe22dc43e021ddbc842d8f8784dafebb1d77968011c977afa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1f3fe92966451f681ec887bc4c4cfc44f50b539fe8b7f378bcfa463f977acd97c88332ae8d39c23aee1325818911708b7adfeb797efffa17445803170deea3fa5ef5a09555bc1d7c4a3723d670f2ae637847a5b7e020b43fa23bd3e6c4498ea3ab929262d53599a6bfac5f89e8c8a61b76df3e5899e58376a90bb0e6265ff1e66da0300f060ff8b2a26a56a9357cfd8600e83617dbdb6944d1ca5cbab15cdc8ce8ce04cf211ce46b68fdc1c39f19a61bb1bf10ba84724ef000ac8057b6dd7772797fbbcd074c1d5faff6429a21ddb4bcaba720769fa793f48f9642fb95dcf4698a5cdb397769b10a27cf0ff97d8c6bb817ed0e60e6a734978d905658b2170d9743e42b067fc09250b73960102d1813fdfc9ed05f4fe58b9b2b75df3d424d25121167f0b031725a936c10ba0bb2e112daffa6cb6977a4e95071bbda16d27a374bc566a6378ec42cf8086cf3f22e45326ec2938b4e3cbab9a8b7ae6f265a6c9e9da43f4a880a228e6279b17948a221818ed935c7b9e6670d38452f836f6683c9bf4edbfade5b482d4928145de5cb8e9714286025bcf26ba81e9891e94d3bacd7cecc7957504744dfaaa95cdd94b783d60e3669d70133f090a2549c32aa27d5ad6ab7eecdc9e274b9dec290c03b4a8de59ab9614220eb925b9a689072f75bb37a803928152b163bac9ca1a37517bc91ab67b85a05b4b890b1197fbb4a549955590e28b7320619b2e0ea98659935aa3f7732b5845de7dcf35f163b8a1a7fa4a022db3301a43c88e3a82b892bb65d17bfa31a84b99602409d322a96ad087036b743cb2161e108d5ded3de87e923bf05f1fc33cc32a32ddbeb5ba834e713bfc3c0cc6b5d64f387e16d73c5fb3e9f2188f66109baee7c3d529749e3d22415f1dc9d3a968498c1d8ab7f5f06e1dd5493d20ce60b41e976fe284abd81a56bc20fb647392740c77a1668b8ee9bc50b2575e6c3d113ba0b29423eb0dad479b03204d9b4b0b69a1e1b9f3cb7432fb4940b1606f42589350f375c4dcfa9f47fc8700d292068d466eb6ce122b7a3f38a4f6aa7d4e4d8a2d6ff18356502f2b1492e7784fafa8c0e0354965194c8493833e298c8aa34090982b69e421c0abcb7945bc03cca956a8679e3bd4561f2e05fe517ec37cb49b03a4d0f1e3aaee24e359ba74c05123cf253b38b1b6396a84d2e8731b72a5287d369a4b8e3e56a9cc2b8479a53f82bf204ccb9953d02fbd971035f32741ec52ae30900b8e306b6b628e0f25991113193f811800012eb2f7f6dec19f54ebe9418fff5dea83850857f52e1de4e0a479c134283406c92c0a8f38237a2954d946788bd41cb632b2f532e6bda04238b3da2ae0309daea415b3a1a28db3acf68ccb23b40e7b1c238d2854530f786699b140bff27d2b5111026fcaa23060b47f90fbec67bf4cb9b322bbb63c606c84bcf5c9c8194131619f59b209aaf40762d4a6dd479f14770e1809e4807608c2cb39de2810304d89a6cb8aa1e1151731dd7907248962bb3d9cdcba3df59f49ed8872e61537e243d8795b5a21a277832839b7e84b3520b644db746845b78834c9a22d7cad8cf88996ecc7f90ca344263760dae64eb004b52139767dc085018618c6a577f33d4c1d487a40d2bc6da3182fb93bed52dfea79c9f323d367c76aedc2293fbfd11d34aaa73160f437be2baae6c5e59ca4733e6cb77712faab3aab9d4ae844d30e719af9191476b05580806610ce634cb76ef7d79f3841a79e1ce0310b79a0ee1b4bc15bb814fe5a6737b83c1252f68818d93c28c3425459d2beea41dfbc268a9c53d69ce796a60e95d377e4479bba26f3eafcfce5d1ffde1db767b8feaa8088829a59d0ac8c63f814116c48cf95f80a323b3206e266c343e45d70190d8649e8630e82690288f0e678d78eae36d19ee50698f5932ee084335cd81d854a653afecce12db2e5ae528d2b8a3fc9e36a7d0a76d66b1fb05afa9f0a99347ed21955a0023ffd6c8aac59267852dea6a258d352cb7ae3f49d776eda4c3f925e39b6a1fae8da997ee03680c2562fa628b51dd4a61397fad4f79040b516c71ebc429481d26a09c4276b0c1a848d58ace550bb572ee95b64463dcdd3d69373ae5120809ba7d77dfe7d1afb9dcae6686bd840aa2e37a8364d4f005c8f4bbc88b62dabb9972f838b9ef40b66eede7bae191611530c0bc43014bec5f933d40440d26c90ba4a055b1c1f3d75c0bbb9cb634a06c91291c43b3366463a2d3945f09750f3ce7189d9a7c311275eafd8da5027440750b737b5cb72028d91adeb166ce1b88c0a2bc8e60216405d2c8a29ef19c0a2f16654fdfef34c86a4a2c8811565edf8b9ec8220a8cd7d0d392c72e47db822e7b84b36d4965b5b53a9d3ab8c55dfd5fd43403d92ed5674c0e64f26866a36594e050391db48e6e05c780ed032a0c6ebd7a810be10d982b737a4e855a754a42e036f4f087441bdc119e4ba2d9df1dcfe1e6fc2bcfe69180582a68ef852fe1287e32129a3575004a29599038a490b68a6d6cefb88abb5b1a1330696a5a35dfc1f3550179e9d2efcfd59c03e121777de668b89166b6eaebdb4711a45d0b72f4ea01f2ca23a3d3622d8e88ddb3ed32213244619cfd28903ead3f80387ae10351d99f8c4ebaa774ae3fc9cbcff135f70efed12a3d1d108d5e8171662cd24f0df5fa51614d8a9b4019b96bdaa50bdfcade02da69f1012f8ce2be501d7e2adcf6359146a873587d33e31c09d483b2f2a526e30b020d0de4464a638c3358479b7fe912196b670f439de1095b8a248f557b04029ab7ccce7304590af56329fd6ffc8adb4dfc767a108450f5d0c59f8c60de94a4e9760ef8dc47646d54dd6597eaf88ec45db188fad36a59da1ae6ca930257e284f67ad63014a4c57284f09e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hce184e8ca27c141229c17bf1a9cf1b55c1bb60ab3d223fe8ba198344ceedddbf8fb68ddfd9d50196335a365af334ee2a93f39279d6d8b11b66cf7f3949d7671488dcace74c8070a784bdc24a743c9df3b55b8c990daff2c5b41f01875929ed7c7528457e09b0f8451e70353cc49abeba00b96bc737ca926720253ceaa63cd420833686611060534287da8ed9df918d8123d9fcd36ac3aa6656a99f2a4ee9cbf15e37bcdf03e267b19861f0ec6c055e3280a505adf949cec4e5c6dd47dd89fa40b5967347394021b5e2ca8da952948f6e9e7b99ca6e1d35c6c6894d8b8b13cc5c70de02b4cec77ed2c9037bdb6d572fc7eb5407f84da1a87c76002da24e21b1d37e007a48ae0159d087fd6126ce1b29fd8c164be0de495882d91a761d8b3880406715a4885583c0e9ab0f2b537022afd9046b605a0b9163a5de639d0e9c4422e969a86f134015c6f5983e12223396abd842d46898b319dbd2a9b9623b8671c30cc42e899ef183dde463b9b61772c6e92447fa700342455fe75308ba0ab1040611b45027ab94cb868da4ab8ae381243e63f1cba9ac2bc434fe3e30176e354c7cf81518338aff8481cd2047f3a0826c2e73b873877607a1e640419066f1bd21869ccbcdfcf9286b486fd9690fc57b8b943e3a500dd5aa89c733490ec781348d104024592e05c7b1c64fa77667d9de753aee3af3c553f99c75a932645327add7cb3ef3ebea3c9481620bbde62d1b790bf4b8c0fe4fe13febf4098c350f28391f004c742174bc665b0a8e4d01b6f79f54251dc06f544f304cd170a798bb240c934f6a6257eb9670ed4e0dec61e3095a3b9d87f3bcdf03d17f05415a212a0ca81ed9547d930008a0de5b35e57a9221432e2f740f782d0cfa702a9d5a61af52fd7205d9388151d92c9b340673a8af472afd4be50af5a32bcfe3a04f0e18f335fc3d09814eda18213f16792ad4fec3b5d5352c911b27029edf326836178bc2d3b44b1b62b285d9a0868ad3a8f00e6cdf6946108db7c8a60548d2c0c582a5a76cc2393dedfc0bda4a704944cc5da2085c0f5949f9bee89350f6effc0a0db37c6c66c3347d96721a47978358ace586aa1033d1d83ab6241e8a735ea95eb6d7040874375573ea110461adc72ad731789aed0a3f76731b538ce20313b29cfa9aa1845d3bf09ae57b95fb23f8a223315c10ff76c1e53702b7457be5a12d13c7b48eed47bdad489613ddf60e86ba35891b08b043638f65eb955c2d479ff8df9b761c14ff0a55c5730a781d7bae92abbc222c8588ec375ad17da4b880094c896dee2c4740ec1805027599657070521ccfa90e1315aaf5578480b1350b3da74775f3db94321d0dff1cab790b92c5c3beee24a30682bd1f367bb1df2a1ca5e91ddc450f44a4c32195aedfb76747d375dd5310a6acd3a89c37532a69e1870f848a151842dd8fcb2032b26710a5b7fcb07baabac7f8c9c5e29aa1940095bf314a6111195bf0bd829d6aca0460b39543be468c54d9c33f409c2c9805299617146dcfd8e4e365fdbb19000ed12e186c2573090d78e8d824f09cd556b147525ba2e898cbd757673b5c533f1705ab516b5182d78cfc69a4a8096eb103ac703f8a74b2ace941bf6267224dcec69fc3ade42223b408634b833a5ddc838766e9550694fd2dcffed50f548854c2d0457e33cc91bf8f69f5f0ccfea0211e07ae4414a0908f63b217c9317fe3ef17195107c23f40558c04cb4bd50f4d44d45e0354f9b38bbcea70f7d35b1e7d8aa5d8d0d9984942e5e357afaa45108a0975a18944f037f36ee34a8ffeb09000266989887a57c2173187f47d3bbd13dbc9288c02f2c3f2f5a777c6547b95e428577f9e00b354172893ec175868877419a336f87731b9d0849c38afd18ebcc6d95ad609092f6797d20a2968f9d911ad37d57a275aa89e8fe94138fcb1086b72da15ea36506f025b2934d29120bcdf5421182fe83c7d96c92c320abfb7fa535760272501586281970b69cedcc02bfec905612a4e5701a9e84dd7e519f75ef93ad6de99e69125180da7425644228a372ba13bbfb0b4425a58518427fb4919e96fdbadca7e6c34db415350f75282d2826f3f1abfdad925834782c9861078ec251d3c170de0f1efe961600d7a43b4e3d74c613692fa7afdcfdc837d4954f7413b9e516d7971b6dcdf1d14c4951d45b308fd65b63bc8e9820151eb8d70ed5ad74742f31ea4de3799bfa8a7f1d5423fc292b0486598edb62449761f861c6bfa08c59f5e20b8e88b75deaa8964c1ae45cedeb946ec7cd3f47f6d8a0d5c4b9e3aa865c96928b46b866300d4d7ed2ef0746fe01b2d29d8f95d9cef53f91b6517e221f0be34c51ac81983133b942ecfa5c3b54811100b17a1e1ef12c6ca086dffecf0b8aed2ef28ba26151320ca41dbbe1ca47752aa7aedeb57afd32b2f334257eb5163b552f5a3fe76161179c1d5faa683f5d5e3a9a286e04c465525eeac4607def53454c874ec23b01f21e3f9cac571e88247675138b63d50d54a6d3308a2e2d48541c16725adc5a494440a21816de2dc550b445ced37d232b102404961ba825d6c1e5ee777ebbd4989c163a262f556ea40b603d5fe57ec453840e4dd2f0d55987c7ae7f44d0564d735356d9301cc1c5d3ab869eef7e52a3714a41405d7a5a97508c302ea7f0177287a70346e26198a5e96de2d794c2d42731401eea23238b575d4b1f8b16bb47fcaf6a7cd7fdc4ffc877a2f918c6765b3fca7fc570b8fc9fbe4aba8a1c058069f16921a23029d894c24f7e28d386e8c848f3300f21ffc5b59186401482b4f928e306ecf0e5b2814ca5f47a31e160642befd54cbbc22c3fbf318d3e0968c8c4cab6249578c7f43a1b54e1275628da743b06b552ce1518e3d10f7bf154bc6a66;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h47b923ceb575c31b7180996fbebbfad115f09ad66d1ea14846ee99496de25a568cc81a40eaa0b7c4ef48aac6d1c387514103b0ff1ac076fbae9bf0079956dec85178fee9292d92a45033f40687163e35e6892e8c1df361ad090d37db8ef416df56a154f97208a5a597266b5d6954f85af0dd044b37233d8a296cf9915f8ff030af5f806b3bf3c2c3c7c0d3bf782fdc1c84d64a11036041953f993f2387c966857167fbd696f30419925648223ede2219e23d91dcc0b34e7f97046888904baf674bc20b9373aff69ebaabf2eef659d52e7b5c70d8414bd82b42009c2da90a28efd0ccc46aa221b55c76b4c7cab749f6195a6ee8c1afcd3ba9ddec83480cb8deedf527f0a66833aad4957d74d32b71cfa4f8393edcd36102e127c985dd5a00179adda247b48fe4a6daaf80f483b13f3fc4a16f16f1930154b8e617899eff9e4694ed143ed0e0010db1294567039ec26b959283bb09530096813ad8b305a8acb5b2f0d170b2220652fe5299e65761de6a5f6be5241f71c61167eb22a91432339dc1275ecae6ca7e8a6343233f846551ea132386b1c177fd980dff618068ba25909dafa70eeda66e4b404d64b72a257738690bb6e33abcd574eeab76b37e6df120eaada694eca1b7039b4f0473fa66f907461233559ef89428def7d5eaa392df0ed7d4e3b7292202cf231c9aeb9810ca45dc88b61b74c20b06915de7e5ae627e1ad97477a0a84ecf6fe16f328a530dfd6c175d3c1a27d95c219633df5a1fd6d6fdccb295498fdaf74e5a92dcc40932e73e488837a11d382387ed6000f7d07b63b2d0dd02f298740bdd4d99e8d6bab40dd4c071b350fc41d0a3f76ce4e0c4326ac0bc84f9cf797c77dab8f5e89791bdaad46a83ca7a88b3f594c9955e99228f00f5233dfa1a4572ae416449cc80ab8368f821e59f2a60951f9263baa5df8ad5884e313077ef1ab6282c64c2caa4d16a118bca58b74386077540d269dbcb909c1d036a914ec30ff19522cff7611481c3fbbe82ebe807c31412580a06eaba37660372ecee8ab070680b6d8dc5820f6e80efadce57918d41ae95aebd0e3e153098f3570e53d7bdb10b7a76e66806c68e727850d418f03022b5c4df98c843277a2dc838ff9928fdfbb58104c6db6d949de0af8327462f972b49285c6cb18823920d230e3f696b1b7a6930b326bb330da3376b95942de5c37d45c612152277bf5ecef0baa7a56db7b08abb17be9d3fd16c1467c429649d35d9e0255cc4f8dde4f32dba84e630727e394bc219bc3620eaa62e015d676603b6e4da6670a6ab32647abb375aff5dcb78db2ca6717a679f50c851dbc7765c10f93d34cfbf10272f2703696540d1eeac93b4a3c33659324e7d5b94a3c32de213ab6d26d79b40f32bee321babbda3bf7377d476a17070b6b5e7584d3256642bc6fab1ec7eb543bc3a846bf3d0c7aa1a9b44c75aedad848ef7d26e2ff707b51fcbd3295622448bd419b8386670720c4b76e34a11789632a2005806b9676690ea63a79f33aa3fd39f6d2bb0df83e51dbeb5d4f8b3508811a33b1b41169eb1287097792e5d81d68f7106a5efe8ad277c3f84068baa940fb6310995b82170869d7d6aae9590f7f1b9ffd1f0129de492e468ec96ed24317e8138f6404396e024b0dca1b2ed9ffcc46f155f1a8e07b98bb6f33eb4028696ee59f9c1c9f43076e3b9f59f10104a11e1ef860d1e23be2d5956ec5e74e82abb33ac99afe5c2503eb6ce35ef29e4ad79de61524352abe228ec18e7e1b1ffc0d4fdcc21d0c597069f567bcffad2da43e66b4a49be9656517b0ec59e62023f06b9e245c5d4214e4e286e34e3edc60ed158c943d756040b9ac78830ff50746190a27c5d01f3a77b5b0c64ccccae9531e52bf83d165da3d639490788399f7fa995b77b6fb746d98f01d7f61133807d3c8908db106fbc9f4b68dfd3db4e45514a88269ea318a734baae2179ab12e2a5872156717baf89b77e1f7f92fd0feb77e34d828243919768ae8dd62ff2228d2536755da90198d2d96debfd23f1d3f2969d154b88051d909323f4e7fdd25def382ca7bf8275aa5f71c3a486a3180210df1fc9661099357aff694ddd6ee2c39bc5fb2f4e952479449e66aca9e47154e3d7281bdbf211172830b987b9c3ef77c1df1c8d64a9d270a230a0dd6d3130439737563099df0dd0f6c1823530da17b5b7bd6be044b0ff6c231523e19cc379aa23175460b25cfbec7cc9b11532b2f3fab89d9ef868b04c84c9e1888ad8b56c79792ed5e452ebb79d661627c462f0cf682b4b0eb389270439a0c1e29585ff005941f58328295a831e7db1344ad2cecdf3172a8976bdc63024dbc7b9b569e5bb27ab4ce3096471d4682232677844e9821a392be965fa1a70a997d2ba8596ead3975bed779be6a6cab8df11df9d7b6eb6166cb1f284afbd22371e5e2c484e3a40d8e0cd2efb3988bbbb23887f917689e1edd25034261666fcfd39846af12cbaabc96887b9a4fc3e92e81185a2a5e90857b1f1954f755b915ab1f21db9758c02796b1384a678e7779139646567a7a5480aecdb9c47b78f187c84457f6951dbf24b5b175912709f40e936efdbc7188f12fb8ee263c4474ebfbcb119c00e95a4b3f6731f882a8cc873ffa37f3964b905682712b9bde2040daadce63ed9b23b7e8b67e6a137182ddff97ce33e8ab36cece710a50c8d72be488decd479527ee9915b87525a88349832835ba235adc6d628379d4e1e128ffd2f7f1920e1a46af51be221eb0ab2c27dc3afb5e4ae1b9108633a32ac2684bfaaef95cf2c68944f78f1a8c56b04263a35bcfa1d4728e074dfd93b9fda1e03e31cb7e7ff2178af3e2e7dd1ecd1a154c32a12c00c698757c5a1077f8068f92ffea021c4703a17b3f279d3ad76;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdffe0f8441e26096a5e9cc9734376f62704018022b1737fb61bf96b644bc379e29d59dea15442d5367c5aac384ed0cbdc5452e73f76a721ff6adefcaa03911d83d1e1e4246269eba430f06b2dc2578473d511921fad0d7d29a5082844aca240b88f3512485d07a537912434d17ed67008dcbc8873b354de9a2a242f7464691cecd186750a036c58af9f72d9af395293dbac092b4df1438cf8adbbe302989e5c3c8b912a040d94af23756372fb3bf18134b5a71678f0038de5692dc9e21da378d41dc1e23241a041d223db6da8f884adcfee66d101277395b0abadd04deefa1dea0c06e9c183d1af9ddc3400aaf2cd72176c8d6ffb2728cacf65715c343d18766836c58daf294f2a648e968da9b51507f9b259b116f62d97e56b834c5c30d75f00106f3b424e2469e6dd30206ffcf946cfe1d7ae21846d0088e0e8ded7a23e2657ee802b6129f1a36ad1deab09378a14177858315f5c62456dc417990910853436022772bd80c5de31408dd7f77f8562c8aa29c1984960f2599c7e5ea493c17066d3dc22ba9cae6389f9afd4cbc69717b3abbf165151dcebaa6b9edd7149b321b62d653fcf1f2e3c53be12309be6b940c8f46bda09783bbc42f2543b3c43ccb0f20097bda331b5a402e59de5a20bcb2c482187999457e59d4a11d28bd7130ed25bbdc7baa5855049637a036908ba764780c14d33df9e95ba0072ad1f927e99e901dfa6417ab29568a1a78f5f5bc0edd23964b114f95ba3528242fbf37358d4c430a816072807b1ddd2083bdc7034c2472710389afeda522c10fdf264ad063b1e16cbde43051c59c59e497fa71d9c4fb998bb722e306344a65ad3aece45fc5fc5f7613f322cdfd55ffc450b1ed3dde8e1f292b7c87b35a4c57e14aeed899ba8714951169806e7f5370d22cd077349b321b5811f335df73ccb9997b1b10c4880e5ad6be2b8756a82d5a717dc679c3f85df4a88b03835cb56700da7d692fc3d8b569f193f72104acfe252529cd96b3724f4025e80941e72a915cacdbba12d45862568fd165ead914b76cf5fd74630adc9b72fe377cd472a3fd75de3d76a4ec07e2560f35d8ce1d60b57b6c7e8c6706bddc5ee289e3ad99de8d45e78cb383445552aa49de2babbbfbe4e98aecf8b5840e5c78aff4cfd7495d12e576c32ee388c826baf9f729a1e4bc8d7b8cf62320056cd5dfe370b2d23cb6bbcb7d6618736d04772ad4892d939d638ee77cf1858b3261e0fd2aa210a75f11757fa6c8e4306b0c31821304a96fad9bd74e65485f4041d30d52c8031a5a264a0915e43f610709f6a0d57f7c25465487d848d657eefbbaa0246978d9fb51652fb8d517f57c976f05bb32a85784d715c9f46cbbd2a61be089ba4e71b66cd03f696733f11e688395c82e034e1ecf0f63f957e596e1a4fd67d3d06cc49240c40ded2efe3e28522752a88362019ac11b5b786b83e9dff7438f216a5462bdb75ace99af1980046531f225bc8ed82fc69e55c11f572b92a2dbb36a6f75c7c24f09678f12dfd699fab63256616f381783c6d4c031681a8bbebaf20ac659f6d67388098002e08ae4f4529f842df58e694d096aaa3184677f23fa988ce46708f554c3271702f5a96f034535ef1725de982bf97cd9046b2b224ed39ca5a756b7b60a40f3b1999d07697a197a1de6b86881046454c24cf1d918aaf5a348825f8c9b2e700ccbc1ea85259b02434a82f4ad8cc9e132719b2ecb14b990f63f66216b6791004d6c78b59a101d8d104ac5ab37294db223b1b3a222cc0c90eeb404d9fe4405625c5758e037b6112a036be04c4cc5cf44e0290b2465ee08496a42d48668416464a1bfbbbd550a7a77f5671413bc2a564c874bde83bbb1b4612db298c6f788ea67d9d5fc94a3d5c0c83515f17c3ac1a1d7579f49d749f9d3b51b9ad327605866955696d5af23a64ffdd9af00ee4f3b4108fa9ba53d99993f4761de6db1e193c4b264301c7c4d1ac19ccadc69f66090b4bb44be1de9d035bb4125aed9f3f01b97109234d4c4a664f44d769ad7e17fe38b773a7a5e454aabb6aadba7267c48b540195e2b921b0fa6629f619b02fbd86bab754f1dd087fae03ae8a2e8247194dc833029b41c42bbe0582c8f26f3aadffd77dfc351aea0aff117aeff05f720f6befeb287d966426a02cc6292fe0a98fd7ff262eaae03773535c91907c315158296c0dd3eb23e273d3910bbc83a9ceb2a2ac5c4d1a3b5af89b781c0f6ce73168c2f389d4f1e44a4b833191bad954d05b33aa1c042c74948af009f7c2e240fccde8d979d6577f5e50aa89a405ed9f42b16010ac782a61cb4f616df865e98a13b4cbc3c49b355b0ff205460503378576d92556eaa7f8bf51ed4943d9dc2f1ef13f12f376d311e346ff335567fc24bac0df19aeb198b2ec7ada18e2cf7378907ba3c4aba04013d8d04e176cf0a4cd0aa907f483986f9b0478ef963127919836c07256e3cab9b2d0ecfa5ec8cfed359d96b086287986655170635b39e30ee3677e68badc1fd510454945b0b6eea5205e323d24325b73ce8ee9771b6e37ccc892d1abe76454047497cac3a06f990c2658f8fde204ff9e1d510e8568336edb3cafbbee4e25139822f68a88c0e839bb06bc3510ae4680c160219eba50b3f894e47c735fbe90587b95a8eb061016d23403595802dd887098c30dfa33830624e17fb974cb4502718f5b89c0cc35afb9c1e9296b035192ba0945297e9246cb0606c59d0daf8e03c920d83bf69991533da946bd6e8fcac23f97ca29aa68d9c6fbffbd5814aa764eb57f0ae5825af0dd95d0c1a29e8eb8405dadd3848234cdf321dd70a694da45cad66c40a70500225eb1ef2ce52c661571c31a5d0b371c3107b5d538fcd5782cbb30a23a3b17e94aa758689f8eb91;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5f34a2d82d6e2b2501914a07e0da0f00548db4e9425ab6eec8608e82c9e6b604aa060379454b7d30365afb06726ef7c833185b065a6fe721b9478ef1e0fa9103a4ceab93b4818100b9bf6e51fbdb21a943b0678e501d235d6a2490deb6dfb508b459b2b3a88dc596dbf609e4832a2dc856604917075416e72c3ab5e36685b0080b9dd6c6cf94a535256abffe49876057a651dc0e47f3d449eb17db56e69263832c084b5d654cc9dd101cfde4ac2dcf44c4616e94bda6ae30e9673492234435c0eeb73886cf7eb72ac3e19cf861bb08d9ed2dfeab1712845c097f05a93a3f45895d145e67ae177f76c7f06cf3e4d7d60628e02948fd8d5c7346a08860aef7be3e76b4200e25c73fe622e0650c35413f851b5a8ca75e61b61654a134d9acdce577ba8a498d9843d1a149657808af667aa48b1509ba75eff7945c99e02df3357215aade53e044d9321bfb9ccef7b364a8c6798856067490ae719c6255a475a115558ad6f058455b0e6109d2408a7aeccee0fa3cd71feee7c93068b95879ede1cee5489c446f2d3c7173cf048f785a9b1edd3ad0f607e17afaefcd015582ae2aca99782951112c8a9ce9afa97a0675838bc2bf14734446bc57d55a8f75c23b1a9bba4c7784ce6d4445c840b975089e2e52a1e9835844584e96b725052887fc2c92a923866a3bd1027576946d3957dd3c27720c2ce4d0cc525b0f118035690d476e6d29bf393426cf0fda631d0617e38ac96d8d48615b2e0d00a37c6ac796ce51cbfbbc3f9860b2d8cfc5650d8b94de1b6d0dcc52178eea16d3a45a60d00a067c45bbda63bfb4930bcbc3a6888bd6cfd290d096a1ef5a8fd9c872641740ace819e72e09ad71278e24e4040f926b43d272aa196a0ad85291d7dab07ab37354df62b03ac94276df1f85d335989a67b37e1a02578af672570144c919a9849df66a1e30822fb84ecbcfc13f2c2b423520325014bbc6540a7eb37a39342432bd04c4dad3a5c85de56f8512de464c9079927b0b3cf371f8dba81cbae7e00dbcfe8049d29d08e027585d2d7e532f9523a93402c8904ac1c11fe16b8d422d97ee6877a9983e2b01da09a2e942029e123a40e7b1d7adbb10cc87aac54aa16fbaf5f10b657a44ad8796f509e40f775dddd060ea46fd4e69f21e8f042e4197fa34e448b8b801a8fab3122c039c010b83d505bd08905017ceec3a4a99f6bba40e482732082836e1009184a4241fa3f4f2fa85cb37fada7fc5fe6784f4df213a9cfa716986ec024defdfab78b793e32c5dce544fab519ea31fb8924e52ddf16186665fd41ef5d268af0a1c1a3348fc53c327bbe73b6ad6ba307833e81750324ed6dbe0185881536ffd4a8cd87294eb9fa1afc2fd77a70d6bd5c3f759ea36a569d569a0ede73198b26b2570ee2c1cd2120f4b5dfc132093b5012d6b3209258e38453c1025624057cd52dc5f1b92431e21e96089b20964eb40b71a03224b1afc23da524a3416d719e26619731d0493a04378ee61de733953b22018b2961b8e8bb60f5a1a0af2456330e839bc3b32075badc79b8259a62e0ede7b6347a2f63a5b69e62a32ed9f62b0aff88a4febeccef84606b48cd6603b83363a24e2c2484dc66a7bec49ee8c2c4b968d9f20d354fe229e2aff2d2662defc3c1dad425c5f17ca2273d5431366987b6a68ba3e06064eb9f52e4c753963e3cafb3786906e08a066f2bf9a82bd89cfb4ce13aca3c9695be9396e16d4046426903aa39850a9e21e92f93cd3caa38038d114e55b072a72e82acb81a1f5c686447a2543df35d6b8e9acbf11fc0d2bad798c0fde74a2ff05b7c68bd788da4c8fa5818a03e1b3e99edd50035b4b3b53539132189beee8df00fd74afd55aa90fa684e3510600730ba1aeba2bde8f11324caa3eae015810dc2a2aeaf5197830e22697db1c8e67fc4816c879f060c22228749dcb99d1bc472e94a896098e9e8d44bec063f098b672561f94ea4ba17ad8415fc7d7589d37cbb62383e567efef8e82b49e262a9c02a13e7b579be6d0e5242d100ba069947a97982ddf5036b8efd3e15d09517577a13f5dac0e107ba73a341450338f643a1207c3f29de094566499e3d12e71e5ff620a4119511a6d7f8e6f739f4197987cac2e59c0840143a4981f3e07f6868c16d1f06e292ffe107aa550c286bb9c3f9f18662b303ed14bc4266a0ce46d1ad83e2266744ff36f6fd0538068f766fb01ff2b3d42048486ce65114fce621457ef091036639d8e47002d46ddfaa9018177eaf00934a6238aebd794ed71cbeb0746b3a41e23bd148b604f866af3f3d28a8f073b936e0497f5cdf90c433d31ef3c8e5f4eaa70e7a92c470c239b582fd4b422c0a201c5d305f8036a5329e5ad6e339dcfab9c34d7555378c7991bda92f8bfb08b12c893e43585a8f0490b03fea50dc88fb75952a78233a7a15740a5edcd2cae0dd31fcaaedf05dac02637f6ef48b70b403d59d433f5f44e829a2b6863d15056ef9f0844f906508061762765b1da18da575d1bef40e4a7b76b3585f2e31dce42a1f90f505bf2ce415b7be3b6c239cb9a6e5e28cf10545d69a838cad2db5b774397d56ae7aa7e0e878e9bd36bb0f325723a0176b42442c2d8143b8f5a8df6176b0d76cc88e26012210a578bcf909b50ef59f6c80adb7c9465b9eda6ccb0389c1fdc4b120ec8affeb1a0cecf1079547755d1a00a307fe870ebacc3775027e1bc34c8a495fe5eb9d5213d97fac6b10e5a9d4d959d4a6a4fc014d4db1bce94d46030e62b2c51639b2ef94bd810f83503590cf7d977ca5048d022088b9326d19205c6f60c9c9cca1257caa216244a1ba3ce9847eb41cd1f9525e166961a2be9b317db7ee779fd620e147cb722b215cd2ba6f0de0a4342559504432f4292c6131c84a754;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h86db731831544366e209ccb473648e14988c3ed15c960724ea3271d2862c21af10fb6dc6ffc3a8c30cb905c14775ec906940a26d29337faddaa664edcf501c8b3f66afcf431a4ebf0ce66559866d95aec390d98b43710a9e38a58651134952cc6376477668209933b500968e72af3b3eda12632f6416d60d3fc9d76597890960e4bb8c3dbf62a63058a9690c341a31f73a146966e1e479177d3879f1903871c43a4c622987c627f62694618e51ee320b29da1c651006973b07404fc9355993886a3d1e24c0387264e517ea901ad20652d1df68432268cbc4465b2426a788b97c2ca557152f28f01ba1da6fb6453a2ec2d2faca8667f6e331ecf0968c815a12e5186e2db7175b4a07e4fd82d1e2996b5a94b497f9a15e7ad8c06599ce74c0a61fce4c386f36ee36fec4a11ac42c48eb1484102d20a02b473829e2682e51c779933599db965dbbb2b0f81b9c6a8bd5c35a5fa3199b74670b4a619d6c4475d7ff1109fa5bbc8730cfa756a34187e6feaaafc84271c88c4c149a7a2c80854f654b675c601f98141c23b46e615a683bfe73d1e3affd3a5b55838d085f952b0df8f104920b1d07c519bfef9cb9ec941e16f36d439b1178852ca03a3e340871a52d41f8cd676671a90bbfbfd8f26df0341801ee618ab88249ab5fe0d83bc3530440a65f9c5677108126e074d2e10f6a4d1b8921e5f229fb027b582cd50f4b64ef5fa1f1523dd0f38a62c6fd5de3dff50314f810c211911e1d35a9fa5e665cdb62c469a951c80f64fe110a61a05cdc291c5b70bbd9bb3c6ad623a1ca1054d78c8f80ec8912d19cf88209d8764c54fed5a7cebca94cfcc664233e44d9d3c222b646e1c2ad32e4cfc34019f97cbd6045e6ec96ebf62a7a6e53e2a7c4964b620c10eaec1423f6311867e8d9982e13ea40ebd64c1e6edb428c4fc14d02b984ab6f7d1d6f389a523c692f982c51c15799b8cc1d12a6b8fa040aab76caea6126c9af078f888e96d3f85979c3bf96e49ba3eb939007df9c75b68f03a89c5007b47aa94adb2ae8dde150a3b24d55f79642ac4865f5829fdd61f0657c13a32407864c3cc0db02063cd5828248a4c1f3034bda99ea832dd95e007a1142326331b6400fcda363d0177eaf323f9bb0b1968d91db974906b8df0c628fc82a68b1b5fabe63e72fd66e6b3578c20bb0f8333ccbf8f816a772a5ad1780abc1061aacffaa98c00883c294f2c95f397e43533db0afe65d8933e4853652bdf03725eb9cb9f983d8a521fc8a7ba41376d9df932bc8d28ff9b530cc875736d3e4f8e963424096bca3b60be314282060088674dc7f8af8eaf52d1a9eafc1a145e7feb9db2d50cd13370fce043c7c66645f47a693dae3855a905196bf7829e60e42d65318510091a166392fbf2c7dfef62c9ce25a77cef6655f373bdf5e6d14a51404f9f9236aa15c458c906206fb0492ed618978df694f9c7e83c23b5bd377acbf7fa60a8543c2dfb75e6d21bf294563486b6bccb7874e30d834b0e7ca03c84c789b42ebd6c15286c74d8a6a263a4793ee3c6b40aa0c314c856b371965269fbf9ed029379852d21e17ca437bae6c28301fccaadabfb7c0e171825cfe2a1fad7211af0ba59cf7329cf8f9efa3c456417b4fefad33e26c2f2f62ed8abe72f62077af80098e5e346e8eeba1f8df5a7634d2777ebb3533e137aceabcdbbb8010eed0014e910b18b095d69abbdf6bec37ce0489aaf3587536dd601912a4eeec6be474ea3394acb1ad631a7abe15e938ad60abcb13bcbd1adaf72b7249fe5af43011766594c323c60ff886ddca2ed4dbce3fd9005a9d30df1de7cbf2ea6f62e4161e80e4aed5822de3b41d4eb78b8154072e71298db4b926503dbeef63637af67fc0f7e5d9d23f10fb15392d88b6dcb59e60298598c8ea05106e0a0a9dfc0467f3050177453da2f3f10d2c50f5c86412d2fe3d1c731051383014b5d56ddbf65f00b4e880127b8fcfaf377ff664d3e03a41895a93317a28eec4f68474bfe11eacc2aff178c8d40cf8379a69195b98abc56e4f4544b42da0694adb92c2ee48b70ae683f1397599c0d6702886c247b69d8da34124f290b5fc12f6919d4e72e874154291141b16ba8209e589af882cb889bce95eb2416ca9c773ea6f080abd1de36c2ded714bce558530863ef54dc60a80496685ba832f08fa6d159f926cbcc31b628de011c345d28714d8d268d8585e779de67acc0de3f622024c1303bcdc8d7cd423e0b558e5d8661738ac363f3fb0f54227200a4e8852ff328c3b8fdc164bf55cfb536b522fc634cf7137b5bb06ee39d9be5478a35e74ec1992a37d29f9db033e327bce60fb757e5eedabc12727b0612d7c77935bff2ca5760c5b24d4b597ce06bba7951a2f5dd7cdc662e55c6b3f5c711c0507f6eb9ff49c63b8d17fc11e0a1e4f2af67c31a978c5ebf7ea6c14d8bd62382e92bf726d0e5cc5d420c43cd527898c6321098fe22cc3bed49f785f4e08e8c3e11a0c2b78962f4f4474b3dce8ca1ff7b1aebfc33319054fe332dc0149c0f4f2e1f8f4f1761d9a87b7dd40aaee4677812f47b69bbb625967b8b02d8bba5230400e26f371a89a627d870ee04bbdc85d201fc8f6702545a8ff90574cf37ffb08bf4fed651abd8684051720907434c266434e7990af51d61ee83d49ff436258ca9dfdb1794e3bb0e70ac639c70d6e992444c4d2a413b46177498f3d6bd270106c1d3fd39f33eafc03b636e31e591d925eb8b8441b7d8deda43882f347df52a8ba3ac64a96a8b7efebaa9e8b324e2e47861dc43f2b979677038a000eaa724b91883e55d21a148c8fdfaa8b104a97d742a097db79a8b2cd6026abca706331331f0761e04fe6ca9c3ad6c43f1dba0fc907a5643e9fe042344017ac012dbea31e05862ec1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha7c004226fa45f92bc4ce05167ebc554aac7faad4ea52791ba9aff4b79cc64163ff9dd4e5360dfa677a5daa36b8d58484d571e593852571bc968f3609ba5d252250f57beb5006d6948ca550e1796bad59fc394a9db84b48d27ab6f380b5bda2cebbaee202097255e003bd6e19350eda935d6eb0f753da9d404d2a70852aa2c139c175a95afdea76bded1a7e4a1fd76ec1b5ab4b9cd409716c811ba78d698c2bafca8823aeb6a8a88d0aa387e3c36d470dfc8332cb6982a99b2da2dc980f1bfd74d76674759684a761e9b2164e430deecd609439edc0c9597be9f4bcbaac6470a5cbd41072291c5cabaa1b680a5d24594950eac5e4efb3b41e3e1e3451c1604876dd1bc524662828fba388f290078065da8f5ae4cd75fbf41992510bb8c8116d83bac4cb99074fe18d4d613d1e9eb361fa1af1dbfcdc64367cc7825d6319d4f76533f807625fd938bfc495653af2fd855a2b4d2f9cb35c768f3d19856c3bf105447009466e5e13b07cb2a87f87c1130e40961d987cc1cd720f5fd06349e0418bd48f77ba9b717e688cbe4f5f443f8d0031fddb8d3e6be28f14048ce93622449ec0fd0c113d0fff18fc6b6dbf7f907e376d849aba72d959b9ff76fd32a28bd4d8dd102ab696531f94cdcf4f3c8d4e76541af90d1faa0173edb9bdea8e53c253cfb68986bb75af8ef04b19c5e81ae63db9990a9b99b13dae0188cfde22fd1fd8f21d2e579731bff7974b55185b283e9649e5a5999ced88277d75d53fc64b043babe5e300d72e34aa902ecb6450e6b3c1d4423f634c323aff3a6405efdf972b439114239b35c5398e7af476a6222e57f97ad9a9e10150db36afddc60057d098e75d874a1d85cd467d563b410c43491f0ce7f132159f0ca46adbdcbe7937159f36d917917e519c83ce1f3c5eecc61b83c4ea8ba5fcdbd38608eade403b432e7c0679c31a4da78cc7bf0384d3253de108fa5a7591bca48c9fac0745b23d6c4e1b44c7e12bc5d1ce280ef3821a55aafaa827caf8bae46879358301dfdd01681b2dacd42fa009f84acc82de710dc9885d098c211454c1f63eb9e95e699eb347b3f80c7d9d6167012a07864f0d9abfacfbc4e8fe310921c02a932475caa5856e30570e58e26e4c93e19c5dfb17cc3d76a57e9de38ebc964919dd9c95a528beb211f5fdcfde35a9b37bd7101bc2cb1750ed370850629f57f986c3a4978ca27f34e210da3c28060c1e4e6ac3d74299d7ff0403a29fc1d29dbce50e9fac07fad501149dbe7d08d41c7dca73922745cd8657448cdb0fb0cac5dd017ed66c37efe976f6783420c905c315d1216872ab04fe9b9343b9981177c79e07caa0c5811f8e80a0acd1f0f5917726c59f5cc2d6b10d86f12b20ffa3cf95613afa2d2bba2dc97f5eca0bedcb4093ad9fdd8236e21061ded489ee7cd6a55de2a9393e2fb085c2d4f046ec3b392836ed50afae799f793f92bde563937f9c39083e7e52aa4ac46ea474d7a15e1dfee27522af4d7f9e22b1139b20cbbc3de7d8f5c823c72710d027c1925518e15de7b46f0fd9c3b025c7a089fa0fdfd7b2fa4ad0977b573e81f74a5f69a795e7c4d4835993a2b3ee366c88681760f09a7afb72010b70bf75acdbc42c6c9b3f161264f95b790e3425d6dea6374492efffa483b444a665671b58805b6e7167f22835084a9bd22bc085896767284d5cfe6726d8a3603902e44616779bb9b9a41d3a63ca3094b779365326ebdf6a65ec1d509d13310317bc6d3e2ca8e590197666a01ad5f0a43b033aa422945a1b9a773e29462d55e98d17cfa3693c5e630b143b7f9a4c9639421a75b08d828eb92094304888f81e10202c64588b06e884a929acf38a39beb900c1893d8e386f52d350a33f2c701e0985cdb7620d85a9370fe96055aa5a6a9baaee74be92a870754860e09442ed0bc939b4edc7391b8754482a3ba6d0d74fdb39c96a23f431cff1c96db2577b5f66da752c9ee966be98d01306f4faf5070a685a8fc4cca1d9cb0c5634d47bcb24b6d1aade539e2fd009a3d9c6990f37d260eced8cec13839a17b1114b7e7f9eaef9de719a0ce16246996c2a8eaa1340b56365f44fb49661fd14914c72c41c326702520da756b581bdfa646775aaff536097c7ff1bd1a433c6400d300a6ce0876381fe2471e2e3d6c9a100d78cd4df35e338d634c3b3c56d8471cdfa454edae54c9769a35cadafe96694e13c02ecd2b8b7e61c928840d148244c40c8427164ffd3ef0fdee04c4bc34938ffebeef5329b6c9a6a94deea17f13e675ecd0d04fe18c2035004cdc7583e80916c1279e536522b16ea6325a280872ed6abb03c49fa59c157a47dbcf90bbea6f6b154b6f22c5fd044df9f990f09e9307a81be42fd355d1279acccf6b5a7f6352c5cdd146a6611907eabe02970e47f7464bf469f7c229fcc8e55fd3d2a23692cc8b056226eead8a66996da817cebe440e6d64523f1a42d9891474117ebd2f28ff7549eb2d95fd7277e72a29a50b44cd537a72ed2a1785eede36b15b00b0dd50fca33c804211d44147cfe986c4b9ac8e22626de46ccaaee97c0ed65b42ad2d4f97dbe48c5cb6c466904ac6b6cf5edd484d01f0908f656a92c8cd36af7161bc2e02d79bc57e08a4ec9e92ffe683ae179f39cbc768edaa1eead3b0b1b74639bd6bcbf2759ac771453a204ff04951303ccf7153c52549660fb42ad49bef0e33b08eb37ced666513d6a5b62f86e500b0a526b38f83d37296b4fdcb465e422b7007c82717c5bcf2290c8572751b790307b14a1eab5c3ec6b4f70eea3acc9cadbc4b63b45176efb9b4dc99c2b0a2199683a4a1da371122ab43e02ff88a715f2c685e72db7627ed7fc90804c3c9293cfd7a3ee73353558cc05fa322d3f6b8e0d9fd7db0065b80d82d1701;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha8077ae961632597aa9706c21d1a3c1d652d8526796b61e0bab03d5cee4e9039ec13ed9d99e5f462493f04efbaeb5bc902fe181741f680e54318aae262007903010a1837cd0a5704592eadbf0b35349a9289dc007e58113a3026198b7b3b4b5f699cc44e719e27b0ebb9096ce4949259b835c104f595e765b0d79cf161821f4e6019d4674da6eb738fe484d99c2be151d74173a6454233afc5acfc0b785efc54eca978992938129bb88ceee8fa496abe19aa76c87ae2a330df9fca31fd7027c49d4d9604de56f7272c95475b9bfe955f3e5e896b1f9e7b0c5ef32bb7590722e6d831496fe5606830f77d1ffd43c24b21b96ba97f4a0799ec1e0cae63e8d832e2374455a40de544deb72c8a54543a163f4f078b4fd2437fbc6de67f25bf045ea4f3451baba87188957749e2418f1695338677c04943a21d01e6d3c55aca87762df3674c087a10c2e79edaada117fd18c4ed48d1e0f618589465d59083938d5baec038ed57e604cb06925251cd5eb8a2a8f87039cced56043f49667c6000beb9e5ab9f1a7414802fbaf50955c83b3c5d6d62eeca89a8eee839c204925572e49cc77206960267bbb54b2b2d4a30e7e11d4e7ef11f9c1a7e7b65893f630f3b1e30fa207ecdf18d1badcb80db7f18bf5e5fef391c3f7fafbe96e383986192016bd0a3c0a488898d5a28651ab78fee5ee37802f62799fbb20b0c6ffb47be39f9bdcfcbdd1850f19255f2b4ef52b063452d9b3a9f11522b26e15fbdddc5fd71679458e421f52b37941e4d3058c99da9b0c95f4602011412bc824ebd2039a0e80a34f0ea0d017db28b51f0bc97ff01433ae265db395d4e89b2515591b55c135fcef60f6f76e51c0d466c2c62a044ce53410c074edd90b18093f14d1546a943a6a8042b7ae1f2706ebf71e1878147652648b2eabea0560de621bd3dd67208b36741c00e820b213127141ede0be8f091fb6ac20ea242b094d993c91895c25abd1c448e2fa120596927234b2606cc590c9aeedfa0066ea03fc99d4c54c457bfc5debff9ef082f997e46478a7d1db1b1d3c649441063d89e99c495afb0e23e384d73f065b1a314b13970c4128b5d5bf3838eb3aa92849810670db828e124cc35d9a6d17ceac126a8f2cad90cd0f4abaa4be45ff3ae3c875ecba95d042332f497f0e6990b532abce84d768e73b932f2524e4db02549340f69c5d9ee3de74ee0466f081e0127e5f57e785f6d125b765e366a94a8681a90bc8b3766738437c24df921d28d95f1104679d9ada78b8350f14fcbf24126ab996eca3865a6a4221a77bad6b5ecdd0d296713070b0f98bdd0dc2ff707711a89560e1ce1ac574f7ffbd54e853427c6c4e318674ec104d5ecc07a2c34ffdcdf5e831293e8cdf7a98532ff30f69eb1edec634d2a739d21248e677f87374bee835c11a866f3199ede24cabfa5b87d96acdd73b663b49dfee39ce385f6aab54f620587325e5e1aa033ff0cbe503562815823dc8fb43fa2eb8815122baecd6916806661050b6e8abae151c9aa11475c800bbd7181ef1d7b5e8edda0edf02572942e2498c6141581df360654ad72594b335fb0268ef966c695bb75397fa5b31d75493d615a9371fac4148926fb91186fa7897f47c346df371ce59417bb4a8acacb648baa5ae49a9ee4932bebbae9f70e6a23cfac2a549e377ca850400557bfdc288264e00399af952668e78b6bc86f67b0d07a708d1cad3c5273e36a11fa77326f02c251b1f6b842922cc997a13dffcafe91ef4d6fa31282d2c06d9c4615c909ea8431cb36f0b9d26aeedb28d6cfc91c48efe546c77f4e9d895f0ed602694746919f7ebc7cdd90b81ebbb3dd1c292e91577ba5346402f76f1d50937b5c24a3ccfacc0513f7a8d1869e106a8108da312f4142ef7bcf9d2e64c2a0beaa7fbb3f6774c603a2573f0811df72bbb41ebc9ecaedb7f6bd8dc87f1ab62f8a0b5a16eea949da0ff71238db4b144e033ca1294fe7dac018977ddff41d832166b66b2cbe56d2db383bc89bd29023c6cc5b25e97a2369c1060a7ee0ccdf9f25fd5645a3580000f12c5724c48bb5bda17bde582b6f7218a4a424449aa7873fd19dc4ea87db40bc29125459ee8d474731ad0a577e65ef0b45b1a8a51faada8c73d6adc511f178b1accdbd5dabf14537843efebe45073e69f491c9a3d75abcedd5a5d81be8c63797fd260151e169c3f33c4dc681f236d5ebc15083a26d73c98c5532c9a211a0349ae36c8230df8683b3ab51c18ad0439bfa354ce8eb4785a492b9a4d31985f1af28bf1b8accac4870c9ddcae9602709ca54860cc769d28632ef3b51ddc248cc748c55700f8ea74c91e0ecfc5f077f1e563321ece75ae00af12d6727546caabe25313cd07199d8fe7df1edc7b10d8434e4d06ce3d6f8c3c94bdbaea677f4e634a72b0dacf2d38654f37a1f7f4ace0b58e54a71805f660f985443fc576ac608ced7d6857384765802accbc219b3e7e9587e8573ed93a12843e793597f77bfee4142fcf51c55cc906359f506fc63cfaeabc7e0c3379234bf1554d74dbbd375b2ef5b24221f41b5b052283858ad1eab5ee066b9b9034acdd7e82cdcabce220167b65e1c9779ff6bddadaa35415ee25db58470b453395ba81505441551a1de01993966ba48243e2f4f2afce58f9b5225039b875d921d1593d39f1291bd2df95de48fa5e800a060768fcd7032f56d14ee044775bd2de5fe6d97093b00e0c44bf89c6a09b0d6db95d87591410aa5b3a4e3819693980b3eb65fb5f8e99fc0d3111651f9bc734009cecad56c94119f265b2257f14248d4dfd1ac101b25d80443ef1272fa92137054891bc81511a4b536dd6c2a0c7c155b50fca3d7a2b8fa3e954cdc33813b7bffae033189bfec215015e2ba89b5027b33dbd5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3352c5e1671d8dbb193d1de71f27e05eef33443bcd23cffb8dbf642c37dd047b822350b8908ca94282e78412e5a0be9b374350fc8a5deeeb2117e28a43044c64177d3a6f6cd6a374761b6830b0cbde0684d7e5b6e5465be86746d7b9ad2517ba9e83f59942d0001e71706973b8fdb6834206b1e6fdbcc8e9ea8b343b6329142c8dc3e7956208f00b76761f3937738b0b8df2218c31601a46db9d94f15ef52b2de89efa19e12ff4926a09997c3b2dbd013a14ba7af2d320c48dd7e4c1a1a96fa57395642a41d5d9ed5532a554b25643f1add00b1d8abe1e3f54927327f1f4f780e6f4ecd691acbc9badcfd1f03bac6cc95db6188f44a287c38979dc670dfa0f198cf6e77742b6ca4c8b2bf96c554db4a8d0eb1b170ad3f178d021bd7714196808a0ea99b84b285b49498c1445fe1cdf0d0c0572728b950ca75d14d7ce6ed6cbd43b92b3ac45048d3441b6683550c840af33a950da0f446e4cd4274eadc8884bdc42337b9779de6dc3d9e52a117cfbf0a95e9ffd8e9857be5df2fc3927ac93010d56d30502a241411fefcfea8cfff0b06a293870e82acf0008e17b2fd3094a531a774bd0029de616bf929b653e4d1ca8537fe2feb8f20af12031559f3ebd92e028c0a38dd3d8114b98237d5b54f35ee0ed3d33206151c187e292cbaccd41b8ef1acb484d1ccfe180f849486d4fd8cb63c73178bc12f3acb90f4cffcb4ec2c997a980a8974f8a18dd1472212a0aa45d281aefe075475cb39bed3de92d2b46d19b96a8b7264443fc952ddb476565fc182b852da9e6425dc810782d776c2a104ef446c405be1720d101aa936bf04ae09841ba734fbf56be6f4e35cdb1980ea33d56c7040f3636062b0cb78f27d28532d90455d6d5a60538d123abc28c67d581601051f9f3c7ad3287aca1b16a5545383823d31e4a20d1ef37bba3ff0609cf67966875604775f2eabfa9b3090d177dade1a29dac25563eb41c6d6a0a508aa02490be9fb43f60dd7320d783fd45b1eaa6dd496e41c7ff8dc8bb166b2165ca4e19b061dd2bf2879a24531a9d47eec298cf6a78f0614ae59693bca45d6b6a0a90b368f61312dc2d3e7ca3e066ce11cdc4a629d6ce2cb2233f97db8126bb6b1ab2799e3de7b91df574d0f7488a37345fa641c4ab67fefeb605c0710c803555fd055c06d8ec7d2725022a8e2faaeabd7a847d2719d59d39fc73b2b4ecaea6719d1be0f5c6b519b1e2a304930fcd7f2aa6318043519a47f9abb2637098c9c89fa1937b3ddc2bcb0a2dd017139524ed85bb0d125b798a34a468fdd971e56a30e99d7883bead5ca0916b36343c3bbb319d8002e8d5b2312a3a0d4e9ecf7ef703fe923e3ac7f77fa11bf99771e3ee027eba8f4348a4a73c99bbe392271394ffd3b1841603ffd7137307d43a99b71b306d687ab816255e843532012722a0dcaf6826d3732cc95a337de212493ca88a8fb99d04bb9c5308cc35ab2d1b55d7faac578c163bb1997454ef8b399c3cba4e632f5b83e86f7d4ba8c3b58a70624765ffc1587261e0ffef7c3cc79e315d57c1a7e9c058b6b558e7a7057e69c3622302b1c58134d835f0bc96ed2bbb8ed9400c3edc43c5c9b93b599529c1b9c8e05fee789ac2ac67e3a137981438a60d5127dac2e989bcd61606c78280e4c60886bdabd40a1656dee16ee4ce8ab6a3982bc0a29e89a7039002e4b3b92b06197c97e6b2ccea9ba6ce70a03c3a33578538cb609dc2a50332445acdd2d5eb4a0d97152ba9c39b3ac6a1814f017fcb1596a8ef7ba4297b41bc5168c3f2ee62781dd37b966c15f9d3543d900d76b595a95742d2401765ca50c5923b3f40d5043fc2258e2419125a6e0235c2c1d6965577f9f18e7989e3d604aea6fa3c40a1f4c868d0a75535b25e03dd58306fa525b41311fb0df96cde2039d43ea87739e630001f57db2b78d93c986fab0c14046842a35975e2945e907359124419b26b4744dfe71923bb22f3e483935b6547a861e9ef84d603792b04424a12592fee30b5ee5ab4db97b2c483cd86c19cf18729ffaa6ce7a560414d8c2dd53b09f1abdd42a69412bf0099413dd05e74f1b436d738d1649b8a9b15f4f1ed2b9c503d44f7aa1e3d1e55488c9c599fab3bb4b138e818861ee9bb629e1377d01e45bb1d77d06f1c4dd3e7c5d299a45514928f8623494e3f95b9453edc2f87ddad29127dd84e2053a3a148f1c8b2c7d5aecbc915ce735a83c29827472d8f62cd239cbcc8e84cd27ffcd8da49960e191bee9b356d4f10f10157efb226b3bd2087599ce00675267237c702bec282c883c91fa8e72a57e506ca44fc52dd50e6acf9edb59faee81426fca5c6ae1092b04795543b36f3f8827f91e98569fe7ecb53f3631b32d8442cc807f663a46118403ebf2a5daa9ffa92a36ada00f7047b78f9d8dd95d413ee355a33dd9d7d1587238a03ae9d7466aa6c63321c20d877c7df40f10e08f175a6635671b958b935e20c3a0f976ce074ca8fa82796cc7856e9f731e18d190eafa566f18ec1b12e5496441a299eeae894978e972258a08f1fb0c7bd2f75a702b7d5d2574a40aba8ee8b28d79327a4405fdfc96366291ac0dacfbd7d5afc56c9932fa59d345f6d782ee9eec21948e6532f6089d8d670b588a49dfab7df4963c0f188123e26bdd263782ee5ea9d092ef54b70e45e21dfc4b15ac68088dc486d0a89bd2cc23967d2487ce0a142dcc11f333682703cb6e7276ffcc64e6fa2cd068805325641770b0d38cb4e70b0cfb9414b7481231f612c67eefb408531b71d46fbc9805ac117640b90a0a0120f277d46864f6d6ac247298c6d29caf85a95ac82ee5f9f97221eafab1b08391d1134983a527d1e848e3eb3328b53179eddbf7b15be7d5cd1676bbb2f272d8d42dab1313026f99429d3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5cea786c9f66f276c234129c8b85dc7b6db1e10547fe49f71a26e97d2481f063e179807a8c28d2aefdd21fcc70c14117a0c638ff3ba6e6eb6a2d0c246bdff3d2336e044a6a5b11fee6b4929e3cc9af22db683ecc22ee409819458570f2e821e37a3cac0ba5ef3d67df91645d64377535cd4462d90fbc4c0a68d8a2dcf8a2cb14827003a3ef7f0d8ab19f5c458a00f8f2c32b2d906135571d03680b017e0c7f444c61ff3a8d430157777739c8c7615be62da010ad7946c8e5f075f7be1ddbd07add88385fa80376d4716b986df7c28e0fe3cab8a8311db38e002fa2b254f1225b709879521dd701502e1a29dd7e7750f4160d90977a7d72ab1bb80a3a65d3048f2f73907ada70f5d91ae8c2219b7e60a413cb16df493722d321ae63261260583e0c2e1f40ab89d60e2ac2e6a132fd4788d6ef2b33191bfc5dbb8c597cd442fc4a1c1ae33538a956136e6d6ac0a9c1864b1a78c92820cd27c71d3280d71f17a8e3b8d86bfe24daff5ed3093ca482f9ff85476eb65b6674dd7447a8008d83336fd40481160e7f76b5a406a08202d97fe647a2003cad43f036c77c2f41d239ef08829b8e1095b670dc9a32739f3193d4fa885600997ab0ed35e1371417def9d8de500a90ce860a67aa0e541f02a29474c5d30c0863779366e5d03bb3e16eb5b082f9e202822d1c4bce89cb9c4ea22faca5459894784369ee549f7d708c47f0957ee973e63bdd5379be4f6c541dd4df252a59cbe6dab5fd00cfb79c23d6f48dc1f2f4705164be0a5079e54b7eb415745454b2abcebd4ab402f816776d2c7d611cbf5f981f1e8812ecd94b72f7455db4882c1fdc48fd392608935d6e323ff5a7d0c3aa69902739dbf76b6281fe7fb025a77f5dfa08aa41551357654f959cb11388cb29ede49944893bbc20ee50e63793e5c4881f24dca3ad685540d10183be3eefb8f44bdbf08402ca369cd799b599b8355de5565c6dbb3259f3cc7982c49418cf007a4a9d0ec88d98470d399541cd6cea69f36cbc559098af481d0eaa2c8eb5c1911a77a26ff58b88da813e980e9f15b5299c345a79de1a6bfc7fc2456deef367d3cfffa5c5d92d16b9948950c11a54ccd2beef77ec88a4ecb32fec738d436f6837037644c9355d1d966117140fd6013432a0e83dd3132abd0103e3425fe1175b4af69297168d6440650ff532351129ec3e8dbfc11e614eaf58eaf0c854932b6f7f150d190dfa2a5912acf4707e5e28f2bf4a0d2871cdd6c2939517e0473f9c51bd94a30494f95eba8982bc69461c7830c02f878b17a22a3c7fea8fa206bc32e8ca9fbba7147caa243bab683d4e058c74b78f63541e82968a9e341786140f54f28a7515e1cf8959279c89158702ff6328156a7243a0b53a465219128bbffb029f6639c6d99853bac2870e3fac11db30dc1bdb15eddcf6c458dcdb68954074534a8180a5d86c127ca1cc1fdf995496750ef007e4f542020f6d24bb8688cfd6181ad514bf5e39492bd944e69dd29ee4f344888b3b50469e22720f1ae2e3b958988a9441ed4871573803607b2fd40ff645936862b3ab487abc0c039ca7294a356b2f1697e7b110c2f9daffaeed8bd5b241da6f85f927b1ed2ccbc758e98df98472c64ebac786c06777edc2745943c7947f7ccd633774d9856c190df41a8c55bde82fe3bb30fa4dc50e5d376d0a332801dff9ef7e4f6590ad40d8e3147de34882def038455e748093c03d9d3bb45f5ddd8af00b63bd070a5ccc2916d5dff4e0a894d5d0ea787d4a0084bd967dd4667c57c87a20ab593244adbbe1a7c7747d71bf7a2b7db6faf1e25ee59ed51411ab2575e588172d04794098bfe101b79c3f509af98177d11141516cc694efa20f4290a1fc6807a6e397c3ee3ff27ff635a09968e7c4607f4f2cd25444c3c70d9e5da2fba1d595c4846f84b768c393d539f2cb8bb0e3957bb0d416b2bc5b5237c1eaeebd3c81f8e515c513baad88b22e921069398c69820e89afa98d2c4a3ea05369abb4c50e9a0e474ee36c964d9ffadebf1acb2f32b2b64ef809cac1ec8b3038be7df63042450e352ee4cc81bcab51d910940de912e58cc81b2bd6272e06985cba2ebcaf6dfe2060800d10c30fd6b2dedd3d1815b16f29f000907a48e44f71fea5765b40fd8dc76cf2337379fedd0ffeeccd207f4a428e6fe8cc2089d7a066437838224b0dbc25d0a43126fd04bf2be28a0f2affa5e460e8d23d1674866ed80968144922b8d1497d6a09014102b41400de7768137e44960d381339427e7fb7e209ec3ccc3b7fca6bd1706ee36e937bbf346fc8f4f248907cdbe588c7fc418339e94bed10f2bd856da0880164e9e090163e64c9802d987f5aae2087256b10bb8f21ea04fed5c6f81f0aa19a3b7070244f1ac74660e2d6a6fe648b77a94ff6eec5e81eee54af5d31dbacbb120a3036a01f46a707a302c595f28423ab296f1e8c93abbbfb946b471f57b43860e4f680749a768b98ca0fec583879339b022fc13f4b84abeb26df24dc3bd73915ffd776a8c36eb89a42594642ca10777f97ec354de937c27786834cf43d6a0869ca100d743d71dbe6b83e2f1e2e747e8c8568ad2c8ebb66422ada012538a0b0b51d4c77be9ea47828e1114893a499cce5418f265389b80d69a7560ad96eb7d0bcaaf3fb3478752799a611514d9c7a37b1e18260960430bbaca687e47a886bb1a28ded165435d1d5562f95821f01355514680ecc169cd5a363941e79903c1d8c6a156565006fb112b2fb8cd2d14691567932e01aa10dad5e8d44db494e6b302377f3f5393abeb5ea1fc56df986b5aa58bcf5c86be8c362379a81058c68bef1c424979907fc3b66be8e506bc3f6922aa07788ff265954cc537587a45f16f9bdece329adad10cfd15e5a2a292fd4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb73618f04a8fd551a3195fb1571da6151f50bcfe98b7cd852c81f252de0ecf7b5389c68bfdf8d8d69402db0da09acbfbcb04ca4b59e24bd33f420993d584027b0ca5c4f30d21cd035a12f8a708df9739d8487b30821309fd594690050468415886cf53ca8cd6dbcd264a5acec74e8ee2bf5336bba66b65e91392c5a11fd02201c0cabdaa249b120d58f67445a2f719d9be495125ca9f9cbed021455178ecee5d6473023d00e2d9e0593d946b49f64bcb3c236e371c8ec36e9e586d0be438c55cb446945f5bb2fdcf9eb6608810c3f0a2c12aaca54ca964310c2b7256ef3356cec875c500202eeeb3db0b0b1ddb8a00ba36c92e8a23b504da887f1c962bda959f81d49e146075f87672ac01cdd7b1442d47ae3f714840dff78afef0c14e47fb3369b9e0872b9fef695eb15c400bfa8f29a35d56c7e118ae549eaac7d2610f7b6ef0ba1676192bca84b4d73747312a4440ba835ad24e3324726086cd6f27646e86d405944ea1e27c21397c74fe5d85cafeaba3e24ed5a2ea9db988bb943d97b3699d57c1f47345e4e3b736f4de0f798568613cb40edebda1f9e7c6a84016a11fd0015b232e11cf1cf114a423ca4b1457c2e07f79aecf2cc50c62e249dda66b2ac96805a58a27897fa3a838871cb98ab94ba8ebe7d0e9ca0f0be265a4134bb504946fa619b12864c982ebb1a1f25e95d8a18369bb20e711307c57cec64174d8d9469d119cce075cfbe543b355fb9da46958fd964d846f2bbf6835d309615ba14350dc6417d17b344a5d02f1787b69a805fa541546f43a0f7d4bcb096ec484ef1a655b438f2df7479c4a912d55b82d259d1b5b4b2d106aaff417c746ae0033a4f1940f444ebd1e4df64749acccd611229360c9242b611784700f724285ad16fd817f199ad602fe367f1b96f07fd8ca8da24324a4ad81db0d1602f86046bf96e2b59e72582d66a33a11a20e617b78db1e6ad35191c8d62106606ee25b2bacb4596fa4c60b6b1bfbb1e97f881b86b48e1b099a0924f2f73f70336053502ae4a311ed50d7895ad09952f5698a7c24dbe20b1680f6e0f93e22cdc7d94e240b52043f65f6502185b853b322743721c046ab80d846dbbdf323ce10088c2cc24a7c2dc37d1d0a7efc053dd7fe20a9679251adb85076d694fb701f047c54fd575bda3b72123186cf9a6ad3b52e481ffe1cbe25a4cd08a2d626a0603a36eb5514ea852e79cd5d603e4b46b6a8f3a366c99b14f9483377f61f3f10423aa846aaae9448a3fe60ef5b6719986645bec9a19e8cad5a77ff74ea2430db294040ade8539178c5bfe3637f00aa17c56ccb100fbe775412b362d609f7d9e3a5db82860f2220c49757eb77f1368c9d972f9c26b9b9eacbf0672f13e2e5a4089448f68d03f00579c1941bd538dccbc35d43436ec93ce9b1f6780491824c84408b1d285f0c57b73cc9269573237f9599ac5fc70fb0917964ccb4eb83aeb80847efc055691c884d520aaba781f6f51ad39d3b9fda4526ff49e5dd910c1994954554ca69fa89388b04ace7687fc86797fc8a9d422bcddd0ebf83e227828bafaf0532430e5f1ed20cc6e689c459c1c680e18bd5546b21939db49c506366d8c5f6fe43ebe22398b5ed97d4a8dd7649e755988baccd019ef1ca08f53044814f8f85c8d374d6cf460c1b82b9a13db4ddee7c4f319323778fb0b66a2d230c1b83b0ae3c920cbf19211c8a8dcfa7d4a1a7acc8e4667a5fab8b6342ddbf1aa6f32de1a70103e41f9f01dc9af50eed612c203fc303c1ef4b932273ef6ca849e5a9d843808fdb4bf952a3fe645276e2c9839e91bb3a82ef39327bc8ef904f8048ca90b8a513ab8fe2b200766ecb61df62db868e884d72771131cbfc36821438677844223ff05f9ed4e61d3f4b9c2f868cdf4f918204ccb3ea7abb6d48a3b9694f715dd821a9eb026285cf11d110fe16625e7e6dd7f3d6bf1b26c33d0d063a62f668fd3219f515848a4d5bb218fbc781824c91f4c156b8bf132e3df88fb247cae994a210f8607d5d89c09d39ff7c97846760254c40f5950240e25acc33d6235f36de48e3becd6489bacfdbb7e814006bb6f31f799b7435d04915879d20d39f8ba89f6aab8d329785bbab0780469286c781f740911021bde761ccf1362ea2e10e0212b15ccd129c0f55475e88f00517ab84d8229f83022de2981a0a7a626ee7812685fc1cf41b657d538846753ea30f868b5ba35d0cb00684c914498c2e297c472d1e8b4c7dcc7ea262a48d8c31b0252d237730b017924252ee8d5da6fe891ff39e5841819ba8e1c69c682442c37b2bad247184c5d86ec24938f5ede795e7663e76499048baa81b96d7ef97a064368435717e64dc46c74ea3144d4c82f252417df638665694c64b6cabb9a1e7f7ea37464645ffe59608845148291ade4221270c19fd37525ae30e5f876bbe922626a813b6a9bf7b017ebf46d8570af69f304e7b59d6fb39ed85b5ad4dac2730e2315b2658b369c89ae0104a2fe23dbf33473a133568c0b8b33e74e9f2ebebdf1be427cc94e0cb74cb62483678b2481206d2d460da57c7afd659ddacc35746b91da033a1e944878a8297423a86897b9657c294be77d294aa0ded2facf768e1b067899b93d7406041d9c1ee773650d0da74668b3d3f6ddf4b82057972ddc81d70b1ca5f9fa828c70aac3d5daa0f8ba9a7820e6cefb17fa34d2ba92e0c13df47442a1a6c78a50764fac353a16a98dd1b4b348e51878bfc0c6f51464b2c890b78a0301ef48cda5ef81427d4384f6de2c1ea3647562c7b9a6081a69e2a3e1bc113d846c56a5b4e262bbccd734ae5f11231a8403e333d656d993abc2f465dda82b29f374f1ae3082a2f9e2610779ab671a82d9caee7eda1b7ee2341c4a2f998ed53a44b5bf64441c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h96dc1776c3a44e619cfd6feb3c331018a1763e4040ab80841c3f2b12d125466af3563fcfbbabc548a11206d882e976586fe6fddc428c2d42a8504c5ef247ad60f8897672d1159e2d696125b904ee0f651a3118ef077d6e2127766da1a0567802b4e3f859d7930658c6c7045d68fc0a87727b42bbb1084c5982feb6551f8d05bce57ffa060396b55f8fd65186d014d586f369ee5a3e570356fa59ece87709d906ecd8794457b7c9444f7e13efefcad3aa15d03ad6187d1cdfc688c6c4addeec046118f0ab223e411b4e9977dc85b6c8f425c36cf5f270a4a37b1fe5f1163bb999ea90f3e220fd9ee08edba9dbef9b20740e2397f826f3c9b443d17db7d983f60389b58a70c4d0e752a60c08e3dd61abb985d41ae0de47ac6331ea7cc75ae53f09402b90824339192c8ef6cb818a43b80d802b712ba0f5e038875ddb75dbb7067a79f7bb8c7421c05af76f6712375261c4431485e3098e97b81e79f29cdb4c0dffc9a50ffe8f41a169ca159bfb956442846d2ea433cbed5f93131e68908ab7c45d6ef424138566526a4b8a9d18014667830ab3d005ca2e1f14caabb7d7adf15893348bd9d6d0d9217ec708e476bb4f3713de1232746564cf4d87c302ce10c15364dd324cf35eda703ee05417fd295edbc5011a428eef2bdf71038213b068b55cd4329b19152b5736d9eec5a090a68ad90b966a707f2b0fec8225dc1c049926bb3cc7e5a4293ae92f2e4135d43bcde8973108756118f9a75e2b70292ffc6b0e7f356cbfbe1d23ccd15ae71a47d98a6feedb13fc59d992d7f73d71a3a1e046c252e03be878bc6fc2bdbe25d53da6b403947bc5465760823a8ed1663be2c045e3be5d6e085eebf12f093e0dbf7e34070f3ddfa71de4bd2213d0f97c0954348974f631388d49f1668c7e72b1e594ea4c7040f9062e985b5ab7ef4db55fdec8e4c375b0bccab4ed0e0c1074082a253ebf3244f067801d2fbd84e3fac44fe0b90e9304ed25d267be2185624f30d12e20d0980ae2e25b9f8d759e99b9941f7c7fde21a98d194a5727f60baef6062d737e0734f31b51a20c3da927f0491c4d7e86bb979c56e493364880b478c2217cd2c7c2db5c7077e47fb60876f0c491c54266564240587c02ceed153ace19c684581b8b3be91a4e9a8817319e102458df49078df1cb2d64e05d1a03ce80346525fef2c786f0c4ffdc074a122d60fa605e09178a5ef2c7ed086fcc21608661377b550f12ce6c1810499bf7c33f6f8547b606d0ba6f590af0ade584fffdb00f8835000bae7bb221c0f00e12bfe9fda779f047d11988e197ee8699107836a0cf9fa57717c071dec6b7de056358fe6dbe8948deccb056987a6174b728c2dc2d9afcf9212b62d5144edc7a5e0e13b00d10fe0786de58e8f7a44c0399f0ef8942c7374ff6adccea44d88ffe3767a1d0051d928d0a5a52abbc887a77d72d4cad6e044ad14c17c9ad0dfdf705bb7bf6cacc48748674b9c8585623e477562df444bafe9a5376ff141d2ba2cbe28cadfbadee0baac87860fb922a0e11bad0e7e66cd6e58cb1159ab5de1851afba6731e4d8f371283d4c8e0a0b8c25dd66911f3859771fc95b4ca4cad4a4f6abc58a36027504c55df7c2a09aa1f7014a2b5b2489ec37f86477c170ab8a0d5dc0e9a0adedb7f0bd0cfe85f083f90bea15548bec6364da1418f1e3b860cfdd2f20e8e71fa67f46eb54d57b5e4c99192296a39684e2896890ac2141cac22775591301e1eb7ef9a039a78b6ed52bd7ae9f81f68878d4ab59e46d30bd6eebe467066314cb6100bb47050b74f1e0e3125dc49b70b2f76a1e60ecd4747265d096bd5d08ac411adf987b3da805eca8c943452522aa61c093124c00b0cfe7b5e9699b81c35745c4f615f2208341dd1be6bbb7b33824c043baa02c32fe5e5b70a7ec13bd24fd1f7011f7fb6f620c35b9e092d62a2a43ea1a69e56260d444d7f91e19ebe09ffc54aac3d83604b1e6e0dad9f3b13fc25535496fc83ccf0dbaf83077a0c4ee5f6c2e8cb41c0f41fdb026cdb17c52a4636f902337513637990b41ed41dfc5619ed69d229c38a2d13c1a5d5c74249f2e4736ec3a6b54b5d7906e07304f5cb9d0d0067cb89ec7c82928a4584905d18672de92c1702eee7812b0db2d7a3e6dc87f60a5bb3e524444fddfc41d9b02bbf9aa26b79ff3ca0f84024a6c14b7fe242ba98e5a499ceb59864a2cf9d4bfb532e78ad7b1019495ce0d39cbe024dae38fa5ab1ed2ed66a0c5b02614ff8a37c97b9b827b35203c9d4a2de0434d244bbcc1f66259a72d0585fc9732d1b73352c82428e10d37d4df5b1d80f717c4f771036b8d93a019f136ad0bb6c3cd9e45910b2f0ad697ddb0f236d1a189e3f436edd26f8e3708717568c776403e12cc92118ca04c982e2af88eae90448032ed65e87fbf5c4474df9866c41172de4d14fda6ede99c4efe3f3e460afee21af3e25326aaa0bf93536e88767c1777e68092c49c8cf96b4509de450c69513d0c726fc5e1d1a878b99770490c376efd14920df43c0828dba958e15e969f9b1792ee64d10c334b759b86ea6ea13194ab7ef445ef1e74a3dd0a7b05f10a44c8ff2663025fe077095e7c572d84e87dfe3cfbe275bac7883f984291551e2d352d79a809f966ac813afc0f6c3410fcf95fa9b215e4422ee996e466b4810b04eb792117e80e372e8de733cd3b798ab01f13587bd900a23a471245bb6bba345d404b1a24bde711220d2a228c78de63dba7915d1693b255063190199dfa04c7c6547f2020ef8499b97cd92565b437edc23b9d53ec9555d2e1e003767aeeb94973183fd58a3ec2fd6ba13904a85359e741b83216fe379e23a29792c183ee64afa21571f8658b6555cb5e64626d621b85a391a808098ec80f272e608005;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h417034000fdeacb1113985424ba93eb7255615be0107aa069d0755b4317b2e303de57f2a0a1c86edf5cd068d5a22524028e400117fdc63c56a71f11c0cbc778f977d20e2697962edd8a38a2e748f603b11ac75bc92f09714e70826b67bea60067f3f180c03f32eb450dde6377c8f778c6c18cdc63a8b21c5490b96f1e10ee26d2650fce4ff24acb7a2f1a485e4fb5a3841443108b909366e086664da14d26b514045cfd15b81ee909eb2622826606527e062965b6f529d2b45a9e7b79b0199ed8f7956356738eb1a0b21e08bd9aa31a9fffb36c50194994f6d536430e170330150ba70b564686d3e3ede47be4e8fe1f957be097ffcb95da96c27631d1756f27da388c48927ebbd061aa71e0f3597765ed59ef5e0aef410553710d91faeab35292328d7c6d499e46e93ff8359f484941a0aa657328c9c56d6a1a8be10dc50bafccaa48aca468da34ede384d791bef009782683a5b04e005afb8396589b3eff239a463741315d0dc5a5732cf3095de40ad3a41e35379834601ca064c00e6cb057714d74635f0996c5ff505f549f255bd1b8b17388992d1730a6faeaf199f761c335e768271264de7a93f91f1f9fd08be9b17cc48a1535fa9a77f4091a3479d069082e98e284a26b374f419e8e21cc336c3a18fcc3bc16af3ef3b01eb54f8bd045d8563f6ccaa1102ed55329121950597a56eb6fdbffb2c09ebf10aa8c60abdc586a3d59f306da08ecbfdc0b713d86288fefd7c0e45d34d10392bc9af26e18d8aaea397942b83f0a0c7256e65ee0b7a7c0359985c5d401e5f0234ca8dd80fd5e3be9e93649175eb9f04a295fa32a1e35007506062800212c68da7c122056ceead5dc8eaf8c188d9141703bf612796ca24c5ad0b06c1d29766de19dfb072769b66186ca883de6027c22ca5539f4c09ac95e2fd8c694085ed54f7b9454fcdb8ccccb4a84b1893bbeb3c5ec913b5004535c4ad588809eb50055302b655e8635bdec8eafc86274014a36bc119ac752a19780fe0a3ba2d598ddec5224f9d3a551484239bbc727ef1e28b0d25373334ee71fdf1380fed6f221c82d5d40cb3faf41b819a0a7551b4d350d8464bf8851fbf05b20286e4b483c26eaad285a62cababf967c9ef88c755ad6f3b63eb48a61a6e9bb395d3018fc04c83ff8ee2c95a666f5545e3cd3e8116934fac67a2f7670ce3bf83f2fa8f63c3947cd39379849a3732299ca5b09dac1e9ac8a61c2a4c8aae0e64e1fe30632943d96f14786189632b91b27941f9be2167d82edffba09e37370205c32c7ad13cb0eaebc01eaadf6c48424cd1b562e2649e97ecb58df58d3affbd10a829d1f27207ca1864fbfe500acfcc112b7efb270905e4a56a6421700c7e8a3ccf7c778f55689c964d277d45ce99a1684b947e6374c9900e33cc3ad2e9eae70dc13581eb068ebb4d667f409a7b6aa5055acd59f106e506e6a6da09deed6451601353b04c4e208cc5c342a33c64fbf1285d70ae41fea82e27497049153009c6393ca8e17c548cfe2e29c1b345fd4f73917b40709dc5efc997c6bc5814af6b78f8bd7696952c71e0449cf1448bd0429fab4ffb612102349150da53baa8a1a5858a572f48fd3418600a7c52b930e4aa58bd266d43a520e618c6865a12305d4c7b376f61e577a58fb8e23bf284409102c1a96cab9f938b3168bbc94d64b22690ac2e2ef1727cb22026f3dfceab632425480c8df28230dce064c0ee9f2be0ee8d9a7ab55f44448a7656f86d4f136851fc867f479915ccf96503878a6a829dd741d2a7cce2338159a39c44a2fa62e2ac4d1ab06599879599eded265aa3c6b2de2e931c2ea7934fd056acfbba093ec6e434dd51d1b125bc2ca42e1d6fa2b77ffb7f2125460174924963c9f2eb1c29c3110f0817c7f08b07c2801558670ed8654f24487930034916328eb0d18391dab3bc73ad6cdc6fec76985f0c4732e2cfa864cc0549a0a06ac0c836e17bf5c788bbc4f3f4959e83c3f3c51d759ccd57b4da708c3503a939a9a172de0803da7726b088205b2a8844bbab499485ac6afe46d462fe2b39631bf956c980c6daf1a37107bdaae0e7c0d3f410830854b58983c413b85f183a6413d9efc3b05615bf8a69f8fe91176472c81558b32a6e36803cc1264fbb885d0f8d74a2f801c519129c143c3ec106ade2960e3a2517a993062de77ed26133a7a0acf53a813339e816e61999ed9bcd5b3e237ede5cc4411cf08046fb5c5dfa7f658e5851b21d12c8de22998f84ff8cd3547dac6e1f27655861c704fa7fa3e7d47f4799b8ebe047dc5289020671976a62b51d25e7f681b7133b35be88d995648e5bf5959e70c291fc974d1ba2c160983f94f0fe36cfad808b73109f6a296cda22eefb800b0001f61a75b795a4aa8e59f3ce03fd5e82dd2e6a5bd7aa2b5863635758795856a77270ae7183d0730d281bfd77a4e3497acf7c634699739e4fcf13551618a8c2b53664efaf68049d46ffbef7da774f43a151504d579dd0b4b9651d4bb6c0084e82fb59939a20b6a8cbc858b71a27dfc07302dc4144c750d5ff23c38ddbc5031d351514e1c88a113178d1d001757a02ac7503e4914be12c2cd4166a02bb29f4ba903bb2c1d33c4293c3440ece5841b43c84c83c38f199187eb35ae4692878fdb163d242fb13aba3b03e219545e0a7576079e2bae2b80c5ef504b38ed2117410c3f3dcf7125ff7fff70bce020a7a4cf370eb0a611ddf13c73203d7a074dff9dde15a666c2136add529db56c3b8a164e20289d2fb6f46126c662f25b74cb49a4cab570404c463a6b1ee6439eaa527be4d8c1e73cc2045371f0adf82e6656ddc5695bfd40d4f11a338043292b59e84ac553e8eedd0822f7565aa6bd52f8264b3c80380138f8475288c537a1da6361bfc73;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8549c48668c62268b5f557edba654e425d72def12ba8169b4807c1d9969bf7cb52496b31bb0961a4697e8b1822c87cb059f9f4fd2261f0335a754047e0cff46b20cb5d2e229d6e2324abe7b26229ace8187aa10690bf4a106f7a947f84d7519646193d028955718716d5cc1edf931ab8e4646b88f6ed310cdb8ca67c36b74f8e8cd2e08648e9f99250c64568f34a9049519e3f1f88a9c95791e47f9d548d722c8791e633f4d0f5bf27584f3e210ad8d71373676da4403c7c1b0345fe3c10cac32a6216183f572e1e0bd4ba626fdf5ddfd086ee4e2dab076b65b29f48e9db522fdea749ea6bfabc441318be8a20bd0057a1683469fad5af765f6b3cdfa77e85cd94fa68c5cd414c1ef474b3c0a3dc2dee3a9b4cee2cfc7a2cc6ef0de5cbbf3208cf75730e4e4748e512661f0778c0d3c8c523fc3cafdb69ce40ebd443eb6436e4274e9b76959a63cfd592cbc6ff9b604032de4f34d95d925b612dbf1d002c9f5bfb2ff322e4ee52491290c2ca47a9966490bf47942b6f9cd1e9b130e2a0d4087ace5305b5d5fb8cfa877b251df076afd4394f0740d86a796d73a46d25824cb56a49b25c9bd6ad9ccdf72467273ab0f1f39400032345fca90d4063ffdeff4612112a0d4ccd85f1e27c1ba1a6ae7029cd7fdf0eab91d29d70a5487af6f0dc91706cf1f64f007317d9159f9e42e5025c99d263118053820e2aaeae8afc6a3b0f3af038fc7e6bca6570b73c1277c6b18387d5494894247f77e7dd9b32fd8d1c51eb6307c52291d070ffbe5679d193fbf60f49ce41faa745f965511ba18d06366b6fb37ad7e3ee54c4bce19b202f9c3254be9a145eeec9c3c681cd77b96497723cc10921bd5be40711880ee67d848b6a0822a7935504b4e1336223eb92f59480d2cb81da55112a0c8e2d672e9aae9b89381307f2d661514bfb942a46b38a1a2841424a0496b29e7381a4500023f5f6cb237ba2b6fe1715c9a66c9f4d4728874c458bff7af16a109bb2fdb9c34aa8623540695740977a7d8c41287c5ef43e363c8b9d64f6b50afb7aba26998221eae3dd40c72f445aa9b5f82591e61d89c52410894daefda7f52b93a029d15288f67f20feb5d666dae9a5f84ab525321be696a2cf428e98ab2c166c13481b2b768f3e6e19d4169e4f992c4ab9c11441b8aa818558c604806b0567d62e62259ac0a4e3cf33881e571c37fdfc6a6976aa6fa9ffd7e7a4f032d438c593d5074542129eb9b5d57e5b6dbd13b4e1671e73b8f94ce90b890a785c5e34021f7d54fddf23b70959085d261cc21c5b07405dc06ff37699f3e0b3ee3db2026d4c7426e93e2c24351b533bf4398615f79b4a395fb5d2f50242465c2d0765cc49b2da0de5f659a25e7648f685e97c024668dfab44e4b18f5fc77f3f7fc7c2ec75d11732a0a909f014f3e0b796299a919250cd327f0f1742446c647292e1ef1ee2a50eb001e43b3def1f6fbc9ccb631995159d4dad6cc5be5c4589d6916000a7cb24f04d947ebbeeacb9563138ebd96587ddfb082bbb7e4d1ace9345b815f86d6988fb6248f100b933fb3cd80dacfddaaba49fe0ca4f6791a3611cc86ddd7530d836ab5d169304975e7c20b485165a06e63102fa45fbf996d46d4095c18fd0f58e3192ad8cc4a38b32769dcf271d9ee72e02adba0615a87a0ef9d2e09578a0d32da5df5a3248f554b052cdac3966eea85bcb718dbd75640ba20de7cf550fd113e6522b72df113f8941c1992a2f8000905c02796b3f1efa4c664a767118dae33e883ca33980839ab2e16d199fbf6398e5cfea562235afbf3933bc3f795737dcfaeb430006d0420b17caeb720aa1e35c5f1d3f6deb413d3743a982a728ee8dc213430b3b476d9e0990548d7263a108b37c287743d2cf1231cc12e279dc62242bd7b5c2b116231d7aa7058216b26f8319f9fc6538dc69a8a3269646fc046ae8b6a82a71edb38740a28484a57e21aeb985f8538852c0d85a8db5c392c51bd6c2a3a5f16274877e436603d93c32633fb5d10b0b54423708336728587f7ea8adfe1efa6c8b0df92f5b0642415363921838f61ba94de2ce9399289da5978de3f33ba228b6acc6e662a1c98d5e0fbba1212e1530dbdd48236590185a90c1400afbd2604d7ec5e4c1465abef349ab873b1e4e012b56aaab2a9fc7daf1de49bf14cb5f63e22903670bd541e03291fdb0b6d5777d5d45cbe98ad2e7590c0bac47f51cce04c800ca558bb6e1f0ed9e86369ac313e23811bb93047b54e71e952a3a6bfba72aa492e75bad9ff0bd501bf1b323b051f9eeaed47b4b4fc062f84f6a3f1ca89c2197fb568d1409e5fb9bf44adcb5d3c1153990c08bc545f8c91a0655fada8f143b1e94f78d75e9514464ba488853a9fef68214701769783c2fa16ac3ba07246b20694ba2cbac18087645ed32c7d1441e29a6f7480f11beaed94cdff5c2ec1519c215632a44011bad6c3c65dc0164e5e641d17128c1b9afcdb0c996616de73ad476c2745c0c3782a611022c5030ae870d09861afc3f9de05ffbef26392276755bc0c8c19899939cc487787bcfedfe084cf5336b88dc6e0dfb91e9a0af241fa65cc324e23ad2be061c62e31ae6a19ec152f9daae3e97f887bcb5de05dd168f94b5f26b70a74d3345af0c23cc06331697df13b98ce28a56a85bc8912f484e7f1ecc596e04ca223f98343e4c471190e39d945520bcd145d1a5f0f75db418da41d2d243050562c91bc050823344894ab08cdbdddbb79f6a6d4818f043a8ebd041c232ad1ac10668dded1322907121d5a82ab1616034efbf9105bc9185f0e2029a3cf78be26ca2cbf643b123d635184529426ded5836f28fa809eee34520c86ffd0caaed11d1949ea8983e3f61e2434b7145e2903e80cf678c2d35a36c9107fd5a59;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h81f7014a7af24c5cf30f0e7acb2b9c8f37158d7152079796e2c7e03f5d1c41af5fc0bab1badc9a11b50059b54275bce1120b4f69c60b15009162c55557cd65954e9a2c3191cc829eacd5b35959d54b86aaab046512405a2aba6f0dfb96791074f22d4782d76b97555eae7c57a16d75ddaa49c44f8b6469bba176b961419a1ad1c6db0fa225ea90ce67fad15c51d8026b471406eac4ed9b81069e5eeca353cf15d925c07a910004b6a00b021b53b858fb81946ee40fdbe95ce0fb2d040920450aed77841d47f39fc4338e92027cc0a80804d3865217c8b76470e11cc6d681f9d7a897dcdfaa0ba955e4caf738aac439094c343ca4e77e53ac09781aaaf6ea2109397ed568c13fad7ab6a4967c275a72beb68989f4eed63d93a5db568bbd8ed5efc5d0a0c6f1fc43c35408c88af07b5c3ad1dcd93c1198e5529eadfce0155f107c1209ebd20750be4f9f5d1799bd267f859515000e3f852f8e8ca8ec938ec9f530d874f43ec664b3e9e506958fa3378ace1aafeee534a8144fe7e2560ed72c23eece66f91615cf3fa161146006d4c289c96476ed391581ab1cecc3a48112d3838ec76f794cef722df2042c9f7121147fb1703f9f2dcc14a3e9bcee3da9903326ae54b20bdb930a274fe3c19e5a837e3a269bdb7af1ffe996ef05cd5f89294bd1000785fe406da295ae72caa8ddbdb7e6644f9ba7e62635e154cb72c2ef366af61bd6a448835829d18418c66b53fb70180bf2eeefae80c43d4ad8cc944185c2a274d960d111f9fef0bb56c219b386f136f6b951cae5ac55ec4d260d3c2dc93d2e60ced17f48e4a5a0c88990839eb4018f216e9f3e652d16f3cb76a3db92c20d54685bf0adb2bf3cdc641e9e186b59a0952bb05bc066118b437404003d6f05b4b99a040808a647461e6dff8358bb6572efbfedce4eb922258acaa98c1ff4b777a634c3235e186c091a276d8d012abd2333034f8dbb5f9848ab277415559b3bbdb950fa217478c8d893f3852f457141f33dd23c7ed0bedf37aa252992a2363430c93a1ae03387869fdbea537a121915b47af643c928875501769793c1ef3c90bc17f9c89de70d33b088222c47b46c3f8450676e30ef4b9ac76e0c1acffddae58adaf20cc2209be8c79330d555f32d4a82e1386bf4808e0a363b960bfb68bc06bbaab73bb8250466cdcbd9c6a138fca2025149df2a09482441c125c292bd0ca3d2056315bc8adb267b467cc9807b87f07fca2ed414d2cb0ffac542c9a48645f0b480198aff52d82b8cc7082f7360f8ea9248b95b7cf79638508e0a137cde537ea45ebe2ca9c88ebd3978202702fda9aa3ccc392d844c63eb760ad62eede466e61c006d4181dc490b32ff03975179e44ec8e288ff00fabdc92952458029002733402efecd91200d3e39a71ce770f036c41657ec26b3b59150db6333408095be42543d0e5d2a29f25da6da4728279369f150be37775f1d3745e886fce33bdb729b1cb50b83b6f290c7e1bb95c28a17b452ff2270485d3da2d4adf637ec6ac36a0885d72a75c4c2893a41b3da657acaeb9b9f77567a05a823485687a2029364f7c2b45d5c88d32d0fcbbeb0aabfe115e5381158a5f0750f67584dcd040812e1e4517769c206a242a7a36ad0b21cde097f85bdc77ad4d988bd12fd2c3cd324574b68250b4eb8373be8ac9120bc45ad375143c0d547a7588ec98e1f302404f150c34eae2315f8559ade3742820aa0916671c6bc2e5ca93f501283e3305e90e01e28f9447f34487034c7b121bf383f8424712650eff6a61be6e1554be4cb1a6cbd9e5e4330a626aa9307a1029529adab6d5bc6666ae84d80dbd296bcb21227a3220fb76aac1747ce16e64901906c19e8663fd5663035b6319366f4dd703c81caaa5e1581ec1cc83097be69c94d0404d74d4b6624769c02b0a3ecb473ff7c910f0ae2a8c2a61794e125d60de1fdbe2ff5faa7a960cf42e735b5000989d0cdb8b880dd2bfac6a1d21e0acea34eb0ab1f64b2dec3ba3c7f923a3d1797e51f1a96c9670c5b4faf6b6c18c37f09fb4d090059276b93d3f10de46c8dc646b0322d35d3800c8c3dea5cabc6f19e4b5f17830dc54831ace28744afe5c61d4f5cf068b0f347754022affa28c58b955d1ee0d283a1d0e65fa3075033ac4079664bdc32dcf8be29b3f6788c4a2cf622a27d124162499fc61499b9693d9abed482a78370d14daa42c3a5ae13a2643c7240f7b860363cee9902eb669e0af7630d9c812aa2994c6a0f7e42ab23e0c474cbbf2befa5030a38761fbf918a3976ec90772cdb051035d41e2856d970dbeeb71a0f6a3ea5d4faf057ddb0b1a8e3ecb5865a01178522dabfcf89156d7f0baa48b18326cbf53ea94ec582dc3769f2f05764057ce7e2b88b22877bdbb87ff219c95f9be290bf198c18638186876fcad23e7eeda27508b7fcb87a105723eca7b6ceca00157c93c9b5686d084540dc664e74d58dedc1e8c78e472211a7e94fc26dddd0c55cff9ae428c250c58421a7abf3d0fd11bd7951151a1966d7daa91aea611453acf9f459536dffe985a890c2c9b530f807265d3b12a3e4328035a5a99b1c02651c19a8de86cebebea807427acffdee72ee3f726c0b429bd122dbf9ab736734eae55b3112f3bc456389ef67e24c94ddd0e1230fdd13b0e2e753a44d5d8afe5869cb94bc373872ec77a31d7ce74ef5695f30a7fff6aa9bd8b976077eb5b1faa81bfd4ed50758770db31962e99e07542bf3363b924133424993a00d663cd1fc635e2be9f420e1ed8c6cc0d5f883ef23a430644eae3ffa685d8afa54cf1a3b8318c39a15771e61dab56eed0e59e675b8df3f02c0a0f46fa78edea34a420dbc1f6765ad41cbce3d62b6bde2cd2d6fe4a1a062cc6ee1cf1fd6304c7ccd3e38;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb3b80fe65e57c2914cca95e3696e22fddd7cc27d8518c96aefba0fc47bddc04860e56398fc7094f2a10fdbe9cd6f7598c861eef8b024a8d4cbd87d129d992b3bcee349459fdd9a1d1ace30eef410a3ee3f065d7673a3bfa3714e41bd1a284dccc157e6167f52cad04a1f7b766ca383b74b5924bf2c72d03c06bd23885d6466de5f244b9238860090a3fe4e1c324635a15174035ae8abda84ae46ae81d637224d17eb285f980e36f900cfe8db356db700c0b55f222f49d0c069f5f27044bf26596f1e7871416cd9c2cf6f55f92d841f8eb3846be96f5d6e1cd108b2bce07a3d43d01d25a47f90e219f43734d92f1d9649a0eb758c4ffa809adf63a2ad37eb3a47db902f267f3da69d62d25c45c887a1b4e10d255c69980db3772a72b879c0717936ec9e1877034d1354868e75d3ee7d7818a49b93ac8504542bbbebd6c42ec7adcc2ac4e7e7daef172e6e7fb87318911920a02bd610810c4247ca8db8902553e9a7e6e83141297f261fae5cf5a38e399f41968f29299a3ccdf20a1a977bde6c32f971f6bef94299918f31e73bf56a6180df64f6f376370c142fad39382355ad9ec4b1bf06ccdf8c9b1f8df4f7bf95cd5ab5d08362d1dd4455f1b7050c3062b05d291d500392ddb9ffeb8152fcb4731f831bc23db45a749c0a75a8194828694f73d471e2be348022de8cd983c9945dd2bcf43216b5f137b1b3de8bcb9c1554fd2b9e358d583dcd61e6fa32fd121c4e3fdd74049298f8a73b259d0c022db1d36218f135e7728d3a3a429591f88ba961af10cfd590b7dd5bc09606218275e60bfe1e99572d42874e597b20aed453c436304564493ff9169c08fa88e18cd94c8b2285eb8dc592c312b9b744f86519f3dc45db01d2e39a340add1c51c4c9d70d095a5ddaa49f5950a4fccf99755d628895d2089087733746de129f6dccdf33409e6b49607ab6760a8b6b5d6d60ea8585e8a77ed62494c30910198e538237a9d8b84db691e92dd69964ddb7181686e5d06f51631ffdfe5c7ff4a8be0787cb4a7cdfc31a1954b9a59ef1884c2a49c2187b3fced5523c687d04b805e17d89befe09a53a126e58db5d0097f1e98accb82a29b07e84aa22a45e589ff3c38dd9b2810bf95e812fa30f4f7137632ebcd4e76a75ff9d5ae6aceb57cb62fcd40b322e0fb75c58ba89a768a8a6362514099afc1e21b28349e7de3221b7073b649b0b2fa337c638c9381cd23ada16c981b02ed7a9646a4fb72f5eec391511ce4aad0b8ae3b0c301731909ffbf38c17958097bf2737a6ef4c71c98702c15d4ab30c1af2f5ed56b657d77ad8d48c1a88ad7ef346676a47d359d78420045ab00d52219a5501f8b884fa8d0d2d22aadbe7c7a373fc1bc43aa6104da2a4668a9e9393b99fb5f7ae05cd9275d828af581a3e0d826cdde9477afce4c8d4ca0ed60163e15b127162f5350dfb71a0547388266cffa31b1c995a99519baca14e289ee9661ee5049d3f781d5444114dc1b2703938d0ee385b90e19caca812762d9c5770212ca9124911286873e27974647e5a435d50387cf0c33db3ab92e056157581ec140f696252177efe3d037df13b0cf7f779021132ceca7c9accbe93e28ce33583d4113591b9ea935ecb0286709dffe34b3b929d61d6d04424ec435129dd024931bdddd4847cca55b886ada62081366aaae57aa71c0a1ba1e9586dbe800158c0d1fa5f3e87d70ed3e6fce8995f72f566b16041976d49381fe71a7c2cf954859889d702830f95ad63b7367f0987a3a9216e76e060262d62e0f90a77667f7ca4cdfe5c9a77d8f3bc541148be6b089e0d15df9f4164a6efb1b836550dcb2bd06e157bd9f7ff7f7fe9d9d88b3adac0030c2ed79b7a3d5c98c7121185e757919af1add3f01b8ceee3e46f6d98144751b9738a56d77b4e064c731f19eadaec7f6df070aa0705368e3d2e8e817143150f48fdccd81f9344450b3dce9dc1a696022764f39db0b8f4954a21b4916cee6a71e56a7edcbbc94c243286598d59b4513f4c43eca2524c53eff969158744d7378cbcb199810b3ff265185965a88706c00d0b6c306b0f67ee4fe0bc67223acd59301c5df88d5b3695e34c276f40cfe9adf6d36db12e22fedefd5cafe6c18afdb62d482a57efb882241f0841f7a93e318599a30f7f8d45bf7f8d6d79836354f5dad07d3e8c72f3b157d75f444e2ecfa212df7e40184a7b12c30e024319c4f95b9ab962b7201db38f6423933f995e72f56e7ea904759179dffaad03eec98abdd3f4c92863965126db1fd0e827173bde73d8d175ff2f2acf9409d6091aa87b36a864b8caa34d269aa9246caf4ffbea115cfa83fdc7b1aa5d090d18ccef7ea3a54bc86d24121eddfee1ea35e5f036c952e3731c4784776d0bce5cf023f3b442b1d84435755c74bec412324ff31c20bc5cdc978b544eb5d4ddb56725db4def48873a654ef5efe7aabea9394b670180a5d1fc35b9c72d84f5c0b92d2f354a47e2dd5072bc8ade63eb8008771f8c19190c3a1cc054d73cc4108873cf3af1de8d65215ecf3264dc88b6c771c04d30183c6f7b6edcdd489aa0cd6b9c45738c1987e38f82580f99fad53e35bb7a5efc0608839b7d59e694979698c94d662008f1aac4cf91e52e9ca57164f0bd1dafe805209a3526ecda18f1b7736e5903b31f0b86bc72a3944a3dfa2f323ad586bcc3a6ebe3a68729bb12e0e31d6e299440a7a938c12f5c72b1d70f957c84b4b45c86d4ca6504fd97c3094b5fc25435dafb98ed3982da0128bca3c921561342ecfe4e850b41cf04fa5edd0d750656361b6dd15631d0ab259ccecef912221588d6634dbd9e9274d4d46ee273a8750c0d58a5c88ec2584333fed3ae170e45e163700337c57f7d0f3240a832877c9c3e161d747933eb5cff86e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2be33a1fb84849ec6952b8f08227b53bff9d8bdff0f0598571f8a296c608647764d839f6cb16dc72954a3a2c8ded021c4ee06caa76847012181abbb1909ac81ec181ac8709fb8926095e204b28a3535d6becaacbd5aaa9f31469f94e3ccc9a1fbc20a4cadbf04961e5774abc97f70f4ffc375f2879c32eb98d568a7cd18f6af8b8b03d922f7e51d6f0a139fe80aee7e2b1e9cdbdfec3c043fecb7be133069ee518e60d7bb0f3cd5b84102d01d918792d966e51f149d69da8dc4ffe7e02d0773b7685a258fdd475006423f506cb2083b26b93e39495c10020b3c46b624d27bb18b9ed43c9e86724fe87d67a86553bef4cda635cd6092b4148e90ee09b031b9b79f3575a527ced15971c4b3302721a268eff9f73bc43617f332ac6aad0cc5d40cc80dfd8fa37c0dec57040d9b6cfe32ef1c3a1970c2e8f1b30e9d28e57c00bdb438a818a0cba7cdf8085d4cadeffad9df396f940cd65c7cd591354c0fb46d95b9369af713cba9057615bdc830f483dc7437c6ad2e6d6c026ac6494e7c1a279dc68d08378dd68af461ee4d6542eb7ff6b696908c64a9ee9ac2b1e6bf50df4bc72683579f8d969317b9e23a8f4532aba3203c189709d3fd04802678c07123cd91a68b75d8aeac8c2f00f4600e9bad3f424fd76e676e0b09e0daa8e2aa7178cff444c741e967a0d11b7c3823253f066a04601a85836b01136a92471bf0d3976ec5057643a98b9f02fbe8380f59948a1ed0799f1ba2cf24c9d3b60d20907117aad78542f71e0168744ff5b6f56ab199d031dd42946c1ee34ecc752490038f4fa2ea82144402e5ab338c13835fa1806172626858dd7f38c20e02ae1b8191e95b93ca779d6991b9fb53109a1452f7355fbb7fe31b9bfc0b50457bf3fc5d56068d8d36219e8e87b088fe6d50611797a51e46fa041826c5877c7ac204ac7dccb3e9fda00cf3c7c82634ea7ad580fff786ad53013f06364c85d186067745bf972b309fa502346128c42fe1c93d0b5908f615277e7b577f4bfd2244c7c77371dded9098b62a2a9eba39b06c1883842c6cd38e9c87fc508312568046d93cd01504ba360ab52d38c2ca65326b7ad066f77e0cffc80659430c99760ce4fe62d7ce15a6aec4c5213effe7b418716fc9963fb8160ccf7a7d3b30cf245f0ab91feec6cd6ae8f9263b1769f995916377f433e243fe034839b5b26967cfb1aa9e097465249cb996d0d721f48ff099bb5b63634218bf1474eefb8f857471438c0f9a61ec24a8afbc6e12bd39ba59b2e784c5c4d1edd26cd17ea3ae56ecd9e1cb8ef3021d3feafd6a65c712d11d2e3ff35b4cf8fd7121b00d35bcca19c35c253060be409de893b3bcaf9e8894caf09beed38f2acffdcd2b727eb5889993053bc3e3d75c38fad9c16e9d16d753f36e24afa8b3abe428986f558a8283462f2d2e1f30987ef19c4b82557349850a10a191bcf077e188e9bcfb8516f51c23875b148461f43f46ce9eec53fbab58d649c5c35deed9f3989069b9327a7c94198bfc13089be3bacb47d88d5902d2e95609b0a5de3da2d135d35ceb19648bb3ac0b829ffde37e9d6ca9b82266c058520f5ce3aac498aa586ee3b376ce20edfb17ccf195fe6cdf26dde0f05b9ecf17166f4669f25216e943b6f7d87a549fd687ed2fa76cc7de7e457904279ae38854bf79427d9561ade7e76762501e6ba2d88e933f7e90b46433db1d24ee1ca31e237cd597a99aeed65503ee97b31378211d07989e18a4cf46f1d4583da32d74b93bc62e672b3c19c41ae834229216859abbd8f138a25776e99023955433a23b3dbd021cfb4182fca499446af21cf384cb19750e1355e2861d8e5b18bf804a1f26d775f4eeb27e661b64e1dba5e95cf6db4715096b19582e2e19bc872e8d39ff8e38d9e9b72d33d94d634c173d9deb2b837c57f74e192dbbd22688a2d90acbddafab8817dc364ec9f4409d285877c21bf16279177c65033c80b70cbea3d5f0cf13d46c588a3baaef99c72277d6a4281031839fb696c2b6f89b2c8b9a980d4ad985d68d896d727ba53b179b117e727e4fef44a29d3eff9c937e157781b545943331c88cdd417fa6b3af05659c83064a0936f286b8c26ef0539a801bb573297d46705141d620bc9bcaeac9edac90b090762bd8fba210f9ed382705af4d31ec988f5bf42055d239eae43913fc242ea050af5f1b085bda78ace2992002bd5a8503efc100263a78f8243d56b4ea7114cca90c00bb825e3124e6f30814680b8f57616fcebb5e1ca2f438e989edee70b6546585fb06ecf5c08bc91d77e149c1f0276a2fd5bf5697f04d0bb50d9e9cdd38a843c672b9a918831def6536132151bf8b1e47c1d5639ef64631c0ec1221ecf90c4c35f422ee227ad5da119a5324d778108c1a37021b0ec076079b43f45a4c39073a297fd4d6c71739129a247b39be85abd6b3771659bf7ff3613f399369c689b730e617d550d5d2fb33a7b987170118cb359c2bc83f5f200c4ba1a7013799f374c7e454006719c22739789cc900040c0d772350e43905dff09a863cc3bbb5dbe3c5b12caf3f76b6e75dce2637a0b59330b0fff5f48a5e5eba1cafec727cd6f9bb8e3ef7662b629e95849f7629afbc02fd7b9993dc9d734f95d25e4b2212ba52ea88f7864df3c8aa63ca4ee437ea553e9efdaedc1a974da20812753f2f2893407e59c2c3c077aabd3075a1c91b55c953c1a3c3da1aa200b72f55d2403bf4ee33f9e34a33e1c6a5a879b821ae597b35a20517b925f880155ea5adc9da5996a4a7d96e97eba6c9cd9561ba662fe2101a778dacbf11848bebd64e71368303b0635309fd060bb52a2b1c457b3bb063084bdf37b72bf61f19ab108cb31b41c6e0ede38c352a9c941fb2b958b06caaf63ce6abab4b96ab12e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf7d0496251bd83bf18703152cff47069ce4ac330b47000ab34f94aac14c7c348e031fdc53fd9374aeb14263b80a04c78e77f1991c9be9542f76fc8769028ba6b7baf8c97b819cf6dd9aa4806cd63054a04d328d950868eccf47f770e624e288a66f3abe17fd5ab1b3a15db081a0db636310f507afee019521c2dccbb92121258d8c61cba5b5d8951d49b9f0ed354977683b2721b56c8b7ceaa6919961d41964d0e3800a4dd2a912e09b8b3bf0830f9bf97039df12455cf2d18dac8ddd2590ad7245e2b7d53b15eab17cbcf1d237365fa69e82694daecb53dacd2a582408004b85942604c34406879621667622fc14681b393b6f2179ca5000209a219435bcbc610140edf11d095a249bc9bc0b90611cd46beb188fb3b16efacbfe61a76f2df2b615633ff5b76a81b0f21c812ec8e25a4130e3e3153066179d7342afae53588a2360235bdce80ceb383e8eed683cc2ff0de29bd7f3d17ab5d65527318c4f576d30331a93b9d2df84af20c8458b5f3b30adb0dae9e72e1d7c48b41ded65ae9ed40967a46e575a1bd91613a13dcd6d8ec4e57fd2239c7100e3c6e7be33c8ecfb85092db886ff1894d2330a8909e49cb9b13f88f80dbcfebbd6b8949a5394efa1dab712fdb7e3c50e5140613abdc355929557df4983e72ce88e44cea407a1453651625638f599692de991d521e06ba3d6bd6d9e3f51b180147c5a621e001fc7ffda583a21959d58ec4169c4ab6fc9160ffa41c8bb21607570f2fe4e127e6eafd00c70405b60c9e8cb2e72aefca8a6e7328ed7c5554462fe54b9e2c4b18daa27c4b61a08fd01cdc2ca332ff51e8740837058c30ba2f0176d1f0eb46589de168d2cb9c1d7eaa7a84d4de982eb432b54c7f6430398ab82bd180d550c1a754f01ea43695beb94ec1bf774eea4f1e1a14449a93859eff7c2591cc6b98745750ce1e08c711770a2603ba89dd30b31cc4d72cee1b6849cca026e05a7bacfd6bac94b38087d01840457f9ed8a7e6b331d43702451d399696b4cc656632437491ea23c70bd11463a9494b3a366a15f028d01a02b52033b0fc57b06f895272f0df5889495834538348b26a17728e4bd7d5a6478b733d11eb534747da8426bc338794ade319953191729d06c538acd142f8a2b7b2b12696de9c70aedf12d620ad7c0f954f7235b9ec5be38c84de1d69ea8be12ccfe728ea8cdd3437ae7ef1e47b6faa13f711d58b7c9487b37b7f007f43d5b751513f57604bd636441f489b78fd8c78d927fe34820e2c13969fc99c8d70099974a70842bac75d4c9d662514c0b20d99f2ed2ae33627e260c99d23df6cf9c189bcb1a333913bf6c2b328eeb89980d666672151c167a09c6c7d72731ba80a8b1cf173fddea86eb58bafbcf9252b1cf53be0828e95d567b24c3fbbb5d305f94d0a3ead238eb8044a4094e299ee5d90b78c7ff2982977630a9754333bddd5328e6777b7aac71608ffc00304db72e808dbcf5808f897fa64861c16b211e8988628551bd64341859323ac083dd737d17d2c5518472b2c60586f9a0599200960cd1b6c2ba1d0efb18934ef3389ed6b69621f5a98ad144e8e156674b70cbb9a69c91c62851c2dc399f1dcbb56e2ec6e6fa8e4b8aa27ad848499b6774473ae867cdbfe218470dccc4c62dcff7aec21df94fae24d651323dc200a2c6c0f77defef5ab588b4d405931fc216ccde45e4df52a1ec5556ca9143c3b67d42ec04abb15ffa4e882a4dd8d7cc03b998612839d150e3d77d956c7efe3970307c31a41940c7f3a83b6927d44b5a093e00624da09d2981667fdc49f47094f8156fe77a7190d4d8aa0d36e21f678c8641c099beb013dd85db77b96991bf053e153be978e30f56da4851271c9d9ffaea1a35b067301315615c824d3504d66f8d000c7d1bb101b2a551397db34521e594a021e6bd81f5aa23904e7a3747afa550e99c9563171eefd573046862c701bf13d8458a06e260b6c2c96826f8ecd99d51e20d16db6f5c31b5c2f4cd7c5b93ab9a448edc6be5c4017e0c91a1d88c9391faeeb07c1041fd483331007527cfaca0fd097540b4959201eeb2d4f0400318241e3ffa4b73da8f6278a72d418bd3a90ab5beb427399e1c2f2e58e80c4a346b3151406b91a9bbf75b052e4f3b09c7a8ca2461d2e17fed1cdb81128e8be1c7600e01f9c52085e46a380bcae8d3b2ddcdb33f71c2629a1d381eb566437f5986d1bd4b371d7bcc7fbb63a8cfb6b21ed10f4d64490e3e3488f3c32e493599c348cf05209d442e6e63c4ba6ac2382522d2b8d5b30c3a5bd801143b2612a0c70306c8c8291cdc74f7b8699b39b53ce4f61fe69e9d60ef295697920a0ac5eb08582336689fd8ab20420d109096fbec15b16b11c2cf163abae644d3916b73bebcb941c950aaeeecfaf1aaac7789d9d8c7cdcd5d3d6408419c0298a3f6e6a4937ee45ebc97a9c9d47ad84f14db6d7d4d683e001ca8f4a01fc61ad6397212537ba1008c496090f9bd37b0c2840bc16c2a63708eede51f82757a59d27d4ebac470a9e195816d874541c70183ac261172797762ca98fea7c245eb4b5d7e038a8f2cf67aafd028a9228838a7b8de62cd65fade7adde57308b6e43b8c008c30468933818a449a704657621d13cf3fa1a5d16ceefcb02f880e89417ba08b6461f26cd132bc26a0351257154e301048738af2622724d21581ed6a54cce52fd97227610f390cd8a955b01eb24c17b28838ee9aa62355b86cc8e2b5470041fdb98d8b4c363ad011dca7b17ef1ca1cc979ed53c228d1aefded76534fa5849f38ee8c60cb4488c525433a5fa8537c068309508674941afabf955fcb07cec478c4f68db1133c242c5461b1dfc29b5254572e18c15b954146be3e7a6d388f532280a0b004d17447230312862;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hbbb89d050069505f12d239cf29c244a26c449c1640859190cee76e338200cf165e5f264e46142d69b8e87af8932e7ae70c365c79bdf643f2756dd07c3943d763059236d9158ae502370290a3ca2b522348c8a0746802c888b128c9a6c0fecc9aa5642d3b61300dc68c4af6a0f788900b5d97d1e8331aa399194538bf91483f81547638bf326c7aca0f4f751f6d15deb5edf38406486cb8fb37e8eacca14c61a8f65153753aa09993ee4da4dd93eeed5943fc0d38f2948c58a6c2970db07c78ecbf256454dafb1d135b5abc3250c0c2c41ebbb64d8415ae14b2c07fbb687f6f3377d76ba5457f973a585124a71e5e53a2464b904bd0a97698d24f1995a08a641db0957de874e8c31d1f10abcbbd0cfe6d4c7a174440ca39ccbf693772764e0507a527d647fdc72af30cde208d487d656da9f019e0327cee75c3692dc4bf800cbf1771ed307d9a276f1e94be2018e902175a54b660e2a42489eef2dd0f429216d90d19ece307c1257f6de01a71d27549a91a5dbbd37439204cd7c2ecde4e94d865e68bfab72f41ebdcbc645b0743152239b23c319968b3ee5a2d187d69f715ec4ec79c84a92a0ec4c577c13ccf36748038c08e84ae3157dfeaf87eb1af5fbae16ed7baa2c2a973d6c289c7e9c702616e2c2ffeb3020a86c7de9ccbe8758aaf5dd9573bfe76a53dff9beb00b6eb9dd64585925c27a4e8982962ae4da1331e8e3e5a0204ac1ae8a7ae5938445a4223cfbecc846a0aac517d776ba2f662d74235bc634e7207bf2f7c8e875d48fdf655c36eca17db0a5441d202aa64e6fd6c57b72371231573d64c203e03308f3d711643dc4b5dcb0e8ea7807b4b64888354deb4bbb28ca2fd9b7bd99c9b225eceffaafff9b1ec7833f49c690b1b6862bd51286aa1370a6cff417628574a0bb1a581204b8f736e9dbcbd3ba69731f9915d556240aab662838bdf0c3b127d65aefd2621d6b3825de470d05c07bdcbe3debc93d2ad5e77842fac43d453a138f7e611c1d8dd5dfe2d468c072faf045efa51d66a8bddd3d5926e299e9b9587cb29b9660f72075e1faf83e4e6b564b3cb111d81f301c39972f8407d5966729238f742f79890263d9634256bf14e665ddc717d98609699ef6e68a59629d7bce60bf3190b30c81e6b292402e02377af29b5fe3d46c029ff5b21618be5ba26c943256194036609b21761227622d464f3d7f90ee17ab172b20dafcb1856d93638d8353c5aa3407ff0e1da95b4acac731b5b2f96fd5f523bf4bbbacb01065751382614888d1a75066409078814854363777e357ed02466d77ca6bd8071136c496d7cb0a092b8592e2d96bb7a7247b8fae9893826c84740bb59298b627377b6b374788bdd721fcd08074471b97903e3f3e2244a6fdeabed6d34987c642a0e3557c86784f034ae1c65fc72bbc140a4e61eeebd8651efa2304b4c180676b7570af7b6072389fba05eebe3eebe11373e6306efa6a83da8798fe253043e7dd77615f8f37414c2d42f68f49dfd74fb49a93de2de4d62a897d511033f90cd7e6a7d30412010d8a480414b9142d9c1bba450da8fd8952ca6be2200ff450b523298ca2674c6523ed9e33c61360a89ff8e27c165ece9916013c918c77d643bc11d0a791925944809234b09b0a3f9c1543a991c50f879ca6694d3757b2d2b3ae4de452df2220df596bf3366555b91a6e0e4103c249f32e4e6615dac20f245a84cd3c4b69d666478806962f9cfb5fb5a4d032f0a809e2cfb52b097280396ea20168dbee1e922a514139152da2e21eeefb17b9d641a95b72c497c39bc7ce219fc8653b87578341b42a53903193b724dfd635a69dce4e618501c92b51dfe27ba98bf8101e83664e171de535b41e93ebb508405e50ad8ddd47f8133eef3474a751cc29796eb44eaa67e48e8db7f2af18f315b3184464832533f2583653b5b3d9728a3118b7de89e3f06edd4a7bcbfd596ad6c71886ec16fe01a42706b5eb18da58abc307819afbe4dd294c1297862f32472b227f6c09db4564febd4ec98d74ef183e365eeaea452c4965a73c9c51f452f8e460fde8194826db416291bf7087d64b38ddd485e3d102aa11c6bafdbca57377b3e4b40617374d50e2cc2adb074a423701e3ed21561d8d59514eb3c7abf243c688b53bcad600f577faf20c23c30e1580eb4ffc58cba38615d3184adea1d68b4f61eeb478644b661497a784e13afb6935c48a9c054437eeb92fd02e852957ddedd8efec14ce61bf4a3c74a701408ca9598a42dc2b23a2e00a4347cf66b8b2b861f696af631e6b52294ed8d5ad55dbc6ddf301ba55da1c3b92fff0c5ff032a43d9dedda8e43f9e28c4280988f80f5a9fc243df4384be9c9694db84a66a3ce55883f4c38b593363bb5b27fe37803e074919edabe4d598e73a661ace577312134fe4afac46dc780dc46b5ca930da229883acefd4d036e26f4f0601d198fa1b05188f59d9c020a1121c574e3455e96dfbff0d99fd5221bde5445941f603ece805aa20d43528fda1bbeac851530f0812a596f837b556e1517b7fdb725b90b684e1752bc9ad1f172dac49924d81002baa0b1584f9f02cf1ebd3facffc58d57da6cbeb110ad50b879a02cd04231921295edaeb20bad9b6f5526933a119c55e303172745a797e279a87b5e734d3f33a14102b8c1db63d2c6296165fffe0fb6a72c1189178dad1f2044218f08ce6738e53b76abbfde12003fbcea63751701c47767a5e7509854c4002ee161a6446d451cc8e74a8f72cf116e70b37f7a167633e3e297cb449bebfd549cd6c5215458b918e733fe1bbbad3ceb9778f1a7389589f99f3335f924ae19218d2f41370b1167dd9a2e2857212eee902115e64b464a816b85d6b53c36b01d93874c2561a6f17f6629467202aaea;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h23ca842b68672a2822bf9c731de0bc055a6d4063c7b3988dd238fcc1ed4c86071981584e178268b450b8151d125b0bfca231edeb4c662cdaad4c69a7a15fc8a15270499c1c3d16cd9b17a64944106dc67107516684220fe29b2648fbf84d53be76f1011cabdc2b3fe37fa47d6f9f46e806e5080af892a83fde12d350e3a0381b0a842436a29f2835f0851811329abdfc9ec20caf70b386c6515f73f3d5efa52b27b3fdf02d7ecbb886bb3fc0dbed9d9e6a64b14b36d1d6457386ab655faaf589e5c640d6010b3114d3f5918248a38f6ad3fc2f1f762bd7a7bfbfa0877cb3593e8830db5ed0a6f69103136110e4ca82a9181295ec7f32af6eaef2ff4339e622038433b004300daff48ce01c5e37aab7c79e4f852ecf1d19f90a169b3df8e5fa928cc91c248ea2a97c3a96ceaf9aafeed3f587417517eeb18d83a324c54d63b4084479b3296e5613f89ce46ec32755b2953af8e8c06da185daeabb5405d938c8c56891ac0b7375f7980fe8f4eaccbe9ef1f72c25b0945ea7f39a26839b9242ce667d4edeb8e566bec3c9ee10f95d599d71e23b272f3a53eec364877ec5978cf70c1a5dd57b71a44f45d0e014a2facad375138049786cefecf790f5e87002f8e33f66f3a18975fffb96cd0fcb42696f88b9847dea0b7109ca1ee3ed974b5f4a957f187b364ab9c860c5c6bb414436eb9e49877c88644991f4580f8718b1ac3885c190eaf24e8f8668f6e6c3ab94af5032a6613b99f26f34b4b82ea023f122a6d270e341252bb28f2d0e1ce07ce26ff6915ae2b41590af5c1f46f5e9f1f1e08101bfab9eeccb3e45d3c9e1568e2c084719a75dcdfeae8fb110ddc64a2c5bec927cb8d4485bc3103ad4c4e292ce7f11d960e3b8842c8867a4dda2f0541df8de6582d2229f118e33ffcce1495f8daec44c32d998fe937638343b26682abc89ecf2882566041dcdd0744ffe707dc3e7be4d2cf55390241ee2191cf858d115d9f8deefa8b678e7e411083ee530aff33ab37fc094f2298b58f76bdf18860e613d704dafb3430350b90faee97fd9c55d9c4f4f10d70f6e9662954689b0c7e996f3b257b1a81d470847ab5039c8fb8f10017a60fc6bf4d867fe02e84891ba89cb4c6f7ad367c9c6a04f599511213250c59753a119a4f76df372eb0126ebc3d0a7b6927e0495e71dd8b34de0e4b39e20a3831b724de39379aaf6eaac84d5f1e31b9cc87c6489731a8b145a015b27dda9401c039713e3a77735a7420b26c502c214fa4663819dd31b5ffc9f0a208c2b0c464a6027fdcaf44fadbce57e84e073708fc9f1dbbba5ef36e394b5beb6c9ded22986e815168ee66133c441018cb7221935df9d17cf72f81496450a6955fa658933b788427e801b574847962d594ebbecf1bb67e5fa42150c465faeffd4ac2b8e3a7fdce2b0c78f401d60ddee46c47f413c8c95ecbd785112431ed69130f27263529457e385ca7d8aaf8b2c4b3bb9d63fe083267d20184fc9cbc9dd8edbbafe6ff69f3cfaa40eaf2b57d73733bea6d633998c1a6eca9f87472ec97e9b33e7e43c6bfdfdd5789b2016e0ac1d8a50590b40099f541ab519fff1cad24d97acd538e046e56d02ab03ed4de4430125f2f5e1a9d0fcb60a9c9f1d72744c0ba8bbcc84fb931ea9a81cd6f71518ddbe466e2a66dac669f99dbd1b7ad22ec8778af2700697783ff3cb8881ceb5acf0292ee2f9a097f12fe8eca12540fbbc20497762d70a58cdc454bd1e261eed0fcd8e603425c40b93f24b4e66ec5b1b4c1ca0af65dccb46bee7842fead3679aa4e8e119fbc128b03c46c14edb0a40e717390415e108436ac0d2d89321b4ae372a72ed56f71d3ce28da48b3ca97ae729716c87eb84cf69a12aa9248c0211204d0bb1b50d25b11e484b89af275ce3045a5feb540ac7dd4124088aa2a893f39dcff7a913d5c44494eeed0e0d99c6509c24793cf55d30d16ef0ae5d106076481d548e694c896cdf2a23a22391c40ebcd366aff5c5a23310fef3656ab9b4d314c41b94ff18fe254648de256830490d27b6ce314b471d407d6b2a991dda0af731219200dc899be8df3d9adae2d9ad9b434b75fcf09abe179765faf19c6be0a289a6d4774d92200f528a467751b16d801296c0f8227a3ddea0442be20d5a9b1b57247de019250f7494ffe14a2b7cd3b775fcf7a1743771dbd31a3cddf764a83d3a74825527240f8ba60771120dd85f4c012bc6575251ea8f69e7747414a43df8a175a39a042dc63415ed3488c51c1777a400e1073fa8013a1b99726d1e903e0f4b59e88814b49f2ce43e4bf8b9cd0a131dc57e02533c6a948d093e86b7598bc864309fe75f473371a2fdd500db746ed4f0eb5b8619c7ef7ff47444d17a4079e0b710d0b1546ec4e2a8e987d450bbe4a0192174f5e15e52ac238683df4e71ec7779b5d2175a8acb7313716a3cc0529ae1d088718867e534f97ffe0dd23060146ae57e2f48482cca4f1b4d73fdef0fd8ae9e080673f7c5dc1d653edb1df7e357a99825ecdec5ebab02bdbb52f673217b61d233895f674fce5ebec34e63e43d655d1cd02c492b17e62ce1ce16b54842bc2c76f81dfee4cff175a1207982d07ac40661afec82f3dc2d6d6005e82eef2eab554e9615fd30095be612b55240b38db306e5aecc32ea0df014b315e7f94cba43f5d59bec65ed6f7fcf9b8b850ead0aa02a484e21f26e81d3268e47ba19d7f03b59d8efa6a631deb7cbef2f6db729ff058e76b5b84a05756b10ba18e166b1d30d9dba336c937fa2c43833c113c50f9e756554481e7af7928d2f0a49506460470b2e530dbaf8bc769db5441d36e094c0a90ba2535bc78b3d95cbca6ed8811b8b711f52de4c4d3e990c5dab81932f6faf8bb7b60a67f6d76b7cbb0e8c9671c7ce9ce1c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h402d7fc8268b6af78eeb6f5ff5575557aab49478790e81f30c26dfb402f6d2b745a81346f59ba2daa458992e58543ca7775d094d0be47fe945a8bb207f9478b026ed93ab3b382a6318dd1be74c6fb588eb307c17464280a8a166d06c2e4045cb03a3ea26b5af8715571fbb3e2744e5b0ea9e6b6f74ca68bf6315429fc957b3499a68ca8ba8f769711eeda58977843b70df48d862665cb174db47ba4e19f6334c5e52fb768fb9d19dd18e639be52a6020f9dab06577030c2e92c6771ec10212763b6a59e65e0e48aa7d2c41e785c243debce82352b1a9c5a0a27a704343fe41e4bbe2fe75afc65b7cca38fb76e2a792c9b5db9931b2517dde7bab021fcc4e0aa7e2a2ed612fb79aff22a2d8b4cb56311183fae29db412b905045adf5c2f33135d3a6ec877b41df09b5f1d35b2d98475771f907aa4507fe57201b868009792e5376364237f120a4ee2622e9825afe03ec129ff1455c0963bc0d6e781013cc1350ef5396ad4a21d9438ceaae7e50f3af885fc22a80d6e1319e9362c8b498ff91cf4b3f16e2923987e315bc71c615cd575745ca0bba7dad5ae7fcd4920b77f2517087c13df24d10c525d325afac4c1394f44ca496637c1977aef4fd7344e81b6c5fdec936c07e4a3424eb5fa765d141368c23dcce77d16c6a6b46485ef722dc55ce51f184f6634c60c5686bbd36df8d1d8318bb437b0c7903f0331d36afa2e474a986c87ad0a6ee4554c781ba86b0d8e7f6a722db98e259670e0a8a5234082110bfb7c73874a96b63a5074fc43d5e685f1fc415335a8dc0ba8e35e53f77bc266cc1df5f411677b2cbec654b82a7167ffb0051d60347345ded543c38998b3beb23c1a10d1ff7ff185889f2470a8a49e3a5d31b2f36050ca3a210796855e566cb7ec5286cc835840e06311927a3f1d81705593b46c69db710ccae960b601919287d81d77b93ade14ad1cd754f494c7ae227eddfb50f6bbaa8c74b61ae5623c1f9d43659e9c07ba4812951cc43e36809b9456097c0a1cbb1a9a0c452f49fdc0df8ec7feb429707be0629d0067526b9ab02f2d0faf74fa5a8314d14a5d7daf6810cf53f475b5c1ccca444ebc264b44271e4a55dd52ed807158f179d483d9fb600e687826b75c8af8b01110a13d389518233874fe8f0159eb784cdb4c48e287d5a1afb48a372957d2bf49c37cd9c1511eab677a85ed3acab6e6405e3854bfc1fbd21b83f3ee820bc9f3a6b13720d746caa3d5acdfc1fb2893d635269caad4e60a8634b3e71ed4ec497a6ed015730f27fe8d94088d9ba55be9a8ab7087750381f520dca52292b48a0a9e9b0b0383d0064570637389879621857c2809f0a64798df981e77d36f338aca124d5d54908afc866c3331cfc2553f0770a12c8be92dbec09fd9ec75fccab6482704d0701f5b207f76e8323faa9e28066c68e8cc9239772b73de1fa13b5de38fcb691c60240d19fb635f86a290df28f7b9c97cf1a7d0b38e6a092b41226acc648b231f102cc212115875c511b05cb3512fb2c36bd00afcee3cdd67d248bfe6a525c7a102c5ac347fc52013b23862399b837ee63a996a53fd2f6a71c408b49af9a89d1519f57e40248d0bb2fbeca87536918603f21856ad63e68d22db0bd43824cef11047ba25f3de68215a5e9157358b6dd214fb6411eedc777e234d149f9e0dcb74d4697d2b41cdff3ebbe61c7634d58e5e3c2141633e5aea395f11c9a67a55592f70481759c5e2f9fd54e16ee4bff0c76f5004f0a4cbc8dff5ac694c9634175acdca94500450fe4c1dc97b46ac6391b13b7f199c7ea227638e2faec931034b70c2114e67db5a9dceeabed5772e4355890f3d5182a0cb1ee24e5375a077fd07329538f8e2a900581159cac979782ffd91fd69d38202bc2e35c4b4e6d39792f7241fc19f261237efe18424e0bb87c84e8b2eb4711059e9a3e5034e631c529a3f2fc000ef3730e3757c1dbf7fb277de8412790bdf1f25a4d892bd3e8a7cfa84bdc84b498e0abbc3c9540fe4cbfceb0507d16dd73d4c30723e6b02ebd3d469d5726c47b04c78b4f4fdd6be7f4ac1453a711bedc7005af1b6102fb8f29f3a31a6928f4b9408ac65c0d0831b20861d966ee1c4b224c07ec3c2699a4933c9232c6df71d937a7b94b2399fb3de6f1487a78b128a4c9d2a4ecd1d2a74841f85888e237a4a7e7ec8d35cc8fa34cd0eb82ab127e572763d2602958f0895313192a22086d442495da20e1fc9429c49ea31b835dcb12dcd43a073ad79ca463ed0e63aef0e2c440c94774cc3c3ae198cb63362036319b4d41e2b041f48a2e8c7b499492d3ddd2968b8693630f15cb3853b6776c96b71ded7a3b8b99d745faaebd1f8ad643dfcaab7612067cbecf99b97328c1c974d90e05167c86291b16ff1b27d9cecd09884a5f5976814c718f03d9803d716293e4e2ce91afa4fe8186559b685aea76744d133c23ef5161e9e3352ad9480865ebb23edcfb96cec55d64931142e74d092b370be0b6e9950502003aa68e9eeefbe83e507abe499e58319ea6aa2818a3bd2b635b5a2874aa2520430a1b146f9a35c4629c86e841160051a3fe09acba9033346fb85cca40075002c90aec9fb947e8bd5ee035e891e81cd8b8eb12efe04c7a58288bcd32ef389a0a2ca790579cb4be0456914ff9dc2dcc72e21559c1c2a4199c6eee7ed88d637f104a43eab062a516d646a93b62c63be214d098378412106c69aaac455f035394f16d94702b57de9f79c670929560a61f1c6096329eccd98e2fdf16008be0699350190ffb84df7c82351b22ec791759d5c1eda8dd3afaa182b1922faad330ff67fbc9d13dd8693fb183cf7247f16b01e11fbce44668b81df7e5b13776b9b74a3adfd29b78789a2e14faefda2dbc4e920088523313ec73d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hbf10f686a3d70397495b32d3f318cdff1f5bef5dfa36fd7b5a4ec0cbd77ca05a5420a159a2f920f87991a6ce146e349c794b560f0e9e1d07fa794976f01a3242f483bd9135193501a93cb873715e12568d0c66cb5a0f1b724138135f9113adc6b4ea4fb5eb7b9f7e789a41a67b1bb0b02cd475bedc9660766dd29968a5208b9fb04e9f0e4768a96adf87375417782df8ce6a105b44ab5b87d72414caeb92808d07623e070f26590faa0d4bdee5d5f0b95790e8448b49ff05ace0e9f13380abd76b5bb5988be5b27b1d8a3ada9cea646781cc39b37798314865a46848b148a6a91540bee7aa2a6d212b0c8d36c62ac46acd6febd57b644dbeacf6210fa20ccb7524134b558ffcf6618207b27a58951db293ae791695361170c580e3f8c73946495503c1f6138b978ed0b57169025ec4040390f573a4029929e89830451f8684ca9525d7a17c87a882b59b3ccfb57e3a62f9f342d08915bddc7e0355026eee411650a3f130377ef7f46d7c4c54db0d22f5257e2235e4fc812c0a238ac0f587347d97d1b815b199c5d8754afadab06a07d5adaf77d873b060b53c86732a82071469b5314414c9074de9ab142cd14335cd4caadc6ac31f9615a0c72bdc9cb65aaccd1d7c30793cd841e2eed160d36242090a52bd7891d9283408ef457786f413e7a2175b1b36dfbc7be9b189cd51be9a26133df81545793bf3dc9b62d9bd01f363780e5aa656425f9d44e92c7b6553af59f405242a37291801fec158656d6e39ab4d3b598e2804fda1b0b4c3e3fb72be8afbc199c113cb6ada97c316c70081224037ced37722d461c9953bbe3f867146074fbb90cf8bdedc2a10c869dd12691468ff6cdc519d81694be1701e336d69e98fccfd5fd0f2856f19d89e9cdb604823b774991019adada065e3ba15dd0881f5843c8f1a1f02a2e4fbe991e9a3367822d6e6103173100852caaa6dd6cb388bb1059481c301b9a539c9fee9bbe514615a6d3baf07cfe0b4965e72c6d039e561f4e710363cd97c2fdef48acaeb154ed67b98d425a0daeefce744aad1b272de1c5f5bb64c970500b1a3bb1dacae9eb21eefd856d8ed3e5223504092f0a858f6412a3e6ae7673b8ea744f1d60997842f3dc4b83104a929893c56362f3d9acf906a7aef68720d193d9cd0343b1c107f34cb003f9446fb93a7a342be40dbc9ec9038c29726adfece75009d27a9401fa4af8108684c00b8758400c36014a882db9e605cf5b34fb57804ce4ca04a4d4e98b1742975bc30e40ae878ea5d0dc13420ecd237d30a4d3f6e5d9dfd8eb384e7641a27e666c4be3852dd6f73eccdbf662d0eeda7591405cd93a34b26bd2d8dc04a92841b569a47d99454dc55fa2332d9f9e17e2b9b7c6230a857a6108c614046d5c3eb681806b8bc636a4ea99bc06738c57a57999614d9ecb27f12beb589e6b459305c123acea68937c314d1e95a8255ea9d9c5980bd108d48e862208ca48b7fffd31484fdead6304b90c63ba84acd034fbbb6f53df2487a733eab93857f614fcd86377536df6d0e5c643124ddb0fb317935ee0da9aa088d1173e301f754bd49f0eb0cfbec663908914aa40d70a4423c0ca0159f349c1a2eb3e0c830233e157d730a5ec223845dfbc052bb6643c6ad3d1d283691df71aa2ce85c681895bc33cd1f39e2c68a4f804fcf7c678a7185ce17aeb6033c2bb9faa8c1ff425ecc7a0af1347ef2eaad682520bc29aa9b148f7bb7e272dc4158c83e7eb4e274ef3f2b3e581e02206f322529233226131cfc76af3df14232e48bc7f5fbe4cefde6003db07b13a3b8b7d67e14f37fb4d37c19ae95ab2afdfea6b72819de1b8cede1ec2f4398ec818457705c1399cabe5e422cf1087685d40648804ea2c0c044763d6f37e382d459f48fad1472b6af32a1fab18dd2e436951c03a93d06e50b9d5afca1e7834aa8031088b76a0ce914adc26a578202b6af5d760e1e5df572bd997d5205501b8045738b9604fd46d68ea73999ad7944efdee51b2ed3e4fadc802f47feedbbd7dc4978680cc64e618046c752ea1030102c20b153f1dc8c2ff195ba535b262e667b5118bc9e78189f6529368219195d1ba076d9b1ee0edaaccd98a497087354ee2c84ad7cbec1fbb525324418ebf12f45cc5b6357c302a0a4b7ea0ed11a0bb8d623b35be21d2704c16d5d943e3cbed13773d0e3c3f2c1851cd54b167132244139b87de3d475b6c6dc67c29d43534a2a7e08bad80e834688bfc5aafbd1f565703545a23dcab3a7552c1f27c729d01f3f7abbfb3902a343c19286529a591e6a9fcb395bfb2c66673f7e0f706909f277bbe41155d4f2d56e09cce6d09e4153460dcb5cfe3e8df30e362d5b418606cbe4475c743df62fd7efe1b6c4608101c6c35c292338f27360e0c3ea9151da4d2c1a7b066fbfe3f3cef3a7e3f6ed065c9533fcb33ccc71883518da2ea5378b9698e47615f0a910052d2b1451e097f76d91fadd4f5af1dfdbe922471ae7f52b875eed9c5b6df5260e7b5f3d9c94dc3176d6c05d54bc41bb46180a18c1124b756b954c43fc5f2396f1b19115a3aeb3d33801a322cadc1cabbf2679fdab12dbd92846789b35210f8676c25ed43170385e15ee11603b81916409bf891c89731b3cd14d4524fd6a764b5175b2d4a8023c27fa569c7d2a699e2998141242ea3ca86b9f6cc48095bc38af1054992ab75b0cbe0ce9595c4dd050cb8d006a98fea436dc264ee7c816b907ca9c37fc3f320bc8c2c3fa7acc856213157c71b7f8080be78131bab0829da1668d0fc1d1fbf1246c6c3f0a450d7be1ad12e114607a26f285a460adc412903690a6f5dbf2c19a2138d6a7793e018efa675942d9cdb438520fca10bcaaa7afff2e0a3af9582e74f858f885cdcdb545bf228ceddab433;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h232004414716457a1860a05869ea386f92e273ba49f056150c8db0faeb8b41f9c8e6271dd3d0a20c8277fe486da74708b7d966f48bbd2c6b78fcc11455f784a5049f647c69123096ce30888edc1fb1637501fa30c0d8f57922930c48a0c2c34709225298b33f88bdec616597a4149fe696c580323ec83b577d27acef45232cd40348b75ab5cae8773ec02a5a427adf1c2ec9f17aaefe3bca9addd9c341bb64de51995e01806a032491feaf827e696970658d78558cd83b410af03c1ebbf040efcd3859309bcaa264c3a904ab6b712f14f4749f5526f90636c04be944237ce83f80caef8aa1414af5778a253eb07e6e20f7d5c186e9b4576390c9482e761017f3011ac005f6d472cc59e0bba79c6d0aef730633640a9201d257f8bc7f335e67dc50d0b2a61410d5828dd420eecdbe1d46d0dc8d8adc3bc45c8b161badd3e3b660843a7db5163a7b3e964bafe64eab74467d971fcd739202426c32313c1c40e3daf20f42be1ea0e6095d9f415cbe28afbc633f6defde4874c181a5730860e918aee0297bd79ae383706f9ea5efbff1dedb3ce78fcfab8acae6fa9c220a7597888038780637e470f955329a0a47d338931cd274ace48302dbf5dc8d062b21b0d8f485a9257b1827822459f7a1ab56ee29cd59a6d056b1b54f82edd31d5946a64713814abe5ea0bf615c47ff92549ec61c4afbf9ab247b62d8467328bc0895916827f0d9753d7e7bb9490f304150617a05770ced7eb6f8b3b5e5955c62c39c7cd329ce82e494259d999d3a73005925210804570b89e5bd17c2d3d7ed7845dfa10b3558fc33ef8d84674038d1b53d1606e535238ff2620a6b9bafa25336f92b627b2dedf38750d18381beeb1e286eeebe4f013db7161aedc30d1391bbeb840243fe79f344728df6e2d8578778ab3e3e279b67b19c5db0ba8a9da517b24c990c40cd73ab4ae0cbd5ff2e2ae7538ad012301d593214d7a23776381dd8007a9419eef1c1636597fcc3e0f8abd763aacd20e2ff2112877327588bd5841780d3873710627be204e2706a1748c44585882568593ed0e21fe6df6361952099ef1265e192791430544fcbffd7345edeb704acc652c9985aaf9dce7f6050f0b921dc346249c7789bfeee784e9d4f9db2a313a0f96aeb9a95ff0f94490631840960253feceac0fea74d59d9956bf18bb3464c628560a646e37e0445937bf3b3b163bd38198f688e10c06344ca3b16490f8dae4278ea6f42fe584076256c7092661d82609125521531609a5a32c3c642175be04e76616a476c89a16ca626e1f3c04be7099639008aee1ac32d0b30b2f867eef4e41d0784f366e8d0198c6d388413adda6e86a060dddc3c57358b0db9ce7c8e1073374b80e9d88f6850e4e3650a64aeb3bd5b6bdea3630c7dfae1894ffe8489a8d5b32edf23bb69419f0997d9ea99162c78d43d70247e826676eb07e1b525e920090c46254264daaad5d6bae387bb08b09a0d04bcd0c3ae76417982ce74847e7764c090c0547154472e39774bf1f560a196465e083c49800aaa284cdba2eeb4a68d75767229ab20e8baf1910b87810b70d7aad409a9e76681b9611c6100496105ea9c3e5274695ddb19dd0211a396b3375879956ea4ae8744d4e81bbf17af698f3aa45814227c2aac83899461dc490510b4fba9e931570979eb36a05d749af79d7405c339c527b0887d14e908ae12ace0f7bf27f51de581ae49ae65fa278ccdbcd84dd092c752e6c1ca45bcce3a67891c7b10d83eb163e6808d4bf902347a1e373740a3c46c017b59ea1cb036bb42df9354404c0474eb6a32553b18c53481af8780969f6832d36abf2a8bdfd2fa8a20c33992668ed0170dc8ea3b892f9f35e3007e6a4368318bff879b287316ea84a5b6d50cbb3fbbb66e13e83570b360dee99e7d1981cd494a173ef167b767d2ca26ad8916fca06c6012497b31b6e596c4b6a1334bbc6f01c71e3e7b2f1bf26915d7cc9ef410be18df061c09cc19b3769811121f7bbd38267c8a9154cfe99f8cff401f4e8f58c6301c090eadd57cd5b4c47e04ef3ad15712edbe78d985c30bb52292b48f177e265d9e53e7d670615f221b66d931e82f43fd2179bad6595b6f345dbd0a787b99ceb249b03edc147cf4dc0bf1e9960d7a66676934dcca36890db9a1617aa98d58781de621c2f325d4d6f4ef058eb8501fc6f6a5eb0c05e40b251d18c698d4ade86019328a0e436d6ed864bc840954da37693e795bb52e3a65187215fef5b0c3df58a65744da2c5919034cb3988f51d1b1ad7709d485d17df93fbe04dcc9bf0b4b076523b8e03578f5487ad5811cbc4901894e3e8ee05ace3e2704a0eb620b48ab0d0503cf2f7ea6166f0aca24eef76443164bcbe8eaa194bbbaf0d3ccf1a965b845c4248b03bb3960318de1a4ae9b94eadb0b3c306108438af929ca9dad89b916291dc4ccc5bdb1ba440626fe4870bdec71becef9872f5aeb86283baa6fdf82fb810367da1884d5f8716e87f3f64e29d89c422be8b6e81c46d15e53eb1508cdfbd5b43ca605a5615b80d5baeac5b65186cb2c17f837a490487fe692a9dec2f60b992003f3cc302afb08068e69ec5f9207b4f700f699d5c42d266ce73ac9dc3e214b30e7c7c28b15f6c2e41381f0a66733faa046012086f37ebb6975df92009e2d677e68eaa806668f1fc2768b6649e2685ae5e0579984b04a6146d0a418d3e6c2ab8f03d8c8fe6477977472def387bd6e797add0e17f0ef81d37c9087067841a73bf0a00922ebb2b9989360572ac9d956856a566e8b670962a0a9f7c2bd41d4b23705fc50170ef8f84bc56b94c3f97b911b84e44e33b2512d7874c880b5f8363aa03c356121416262ae77a47a9e563d991623a8e5d5b13bb7e803c58e3c13fcbb9c4c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h3654277b42ca3c5217db26e5652ea93451afba3ffcfdd673eb3f1dae8a5d140bcd4bf2e45e4f76b64beeb789d4fe9f7722856803a1bd3ddfa7c66668424de768984bbf83e1a3fa1d40e18aa236f73cc7d5e9ee97a0fd9de4f3f6787582180d23fb132032f74101345bf1d166f0332e10a6258934cb027545f7cf66b88fa599114d7eda06fead82ff518b9f4e0975e2ca2803a168710fc4af20631768020af362f619feea78db7033b66e14ebf99f74e321408d4d887f37758858c9dcf80526a4542f3d6f91f0b4b25d279242f6e09fb411054bc7d64a9f639337004271e9376f7e735ca285f6e1bae0f2275c47dcb961df44685932799ad39f7d54b8b85c294bef13b6e25b37ae52da339e41bb1494930b854bfa54514500284543286ad7b949d1b827b3ed6baac9680876e592cdf334ec935398910160b04ebf5df9fc7c615cbb8f83edaa3cf42df4eda407402e006ab9e11cecfaf6fe50914e2897b71bb3948cf2b94dddc7645b6343c6de725b3f8101063ee5464f7dc7bf683a4101cce1deeec7b8ca70a59e98661f3ed928c06077550333674373c0f42ed0da0df02f46bbc2219e478c2ee18fd7447362f4568e419e5bb23ea7de503aecdd5fa3d818dcac20448a622b02493e805340da58d50dd918f477e762a92b6da18c5c2ae4426ab8b8bc613089f32b4033be72ff19d17290e18b96273541a416fee8654a824a6605bb38e436498bd8f38334dfed3d2cdc1ce62441b5e0972b98f9143eaf723486fef6f3d01cb5ba294f148700d3047417e0e014796daaef5e8fee1f2b1f67c60413e99026a1db2a387edfd1990572cf1be4f85233cb7c281efdf1f06cf793e48fb91d8be843f5200c862d17e112146a8cfaeab210e8dc10746545d4987bf69366095661ec46443bb57158ed658b5550e1bc7e4697decd7dbda1fe1fdfb520ed34760b5dc316d07f5a3db57e4415108b07dd3b6e72112f65a0caec13ea2de1124827e7c49682366bb5bae3f8087418d9d2e746fdc34749e83c0c17e0968fad37d5d7a1316c3d5541e8c015868d32057bc3db26c65e3364c8f7a3b4f28a0be14c7375b1fa1eb3bf4d2cd48fb66cd637491445f5f2d39402d3530c1db7bdee16083907285a137ddcc127aae9ca92e6d900f8ac7daccbe593fe8b6c0f860e3e6ed0e7f86c65031abda2b28df0380a86ae21f8dd1f3cf877e6a3ffdef761997c974f261f626c430d04358e57a8548da0f0fab33411ff7bad8b973e41295655a2aa0f3b94d6a6742d01e3981a9bc496443412ff6eed818e856b8c4af1111b8a269881261fc345da26e996869270f6c296243b72ee4167a3e89be8cd8e3e6f7daadf250b37c93066c1f566ccad2831bb388d100f7d1621119ce458b280f3981e7e2bcb0018584510578cbb9820b854435dc098681a0a959c934a05f381403e23a7b6b71b32349b9b05dfb18b747fe936496f78cc91ffc5dcc2dcc9daf666202606b0c6efd4091652bac3a107d14c1f94740534a11e6540c7a61c3ce969da1c0625466795904b56c121bc5c35a6da3c8ddb7030ab1d404367eaab9a9dc344df4d45213ceff02b1f86882c8c42877ecad9ad882d38cff62b77f50b6689bce923bf7dacdb3975f8d92498b2145bb1005f6dab843caf636f04b403e325eb9fef150433af141d5d6d8c54bbb4786b2d98ccd8d5f88eaa44a00316c56d83d3f642d18b1adeed17ece754dec65a9176971b453727d322d3002269aa8012aac9f91c2fda7f47bd0ff2576ca83050aaa41ceab1cb6a43576e9a6c360a1bb8679594fadc6a7448422679027a762a7475853350eeb534d826df01cdc4686b477e5b4dc27e71b9abc3e507c83931606e0e25be9633cdca9cafcc1dbfcd960805aefc2b83a2101f5f08c9b3c4a8f9125e44e1bcbb94a8ebd39ef7ee7785f031b01cd201a2e53fe5aad5cda316730d3dad3c46e81430fb50bf75ef8f6ceec185f4fee2f3566c3465010c68003081dd7678ce68d2671b975e8c6ad2a9cc417132f376ff605d9168f54a7aec43f75b517fcd9da0744793290e9c7bba75683e131ba59aa701e10a2538e78834f82f6fab52ae3728bebe494b3ee4840dbafbe32f50417ff7c5476c737f636f283469d73c6bdfcab301918e193ef0b65d69b53bd24132bf3864781efaeda44914abee6c1cc2acaf26115881865bd815657500f6e057625757c0cefd368697a17e7e1751e19073f38177a845d56d096d6e90418fff86966f08e1d4467b8dfda2a4fbaf2913edc85387539d735c8ec8b7fc6d0d911364c034ca7df2f79bed11593cde66cb645ed475bfee89c1b1765896ce6e03c1424d26001f87ed9131c64837c82b6d8e64e81126a7f6309071812c995ec56859c17be2d90110163e99475cd66ee8bee8a552db209a320af924d16abac54919ce0a6a4296e90b71846a683e1da3d16d164ff4c003294c98e5877e9e5d73ec86dd8fa1476e22d458e3dc146f2b6f4773ccec464bdd5ae21a09dc088b6045d6e62306ff92f80ddf70bcab92bec597605c996fdbe79738e98b5e5572107e262c6286ce80aaba6cab7085bc55e1be08a9516ec99dce08e391b495bfc5be6b1fa43d3360db81ad7ef623a18e7c67d1e7ca5d55bb562e5f13789cec7b9b7c09f7ba6843ef6a3608d952e538c94f69ea65eacbae3a59b8a583439f58e6872c9838af3b56bea8bca45a3f00e9e5fa0d16fb8b9891d73eab9b805cb1f59ec0e928dabcbff6e224c2af3cf08883cd3bb56b0cd4c8391eb17f84d92b3bb12938059fbad3e458f305f1f1815784cd7c0882ca53717105acfbafd779d466e8ec37bf4d9c562c2599941b4a3cfb94c0bda1af6a2f950e01419da5ff9a7295e66909ebffe082eda5faf57b2fc1e4dc77218617ebb4b6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5979bd3155d76d39e2729763fb15e5576a393d95d6388817a086a40a93d036b01fdb23f9ce4026a77f13079218761db8e981e0de7bf501851920e195709e7eecac179fd859da731e014dd3ac4358bbdcccb9b0d1f5d5717a24426fe31f73061f289eceb5df8adc4377b582b5bd7cc9bd020fd1752344ae31f9993b253f2e4b2cc85ac31c618604e201b23b77078b758e8fd8eb38f9b2dbd88f020c00991c6367ba2484bace4ca0c353c2e4f719b9dc9d0016bf15c8c9837302667552d70b0f15c03d2c0c3d2544845b685addde540dec42e3f2802ae56bbedf9d6a13da90fa2474f7174fbe93b3a34f909c1442c4542172d3a57049c9641b2c0655328da6150824cea386bb8e7b4a973f7d96d41cdc52df263496dfbecdcce0aebfd466d4452a7d069ca41553262cc7dfb167f37325417c2a8a9ea7e450b6afbca3fa8ac6dbe9a5fefd4d87a7250391ef2428ddbbe7b017bdaeaaf8f4aeb9dd9b71748a97d7eb23c2cbb85856533c4f5f102a30ae5346a3adef15865869bfff6dd4150a552eb173b988b2835165e28e2605193f2dabdeefa6cc7b20d8c2807f0bb8f4c204bd219d6ac78d7551a42d60c21743c1ea7d98a5ae28b67f9a949e4c1682d438210bbda69716d011ba4a8af82aefbf5edf7b2d80dfdd4e981fb5a899d9ab1501595f852807dd4766ad045176686a31e70a69b4ab5c3601007ca8434d00ebee5854824e99910b5c8cab90704306cdcaa8fee3a38552809e605f59a13b3c4a83ff4a78a94ff7507907643e14ed720bef8df183b3663f3ff1c443e1520cbe0eabdb86593a796294c1ce3fdf93a1262b8982b098eb53be26470535e0d01a54703cadbb1c9157c6efb4f395d3fb612870b9c8f64539a4f9fdf78afc7eb3a32456e63744701db345dcc7f60938b4979fd22309f93f677c5888bac12fac99e454c1760879b651470e203597939e5d14dfd4dcf83fd1c674ffd0de643ae6e541dc8e1c9b63163be6b0a5c6807116dc6f8dde44e34296683acc8923b1b191952031f4fb2dd3844353f7a96051e29150a5d92a06139702657515649629df09510d09bdc28de49f58ea0982fb20fcbe98234578e09769a45249b7a6ffc1a0ee7774d49040e412aa48682eb9d956fd7221efaa1f33caa6ebdfc701213a2db2d3f385feb5d6cf2e4c5b499ccad4bfab534ddb70f44e04981b2d89f32f431820838f53287fbd34b7959e99f7cc06e48d5425c9c313a9587a6b2920ad4a6829dae06f812041e5e99dc6d59f7e9c8a9958c513cd93d8b6248127ba18c806031200927cbd5565266f7e4bf7d859f0cd1602e810646251d155a8e2efc5a2e28d0d809310533eb43c367f7eb2a28c88529d11850cc0c5df4eb81ac7381f701844f58054aee54c46ce34c74ccfa05a4a154f696f0518b8a08462a556c27161b44267e7c173ea9b074586d272c67715b445784b391039a7c69e00ed1060188a789bef2740f80da4817ab4c0ba20772663747b39feeb04ac19d0e9c7a37b85562862c5c656613e04cc75690908de8908420743d27fb943f541dca8344ed6f3c5a2b36611b7f48914d1b7e9a003a81633b81551826df6d8f639f12a1fea81ce8286360e9f5b29c1571b463ef0d2ba0b25da34aa77aadbde85928269e4a4cc3ee1e773e72cfc7b8f30ab95cbe76af692981cab649a59c4dff7a0a67136236bd3516a390acf57f5e65200947541cfec76de1e6feaa426f8d5a72de5395c90baba9ba82518a541b28ffb286981064e8e9a5913a9690b74a6ca05c513e8e9d056491c31e0c0fc57882b746e9cdef0db3ab5c276094ae813780218644876ba56834d4504d6e1e314d2dcdfdc3e9f8468510ea8cb3b91c2bce1c4d47247e0fdbc0af485ede44781936429a23b9846ff070349794f73f72b24361a8647b420cbf4f3e50be6acaa7b2b41d1e5e7ca306aeb5e8cb256d0baf2153293b74eabb27682577297d53a0b509da47476eb77d8b316e0760722bb65968a9a78461921bac79e800634719add12bf7fd2796a0aa1b5c816c428984816e7beda1d4d3e69e50610cb91bdf78d1e8c6d8ce5001e776098ef3e94d8babe4a8a63e9f1c8b7e2bd49049471f82316ef6ddb119b11e8abb889c2a224e22f8f7cc2044d709002c0996602ded5d0ce80292e22c8fb9737104fa508bcbd08e45bf3a49c498f4e36276881388c6a05409a6e9cfb7ab1375e78e171e39f41042cc08cb16192f62120ac56f987a1d543d31839101e6083f65491b9cfe383f857b51376fe7218100b136ce8b73ef91ceb0bba7b78d7f045de8d640cc64e0516dcfc6cc2682faefe75853a68214ecd575b6e5218ccd66e4b8e7c38d0e0e5e920a6189012e7bc5213dc816b7398bf704dec3eb8202493dc3866397212c07573aca51d3d17ba85046e8d631d542b4ea3495b11a59314322adce255fd177e84531d55c80d32b3ed22d3b0f56d80fbe6610811af43cf9714f35134d7e0f5500fc64b3b55adadb15639fe714f9870a214de05dc7241c0b71a3a63e9c15e16910eb6be7be19b082e3b659d19bf339052c4d57c373a00b6d38e18453bbba659d847e7635f86d24467b28bbe9dc2792a65c2001bc978d866e90d66cedae26fd75b82338dbb2cd35fb673705e77487ff0a1593129060eb29b531e86774520bca57f20fe1bfba71eaf60dcf04372384f20081881e128823339ab3aee962f44781ed178bf64f9aff1d02e0f165cee3d42025d3033134cc029b72e2223ddbcaafe38d5e6b4284be24a089fa69372e8c55670ba7ab0ffd530ad1a9216d1eaa93a44c8f9d11520e214cc511acefc96588a250d5e685a698402a4a88c7c8a0ecd121b0ab9c67e53bd51469173bd59482b4e2295647dc41912210b8a978385ff65ece33a4fd4da;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h44da81d7d1265091cad620d40018cf1c63985fada78f108be4d5fc013f0c5b4c47b942addf183b36d5a31300f9564b0982caedb1ed25ba8707a8b8d4b188a1506e2639a4f9410fdf53ffe83571694c3faacc7ff8424172aa5f82bed65ab1a29e9e4c229050989a3872376a864a0f8ed156225f5e8a07e70534cc7e8c9a6e40483dcd5b47504853114e047f8161899208816123df1cf8703a6730fefa166dc312bbad78c87cf262cf408b6b4e8a5f4e5ebb7f3258957c9f9cc3a502be523fe95e9e01913359a43cf1d721272d6532cfbac3b514265274a9165c474639b2695cbdcf27359eb68698f4227367f04727c81ec7762dffb8950548650633d28ca1724c94bf4419b48426c50304f35a2e8bf7c401109377b63d244cc6f0664b01f0a51a06166a9573d050a80ac340d721406adb0de6338e3d0f5c510dc07cfb91ffbec662fa6f44adeec95f514f14ee49aa170313aeb6f1f7fa61177f6b6fd029ef0f48371ce828de10bbbe3642898a6f9734d012140c9da0d60237acc61f2f82dde7130d5d35b08bf37674ca8314bf31ee63f139be0efddf57c28161dcc15b5b8da4c8f1c50ea1fbda32a6c1272fd1639b87fd2e7be17d9865bc977d4c75c2c63644bb18078eeea4a6577ebf21ab82f66f11848f64866135a1dc21f8fbef37c5da108e6c5d948719b72e6c406de49283f72f15a94cf4b0379c86d929ef8467992f6efb848ba0b678564b04d95d25753bc15288f2aec84c2b94549cd4775e95cbec4af82a62ef84a36d6d38144fe50b209716c492cfe0ce971c565824d0036b40b1bd0b874cdae14dc709260710f1188c5ab8eb14e8131537326d1dcab27f947e2be980182cd4b1125ef527cfc93b07ac7f60f45bb5761c9f95e1cebadaafe43d17bc25440b53da0647c4b97da5c76d32e9b7a923dd524a53faddf415ad940960f1ed0427562a1683e4ae95eea458d7b47efc0f400665da1585550315c68bc4c24abd35cc8dea97769e218fe298b1c498c2e0c53e161cfaffe27f5a14cebe96a9a033434e8ba7baaf7a8fc508d63483ebdc58c581ce9c0135c0c499d74ae10a4da5c9f76bdf619eb040d8637b5510547fd9d40a1b477915c6ebc39e52aa079fd797c4553199322f66d0f66818089146173bf9b3a9d18e37f5ebd2c93f94739e0d9c7e777ab77fa642c94a4e5dc72b6b05b227044be2bf1182f7c888b134b82853226481d5b6ac1b3a192e68177fd62c3a60d6ec2c96b435aeb2e7dd19eb2caadf94b857e5f23642239fc235b0de9bfddf5dbb9efd1b9404bb0ade59c16ee1337f107d15eb9144083f839d6105c2d5e808b03a5720caffeb7e5983ddf776bafc7c197459067db5ea26e65e252491c538c4ed46c109174d2749a6e17694d0f87c7ca54427d92e80f6bcf3a66f19737f3519c3305584f1f05fe46d8fd2aa96f85114e88e3cb321fda20516fc4588206933892111be64eae85df43b1002e1be9442d6d5929b5ad30c53eec0389bbeea5cbd5020a4769fc29c3c535cf690f67d3610760afcf5e4092c0af65e20add652e74312d8a4d20fbab3d93d61357fbc7b36f357646eb95201868e457a62a08c20a9c603f89711a7cb77400a9eddf9c8ffaf3dcd5e4a0919875fe123eb9cd966f1baa4d5b4f6e747424fcc82a950cdac8b7c24d78f0dc3b19d8bb1ba825e9f15b9f7fdebce67116a5129da4ab7cb44c0868d779f991fe01be323e3edab79814e469472b96ca6e1c9b17351a075c8dca80aa8b1890804005f5eebfaf8f365b65d5058a8cbde39abc7b8a5720916767ffc84c65bf46d332f85e5ef09eea56e032a4471f3f3bd9d5542c21ff0548c86ecdf573a85c64274cb9d49ffc32f65ece327dcb8dfeb16406e8dd83af6b6a52e85d119891717a1feeee700255c8cc50d08e4e2c80bf7aecc921c26ab87f8be47c61ce22bc54e6b374bfd9f5de3e28bc5f3ad58a999c026f3299207f9dd0b82d48d637805fe43cffa347551ace867afa74595c339f8bad8e39bc9e8b7bd5b1f49dd746180440d3ca89ef3f98ed14166c554554f283767f3866e85ebb9e6ceaac273955c9019f95454b4f90cd2290206da539e17932efb7cd6959ae59c9e8088643e302891bffe7305416918c67a70d6b758333e2b1de31d5afd468d3ad2417afffc37554a25ba128b8158945c0b723121cccaff231e889ba94d5b69aaf511b70842cd1c1bfba32fb2a6c194dfc2762d5348ac48c05bfe0fcc70840ec38fa7ac0550b158a40d7f51c9a09b73873db4cd498444e61159a86fd7af8a95318e5282b9b5aa8fe8bcc4b34d4b851f33ffdfec68fb43a5d253872de5bfb3d5d0604d891892ebe6957352c917ad1b0f4c7062d17a5adb8cc217637c3f365de527542c86704c029df1332227da0bd14e90419d27f7fd39b118d1938bdaa0593f0a7da8794a05a6155b8a1f00e98341ac13eee6731df4ac08fd406a0d79e80a6ddaed1737bd62cebe65a6771066830921a6ab0a6089b7d3be2f3aaaecf34015f56e4b2ba26c5ab70fbdbf9937312d89f90155ecb0e8de52d2ae0db90890cd005d6c9b4cf6b6681c777aaabd4a1493faf520061d2840557d5f7de00ea80d163b986b8c5ea9518541a5811c435596e6582f38ecd775c6ba46976942c6293303e1991bd50ac3c8f8c8e351fdba2ffb384b791599301019ced2d2076799aacfd446d28153a69a81a79cd56128b3112dba6b1cd84b339f9a2b06e5966817637fa08a6ee01798c19786233ba614c38f3505f37b20f82b40e149732b7b018d30e75c7d86ca0a9ee19f6daa493f5bbab9a31028912ea9950dfb7f42e83005dffa2e05fd93dab4fcf8ec254a851fdc61a0dfa52c875c191c37972d643f0741eb80e9fd4a98dc79cc1772827a5ad0efc74f7dba;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h18207db2cafc45e962b770cee42f064cfcb64582575e0bc004e826d96a0d4efc74c8b25bd49d99b0d84d125cf4b04770696daadb2dfdbda493a0a50f91c85373633d9cfda56758c88ea6b4595f5e68c2fcae262b9ba20221b464536cdfdcd00cf18f9ea6bcb0132b97ffc4d5d6849b662aa1f29fe50b0bad4b31068fe4ea0df128b0a92611a40eb5d35ecf67738cae6878e850eb8a43324892c939132ae1032d770a36c144c74839aea4207cc1e63b49d4f8ed5a90509976b36ec1d5db737d4a70f3467dd31eb7615c63ac9390d3ed47b78c830994b89c301b63d03e78de9d86b4ab6ac4b29a4c9d81cdc71391e52703f5821d9868cd6ebaa38421ddec2655f5e26846f875af6ada247a50a7939d71290475afa55ee2a797cf2648290dbfa55db7a198b319c79fc6011ebc497d93caa37a8c99da562bcc73dc0e28615d01a73d80978fdb5370d75419e3f9fd2db3a6253cf010d9e0de768c3690cf5127e43dfbcd1be72eb91d973d677279faa9a23c1181fa3700b5e15e8d9dcbefecce7d82058f4c476a4c99c437b2646dbb8d9d46343b8867116fb21d6cd093e09a03e645e3c194e663044f404445a0707fae6ed8117106c38b34f11e27117a7d95530e57f1afcf9eba82ea3f35e4faba97c2e8f7098c201e62acc4265c36db2d4b5376233d368dfccde44e6ba01304e6dd9bffbbe6a7ebece13816b5fe6e0e84f6cb3c34453e88e8c52607f447df1b500096e3a5f5ac3394d5b49def88ab640cbc3e92998716898801fdbdc7deaf009ab89df661ecb85c3076a5bc677ec12618f51f0da0626625003cb310ddaa80f6bac7cc0cd8d6f054fd9279cc1998d71cd8c713d923c137464e2554813d045323937d48e1a0629df3af88f1c452d77df1798a3876f233c6a3424892216b9ae425f0d05edb01d54bc87904f54b3431c5d5888606162207ddd1b55a880b3ee732ea973a3f4c61f21556da5cda560e1711e170df8926254f7a5ed7c3ce406565390c56a3d285d107bc81eebc5189e8c7036d0d6d4984afdeb1b500b682b0a0934ac2cddf93ec99a200582f77c280713173db4d7b2adbe3dd590a1bb679a92535fb4045440358d4e25d8a16e6b727f4c39683d659d2a1b406dc5f5bd498f271e0e80b27fb23e50101fa6b3192a52744f34d044ee7a9157f0d0fb40ac0068c8fb006751ed7df5afdf7612c00efc06357f9cad9dfa8fdd3798b02060d98f392b471e0007078d31c797b785fbec7600b099fa3c395ad8a3f6a676098b8f65dbe5b084bbc591509daddcf7b5253f133d484db512a47fb94f72fa01b801e6fd65e6f507bae94f09845ceb7b9f03ff2f39806ab758bec4af7d9f799b7a8daf031de0d0b73e3b21acec9c2e4c2009caa1d6f8cd2c0e8641e536e7d1ed9417f3afc753e7e93178706f0f88447731b4188ccfd42918239e85bf3d2523ff8d21a8202eb8355b2fddf2d7f53e444c1b62f442b6d401869f40f82bfb867a23bc4f45003f67d0b917a42a030523a295655db3f4d11cbb4a1cad630d050133fb274a9718466f6a7d55d2cee0eaace9f1ee0452cec7482943ecf5224e9bfa44c745139f5866beb8a118d9e9c9c955ad51c4d481ae247d065c4cf81ee03c99f91017b9cece94a5f3e2987e25d653c9374a91843dc2e1289cf77f357fbd43209f7399ccc4c4055fe950077018f97cc0cb8f94fc8fdf55f01ed565891de65f22cf4708c765b06fa4e76326ea1fc43f93595b805ef5fe37c0d806dada0f484835010a3b9ab83fa364be387ba87a498172daef176e2192fda09daadad244137702a4500eae321f4513eaa696a8ec1bd2c2952ed70d4c4b93fcb598df1f0da36bd63a38474b0d5a8de081717941c8f53aae2b0b51874b20f1c00fd38c487d4c0b86671705d94327a4cd80b00218726a2756be6f24d94b86e9e965ffffb9027fc0c3917a696f5b0d0ead5f71b63e0fcc82f10b3cd30394c8afd6dd8af138a1675ffa1877613c9f5377cde1569aeeca23a47399adc0292f3c644a40a64d363300019a1d305d05e4052c181cd5515239a54d3292db9a69b0d885d2b5581a10ed621c00418bef80036c1e5ace40d33597ab4d426d1e385d02460bf29988173af15222c3f1e21fef9975ca1fe3d515323bbbdd09d7ecb45c309bdf3d206aa2c929856728579c133fc02d8ae2ce1bec6db520dbc125014f17bd6f2a44c8862df52c3dbe90d475fc23e94a14dd6b2d48aff632456704a5c9b31080db63e0203c28ad1d18dba06274c2eef2e610c97eaa9d32f0ece39904b7805e4d3c8e6b007aeaa39f36cdc9e62f3f40d1caabffa389c3f965171aba1b389ffc0b7e345a9124c1c14098c36095793b2d2fa4c020281de7018719b41883413efa032081cbc72074f69b462a9d8151cb86b54644f6bc0896162f12e6aabc1cbef938b5b55227d1ce252b26b02991e3d453e3e80e0966e2799555e1f331117c646ccd3e45af4703d702b47719cf36a018054be3c891a9581d6cc136c3e0ec08f6f60f259de1ef0b99c0e9f716197c56e546847ee4b359ebff0b1bbec817f380132630461fdcf258305fac61df7ed505d6e2468ff44946e6a61fa34cea3901a20cd991c067ee132bf46bb63820b71c1143bb4646639d173eaa7886a6f08c053012301406e6a243b15eec5bf2377c65919605eb79a8b040257b6a82931ed2b1f45534771ef30372466a2e0240c454e92f6268cb61b1b2fc571e7e4b49f6558524e454e2029a4210913007f19e7bad3930e732af044f91290a91fa17215fcb03bfe97f96a8b9267e88fb8100eaeca04d44154ee95e4892ff079a2e32347f45910f6f5d2a02759c90256efc3671ef79977246581e992138e9e0dcd2b96c118e0469fbe7949563650eb3f5ca190401066;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8715cc14c5c309fc3d5426ea3d09e23ec4bf3f603a74e14cf5649ec37a7a919321d93c5660a0d866e3c4da78f088fc76c634fae41987c5f885779ef59c8075b903bb80627b4e3dac99fe1661ba1fff08d2bf89ca6da7dff2a21e1d7a28753e792febb4f79efdf2813aedeab02e12d3937dfbad3050fb82f3262b8f1b46cf316162725659807c123cf3fa9d79b311d0d11692bc650edb9f099690d193788d1cc5517db590d5c03ab97c9d9d23fa1fff24ca492ad6c28dd6649b47afacd6e56ce748f3d4ac9161a23ba488a79fe87881d176cb8c854a52d6f87bc50e45dc947a08c2fd3ea4d47b0164f9d7b7479a9d85f1ef8cd34b634002b3134c1f6b72c404411b219c42016205735cb79260d92de805993a3241d3d87fca89f549c418ca6ef1a960caf913d017ddee5499ce323b913bb49acaa847b4743b9671e2857cf6fcae9e69259471522aea9ec86cc4c11b77f71ae9b2a107c5563522ce609f236d4b7fedb29d86d3f3e481119f5034821b6ad2d298ff75d5acf8a480433797cfbf0a7b90029cd92f42cdf2c24d3652df5433c162d15d96a4a6d0be0c1f577b14f91bc99f587fb1b3b3ef8b727f3def7caf0e48a7b3967ba2b600e82b98b418bd5f126a4bfa1ce92e74ef00ef63eac3dfedc9176b4dc83ef1815a510a2660dd61fc3180c369865edeff9bbd5fb7fe4eeb8a79eba72f7b473bd32a9469796b5fdb9138cb29142a9a4a2561ee42f4346f70fcea338a14441c7a2a2ae6dbb310396421a4f9bb53bfce58949abbc39523975f3acf8a804fe59c3c8b4c2e9f77b79cbc00ccea96efdc772e372981d6f0a79ab23d1d7e8741fb36a4007d33535546e4a909fb29cca3c0eae83a1ab3d535f9d4ebd3c57c8790f8613cfc40d31779824fcd4b47a66238320477d06021847b54ffb75709f202e39cda528e5c456fdc5bd13a2934a9db52a2b1e5537a1a2fffdd1cfbd4c8db10c62d0a6dd8f09075a91aa62ea8b983e6a3a55e524cc82b0550bc56e53b6df5ff29acc66ecbafcbd191ef958d95d4a74cdcb6e719005c49e674e8c856673ff2be8a88fea3a714402664039b48a83a09960148175a29fc568792868612e22d6859da124df1345e2d1769e35225d7eb858fdc403f762ff14acd99e44c843c8260403c0fc4327e38083a65cdcd3e7aafda417f35f174c9dd8b303252624d32934879591199e3d1c71d45f2eb417582a09ac325767e8919e7418893036987ba97adce694c112fd352ebbca96eb8be82f34eb9942203b3556003218126217b5a9f22df986273da0bb5d95897b55ea9ddf8e597cb3073ada11b8ee9941fd7438e7cb4e8ab9994caf37102e9cc0af7d1838b071959ba4a7766243c8ddaa59b580ba474b63ff87c884ccd37cfdf6d1b614cb21cbf671a243a1e659ff66ae169ad40be2fbfdb4c50fa7c81cca64dd4d5cd5785a7b32348441e88630ac01f139d1b56714ef6fa940d0c50b640dfe0eada27a8149f725d75cbe17c3822169c893dbe5e6d912271f90eda9be858a5cba08a9355b20b0d0efd6022b6ade30efb917a226640f200a1f1dc59ee8c7f68a197a79550d186fbef496693d1a972a17c4c4a8251aeb654178577fac1aa5cbfaccec629fc1a5eca73e2e6c0daf103ef8aca9af13fc01fa0386f268d2797aedeaf0a96cb9e3298ab442ff7ca2709b7c1827af8b43ef3bcb2c2f9cfdf7fc2608c89060147873551c7e3ab8b9dd05ad4fb8ab9f9a8a214e9ba4a411009f232f01f90a83ae0f101a438c3eba7c425edaeb59b178ec567320f1365e83a6942e8a273cf084960a4d40fd7ffd5854ff4c3feb0c2cff9d6ebca30c5d00df2a68c42b4d86c51c61aa99cad703e7d81aaba5b80f8ef1e355643fef8ea30921dd4e276846c7e9e3f35325fae2817699e92237e1ebeffdf0c943355bc62c1605975ac7d5169f9fb61a5fda2ef81fa65d3ea93c26b2b7d6eb70f48d0ce932b08c6be831ecd1c5e78bddb0e0582572d3931d2f82cf8a64e0bdaac69bb51833d5a16225c1348ac0955f9cea06f8981a46c670e46ae9889141a3027a96eab8398c9da856fce1c5a5836a3b80c6aadea56ccac64b6a30224173bb8247bd4b1c32c3562626cb566e416458a617b5ff11cb01f9e1214316062c57c7b6ca36a9c176ac50810c5bdb86250712e58c0c14abf4056629586b86ca4c58dbd732759e2e0a03ea8335042c347a9339249634ea6627c5ba3368149cc67193f61f6c242ded77e9140296083c2b95739733bd0223985bc0871661a0cc73593a37e3cd68ba4924d9a13baa4a43b8a90c8e048c2ad6b5b23cb6ced73b0e029f359124c79e744db60bb25104d49da50d03c565d455444e58cb4e6c40ae9d7c16e7fec589afcdc076091c052554f8255aabe178a81dca1e198b073b11e7fe0a23ca510f8da10b8caf22ae50fe3b96d89f6e225c0096c6c730830098c659e6f42816dbb4c7c2cedbaca6cce99ab6d49926f48c0f4b7a926c3c43d1d77d3214cd0e03ec9719cda83f7cb9bbae0b92187b0ca5628d676cb6ad5fa03cc0f0a13aa5b4087234bf5032972d39bc477030b9a1678c326f8e9e1b8237d56f906548b726104f02f08b89403d2a20244aa784466e6f5a105513c98aa8ac7091a34c9edffc62985d7c693fc98f298327696e0a064bffd84ecc2708e4b6bbf0e8e911a749398b55726c695b85a8e17cd37d79d8b8e7b153c44c53cdc46761ccdd11f37f939f7335f1faf8cf5b094625f840bce83e43eabb33f1923da2942960c4a14a6e8602a1ac2e8f0c937c34b474c26b0eba0542f29d80651a6f285618c4a51746d180faf5a1f35966ea3713f912ed14806a22b93cb517c748d5b2f05f22b6e0c2cdc38cb95032e401fdfa0920a799a3d1e26e000e5692be1f8fd6c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h92ad702fc2080b95c84a82410e5150ce10e727c95b7040d826f03a42bef17e7ee43f26d361975282c5d05be55434b7e9e8f4d3a01ae377feb933a74eddfdf4754689df3ee74604be713c464cc2178c2e92fd26edd9af54f5eda6e7d3cf62f0af0f5074c78da70e7d7d7c6a54dff4739dab6a384a121cbfeaa5184dea30ed7b518e4416c46653f29eb3729cafd5df9dc6d1caa9a457a8e558f9df7e1c3808c97531983bbb3b33c3e6e19963497a3bdbe3c3183a768c22207b9dacae680ea527ee4f666e1e90b2edfb850b5776cd6c94b98ebb4f1edfe80b97f57e6284fe10b8e6587cf351d94c8358a05ee0f6901b8842e8e0477a5999b26e5e3ca7bcdc35730e819914b1a0c20ca2c0cacc29182bc9bc94b9393a4e3c6a089eebd31420cad23dc2b3470ebc6c6b9d691e7f53b263333fb69e04e6ae0c6bd69b946284f8ed88913bcb8e0c86ad81db5138be190d895bb234cbdbfb55046f59c0408ecd19910cf29db0a2ebe81ea8fd97366f423a87b37ac016c56fad4bf4a94a85b97fc1189dea0508f77b6b1ec7607b33f6e8853c2168b6697e1281372ab65a4d3a24a7bda9eb6e55f805c06a1243e524f966df45a11a3af437e46aad5388089c3b7c1277929ac34eadc23955dee29d8e90a44c8024d53e5165562b8afefcb55ddcf0cb44b1fc58f26d1a420b8ab59fa10f84ef3a0d4bd40931a9d3c408d3452d176f7e563db9e31366fbe1e26bbb58efec13973d859bb5c4ad1ccab20499b52bf1aeb43785b22afe973b0dcc46dd10f898875cbca33ed1b69835aa18537509f8184c3f1d92423535fab38e41d4fb64d090eecf5b006a6dabf801ff3cf0093311f7f89a3c0659479d43e9fd6ba8f0ac9ca907a5a59f0d169952136d85ca3c409bae980d184fa4cedcd84f315791f9cfc0186443268725081373399b1ada5be16cb780490baaf681f4b503d9c0d0e8440997fc33c908d4eb5b1ec7d5cb8fa61dfefcc6d5f2db8c986b7a60d45510d9cbcde676b8da69e23ffe031ffc82dab24dbeacde8b0fea598f17872c9a728ab0a14fb60b1f2b28c1ad749ad5d03eafba880df302dd1f15f4e61ab736af2f91d03545db9162d5b93dfdffb18714a8cda8211331ce28799d5344eca147586c2bd03b19df10a0297580ac88bf0c5cca739fefbb4d2ca896e7429b71af82e90e91a1eb819f1ef94fa859daae8cf7a3bed7fcbd1114e33f15b7fc11ef87f0d862435d9b7769836d8221d78077b94a963c64e825c27c48c0e404af53c947c30d94093064cba5c4b42b672b27827589d0a9d4ddd66693ef052f55a4b462f19539a7a3cc4e20ef7541e206487b32a05a81c91b572dc40d51abba38bdef126b4dfd3e2abb85d1575e0e574d21b36c1e0b6a8059c2ec8020d2b5628783359a2ba9c1ef9aa12ff477acd50ac9fa9db8e972ca528b26be3ce25cdbc471659c4e8ff26ddb519f1daa30eeda7f674e4625e42b3e117a01f904b8d21a8ee894c556cca009b113c78122557648a1debf06608ec9f3837c84500ace4a1084a671679a50b17342e78d95b9bbe85e75ab75f33be4ca19ad8939eb7cf4fc1fa1317a524941405da6e40e7a9e892f0c740b94839771a87bf88a71505d3782071f79be439151edb12785124ddcfeae472790be6a52b4d4bbb27fc58578e26e4b67f5795403c491c71592fda784d25399d2f28def39f7764bf0e953fac89b5fcb82c539964512a8bb24b10eed91a862d7c71de4bb1363753dae59a3467fb7519bbec8d5cfab2b4cd4c99584fdebc4dd77dbf473b71999fe2e40f1aa9ab9446f84702d2c7dc4fa1db7b4cdbb95f3f81c25ea3e4e5d0ddab36b4c2b19c282bd92466e320d41d8ee66d0ffdebb59a2008a00630ab56f2c65560b5d16333879b2909412c196f93877f750c64290c32965c809cca24c35bc761a3246b3a1e9cdc117e442673280767d404eedfc53e5fc37c6f07fef2434395a6892fc2bcec0cfbcfe13c8dd552efe1bc2105d4329adfca2a26a86749b046045c5130ac4a58ba3606a9021d7cdca544616794e45284ce85fbeb55e6b8dcbf4027aff7009a83db69ba792549f8a79d092f2b7122b13ef8af33162cf796a3ad3354f3a096f9869e3e6cb18c09a4ccce81600506704e5b6a2b59a5c5bf3817599e4637f142ef4c67af5183c27fd519e60e86cf1dc06902c5bc4837f0d1723692987d0b292262fbf484f1772be901f6566daa36dee7dc4418d67c24782da223ff7bbec55ec6db39951dde331964493929b461c44a1275862973476942e935e90286265b6850ccb65e432c6c4ec81667998ef6694a0deac9076767e880d68a95e3c046a646f93dbb818cd4f60485e71c5556970059cefe2ed5d6733f643d3538fd31d6e4862b4b6ee4a9fd82e876b15867c9cc4da4df5e903ec32a814c5d32598f50fd7f04ee637b366887e64d72d65139353eabc8502babbbe8573344215472e17cca2cbbc789628faf1c2c741d3fbaf422ef298717736aadd9ea1a5e9d75a869fcff38f8f83569c43127cc7354a66106f120c16f445ca236b1a2cbb18801334ee950ac15a624736cecb1dcbc8a4985f8dd8ecb29f0d924574076841f2c2fd83b39c5c8c53ea1cf17dae5404f705d33a8e8a85188080f0127929a25b0b0a12db42eddcee489d2ec94abd3bfef989331c60a557c691e75cca87e3cf79700dbb61bb9ed54933bf8c6b25aecd790ce56e16f1b748a48cb130d9a4beceb0e9e06c32b2e961874a0232e91e4576b9b53cc5e2e41a356c4a3f234b8fa8a04a6a7b1590d0fd70025028bd5612674f8385748e9791017fcb22d88e7b460b13e152927864a98b18323bc74e77b5cb848b44fe683ee61dfe67bff5cc1071da8fb6715aa7b32a4a99ef287af86f9211eb212756b0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h5dbedce39f2352229327808b5dfcc404649a90e0f769c830591f766d22e29c5ec45335aa1c25a3209a33055e5e14febcb740ca27fe04b7c025ff5b22f72d6a7f7c4e1aa45ffe7578e6a69c446d9e769d5222a115bdb30b7281a6ffb325394875897d20c3b73e4cc13b81721364dbc3bf815c26fc374cca35eefb810d1a439d861416084b3f388a5e1dca4221f71ba0dd9a6ab20c8d4eddc8af66de86c6a57a3b8ad74547eb96a18d148e05693af2c4bb73575f0eca538199cbfcfa7fb94d71c2380beaab6ac0d87880e3d744a9483d32a71af058843c5d85cd099ea22fa806d9fa2f91b4d98267b4c50370e7e306c5418485e8ad4c874db3f344c0387b34488a0845e2b1be2ad5a58d277b1545ee22ffd2f58824fa8d5ac7cdad17d8021212991b76ad883889561c0d9a878d412cd173aa75ecf701c8799946d98e282cc48cabe45ca54b2478ff0f850a6ecc62b9f8f4a3e5a45afa5c6cb4307b2e5868a3b35d81a20f345eb7e40ecde1ef26d28776edd591f25eabe9da161d82b727a699b02841b9b930f737521bb2b696576bb05f5abbe9809aad2cbb1f8294a17a77df935646a926df79846dfcc7cbb6e928b10b6a2a9cec45578db0fa7b40f54cd99978275a3d94cc4131c4a745ecc4a2e0ff580a32488263206f077d9343081cde44212fd59d220ea3fd0d211869915643119c905dc9211320e6cfb6b0e722b3cd7745415d82129f8846e581a6c861d1701ce590317a505a668dc919600b2582e2c7082631e93f639e51936f5f87269647646a1e3acdd702cd8010692e58f0d789c6f5d2c8e3c7895a81766dc63784804f2f08dec3f0647d772b2d7c7c3791d308643cb76e3cbda5381812e2cae2c9a9d7eb3e74b5f76ed88e5ad4d564b1b91445956d52c5ea2206c378232003b58d947ffce451e97a6324acf6de12df40fb4ca4716ec60edb0edc7cc1a76235439263512d8ec0cbdd70d469848d65a8ef771469169bcf471886e48730ae4f3bc4683ea22b77dd1f4ce01b5870ea297771c275ce4199ab38a8013320d44935f810d4e845e637f1c86fc43bdab5083890a66b10be19c935e70d9cd75037fb4fb81853b3cdb2d8e32c4bcc7d353b2363d10b391afa5c84b0de690e3fb8eea63c96b71b34bd06f469340defaf47881793a201fd9a47bd066c7313f53a819e3567f9259aae218700c2fa8da686ca2e7e1c3c04f37a896c133ad9634b7e72273d32a47265cf302376e3080dac08af55f96b523613907d3f0f24955382552c164d06fe6f5bda7aaebd4a81e1bf51bea1746b2894e98cdf9cb402e7048a912dc23bf228d2e15ddf3357284bbe9e109f997027bae6275b4404ae89d538a70dda9bee6ec28571845fd1985104c3aee881e807485d00d6d2b5e76df0b308cdf6017da6f3b4628f305863c3f60e7d6e47f0faba46565c84490d2647fe28b166cb7b19331050ae3a4d41a41cbe2a2ad5d1db822085915b3a387cc36e82475e1b9292cc8dd05378492f13f706d8096269922319a00b679f70b5243103c7dda846556485373b8d35347b80913652e526e570ee14104caae74f465552694923a193dd4c12be73922587fd67d7a5e7e49099aa450b929314eaaff64743f3ea7bbd1ea71e754d3ca8d14150bf2cfef73bc26aee8dc4c9900bf5d29fd895b4f75e45251fa077e797ac00fa1dfbb8536a7cc887c1989168fb12be9a81e57c2419e487b78f7a7bb9c4cecb61fb2be5cb2c951b4ece61913cb27ed0062322475f52632efa2cbb8d229025bde4db2bd1d9ed73ba55ab81256c601bd30a9d58c799295b9f284e0ca7f0f9afda5c27081bf5f0599766c0c5691a8febed523cc1ebe42c3bf48065d2fb280698e6b3d15fd521daa930a98d9763f68fa20162244cf007f1803440c6fd1bb8f81151c62f99d707e32c36e02dc80c22022c225b573f6db798eff8b9c850003eb83445f61415d489ee2b939c8d94c3dd7a1bd6c07a42519082ec0c2eddd0a9406bc817658222f7d31b2dd0244496f945d90da1584c005d3acf8f9eac4eba813e486ddf52d138df4c57062ef4dd92ab177a18da495593ae227bef834ab5ce247f8f39ae3cd80534139cc44617164c9aea1ba5708f7dcf03c8ca9f373e9ac8f2fbfab95deb7b81fac1dd2fb84dd15ed6cf1ea653e20f0abb361453c2d571e2207e11a6cdecb6cfc288e1881674d38db7ff7f5c6d3112f2f58b047841d80289f9d6a9fe563e2f8190b79695faf7ac620b59d8b4806291b895928b2a9499a5a93a7bce6f340489388c98c2d5393ab1159b76241d4ef8698cb4e64968818e2797fabd77588f2985e6bfce67faefe46b32854ac5ce48888635e3ea01775f8037a13cad2aa3b2fa4881f75b969062e4f6c92eb822d0fc14dab8e261543ed8459893ab166316b471a7bf8ff4a1905002c7269192ee5d3731be75234bf7c3f6830eb4a12e2e9ee341a6fc7777c312a81bb25b614cc02d2866429dc609e49ac1e9f4b88c48a018ba5f2ae75b9ba0fce56ac94ba82531fc4044f0c2b3781fadcf75db5008fc58b3a88ff33fa38267d244f1121a52df00fde26ac0d42d402360323e10824d83c03c199f7b75d90a945a31019f7bf17b3237d037adfa6eb978074ad34edaa3cd798dfb32473edc4ad2e42cc4d00d6777028f3d973cbf3291ba93eaed1cfa921d519e14ebb60ca6b695af7c25d134a740c977954c3fc1b58fbeb6b9bc3b82507d805a0481459625e6c2b1d3eca4d78aa90e00c81a4eeea6411220c62fb1aadcf5e4d89bb3996c71e3c0c08bca7f74d7cb907179ab05af4ad5c86b7e90d0e478cd8e0a30a9d6ac5419e9ea2af9bcc59de9e23e141d40029c7e140da094d1282dc5b9e26e944a90ab4b74a3dbefd9185ab81f75424a946b6e49c5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he4318acbafe1f2991f7ebbe0427abd9f8d186a59afc3cef549da61f86892cbc690887fe6a7f80f3bc08bb6dd347eaf2efe274034cad30ccd7318f0e74d901cc68a99727c1e54e464654442cdaffb3790feb4f54dac91e7e8a69434f6ae46851651243a826d1b77fe60906e4539a828d4a1f0c0cc669cd3a25ded1f0ad913b76e6d246c00580ce68df6923b0cce546a8aa0635c2a4de3874fd6e479890a328f001551dba1c3478c73be3460777f78b38d26ccd14d141b2b37b327f60a29c61d3a3ea5e482896f01ec8e9c3bb979e4773611b535355578222286d98295ffc277b41f50738a136600ae665343735fa9f5383aa5a75bbfc6fdaa7728b76fa88bf189061e43f01ec8ac1defd6b962fa5853e63c25be2c302b4918b6440394fb1cfbf1091d6ed3eb8c2cd62b6531e8b7483fd47e614863f84f5d08d9541634fedef2057c558ca8a9a877d5aec1c84ed62e518fb091ac149ef1daed528f2222ff64b2825acb72fcf226c13bc7ee361ccc267e871d45de3b24fa3a06ff9905f67d67a3f0c1e10a3472d5d90a011af5f745b9d1a01c1269e017bd4e0df77428b1d70c8bfd6279bcfc9773d14f1a27138dd308aa58c16857da6dbe7db3d04c3606fa801d4a1d182396643f275fbc05279766628992405e3a3d4d14361f7167f59960e72718c3ea2cf57f870f404f057fe2451877622ea66e797e500fb98d97fbd52632fbb6d63bcc67ecdbe07e220c1a6e2bce88dcb7e572c4b37a13c366e6f8b6177bd07b5cb38292e8dc6de00086396dfb2a92b2f4cd75a4cdc6c1dc6c89651da539050fd57006d86bbd40fa5d3a69ed7b9e6030b914a6237d701ed8df0d28d7971d42f66a19c5c4f25970c3847782497433e0641ed79ec820e64a583c4550fff4ab1767aa162cf973d57da75561bf0e5f280241173a959d2458b796c2a4e10f8180dd6e2a2220f00734528dbc26ce4cca3f382be772a1ba60e3c6f2716ff35631a45e7da0ed76ac51697208ec5ddc445db1aaa6580e0af9d7c713d301b8db1b3bd272864e599eb76f857ad1365ed639b0a9e574310177b1b23137e6bb489b2b264ac80743197cff4521fe5a3fe4cc4f8f4b4ff3d08c612e1519ec521c2cda3288333c8e91d0276caf81c896dc4b5e9fdec33705c8fa867a33cf9cc397e5cf2846377ee974aa8d4375cd8aebfb50e90214fc7f0c6492f58e2ed1b8895102e088a4637ec619072549641281e0d3bcf21868118e45c568a58f6cf81bf425fa706dbc79a0be086ac27cd0aa8ab2302a9216e37a36fb01d53a9270b3ed0978e283eb2ceae2add1c13bae1cefa393a8bc4842396e3fa6faff10c73aa61f4bb98859cf362afbd1515eaa97cb7631e74aa5b91bee01bb7587bee22788af3f4a8999dbdbdd1028cd96ed88ef65621b06007102bf0a67a7f96c952f339f66a4224b99190f2ca69611f858028f37f7beb740d773b2f83337aff7754fd4f83dec83caa26a9b450799e571c339a459d2b0d3104b8b134938746f2c502684932d8d9e6a73bb7c433819e2d7a7d88880ec95aa551bd5abb075555e40776d7a59c2272d19001f658e0d23ec2e9bb4ea2255099d3574c962d6625259523da55ecff37382935eef461f11a500e9f78563ce8cc0d345d27f795e3158de17e6abc8121208411f8afd74bc6b6597049563156663d42f85fba9213237051e95a10786f78cbee7521485ee75b37d0bcfc9d37fe08234bf8e5f2b0e828af26c6f1c709eb66501cbb2564dea022950d1b013b86f8c441edb07384774534ba7fc129b27c3c5135d5097092bb36811a8536b4f9d413d314a06781fd2b7d59aa2a03ea48dbf7b6baf5bf4e022fa24e33eb265a40a15692879b381fbb30c80d7df0f3a710635863f09f18351686b7180d5b30c399a0ac6bde179a1fcc2719468fdc480ea021d0594ce45cbef927f4987a34c3413e7f86bd74ec2be2c0c6d7c059cd5d1a6483c89ce2e3fb439c570bb079d02c9b633e9009a56fc65115fb4443b546004355c5e07dbff17583562092e922985c5f423bb850d5f53e2d3d920a8bd958b3191c6a7949c229793065ad81f45e97b08fc5f7bb47b55c5d56c3a50d5603b1375f9ec75d7fb1cb1a2016fa92e18cdb0d3060715151aa6e831d8f74ff5587e62a2706580331662b4a0857d4d12f3fe3e94647190779de25b6af84053256fed0040d3eed57d649e0d523726847a03b792a1d703d83923ebce48d9487565e4bc173ad3120b285f8296b78b64777069cd8dcc16523079b2848e1a42eb2d8c4ff6816b88935238636154b69497fabaf91231f261110ddab4133030491612f3e7da0d90f1634200f2bb28edb7c0542614bbb486b84c3779d089e476313567485c72a5f10c3b1eeb67e496605ebff667cade6fb4069a88b391606156fbe9f08cec0f9cf92d7bb1b4c2767dd61e3f60bfb333e0b482baf23c1a4fb4ead2c131877fb7c801964bd8b1bd9610e928c5245b1e8e28638f2ce88efe3ad0cafcb988cbc72bc0cedc629521b8e65e372c55cb6a3c4ee9483c0f72586b645f16c2fdaf406ab2f3a252920a2f1c0063a1bd41586f9ab129763c5cae7eb4882bba8b7463ff4db41b62b7c5be2c6f167e4553a204b6dcad43ce566ef1d2572666712b9dcd36aeabcff8108a3f34a1fae6b8bc55df90e4af106343a33bea123e5ec09d867e1ee1751c9858542edd82ae5d699b1319ed75900abe1ebdda1e595b9f0b5d3f7ba36ae265d1a97406f2deff13507091f235e9924b7be4437244e15d4830b7af65ea72edfe14baf8a518708a3895bd800f0f7c8e805bee7e7d5574742492fdac641379b8de5c7f85b8fe2338c22f05297478e6d9ca0b58451e5ece0e25682fe4d9344a766a0f591644e4d4403987b7cc7c4297a056;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hacaf2a755d0fdd9c2035f3858a183516f4fa6f3ff41b9762926156991d8fec2d8d82e1a83d59f9538ba49f732b70d127cd600405bba5966a4db7526b49826a00fb40d508dde2b8bb5b29d5fa06181657b34179a1868c93d9c7fe7f2d0db6acadfaab32eaea5c230fef831574f72e83c20985ae503f96424c22e3f26c95f72d291fc0736b43f920e164048f07088e55fd879626b6de56a3eb7db41564eeba0171ced337cdceb01829b0927528730e30b79d50efa08f96a3d67b1d119d893597363abb2a4a4bd8c1cf3a07e6afa531fa985e86846ea2c095d286cfee39a452ae2a0e674f01e19579404e4ed28947355835ac69e2d0ea371e23d8d6b6c5fc2df42b674bcaa9b1a348725b78e3fe402d11f7cc10740e023440f8d0983b6d628cfa4ce4574018e4017a98896f981adbfdb1cb75f9371bb28582874c739b92208c657ab25a1c67ec5e8f7bae8e03a1d859dd3ac3635b95bf18cc47239f43118c5fb4e0bfc8956021804077127d0ae322fcd8f9c2e7bc1eaababdaf27da94cd8abdadecf6799111b709668b510ad2385648d97cdb0b74f4bee357ac0f2071b00d1900ea83b631cfb56dd4e52427fa576b9e31e65e91e4f9fb20f0b64185c0fe21b87a2d3a683c84fa716ba016b37d6f4ef2b12810f6f3df56736d3b84b1d6a3b04b5ce2dce50041b6eade7d3aa09288854c1339323358a701c14af104d29a02e9a959c59b8e51978a7e173d774828ffeb166d91f50ecd017c18b8f5e55f176145c7354fbe61cbf0a78ca96a56decbfd5411a70a191126fdbcdf6a4f9773ab71065ce0f40831acad89efe1b0ce04cc49388a8f36d9cde659b1e309b06cc1b96b514dbe33b90ba79b337a5a3880659d22454e4f89a8c6d215ace79a21026e81f27c3010884ea2bc46cc446e0f1eebe974a4f5534426bed72f9067b42f565f7347e690602eb72a92c61355a19789423be96375c789a79925ef8ec9fa0cceffeba4ecf4beec68d7e1751dfbac5151c7274b242fbc95dc63eaa9840db1549bd0343fe2da0421f47d3a125c2303ca3ea81f1ddfa4bcceaceceea0514008e4944b8c11fe3bb674cfc90c83751e2a593e24aab03052cef5174d79c004a9a4ac5ebc9465643153769b79253ae305725a0bf3d17fb9b168ed0ff0b3cb09b6377f19661949979f2921b337428bd1a48fb2e8da3d93e989a4a70d5afb3eef967f891e819a48112ef1a05a8a50171570c03ccaa115c5432323cf39156659b543381b14ae7c3629825f7820b536f3bb3a770c6683695a119421716da86d89001208ad441e58f6788fede92e553c3d6b8c7577d9499b31fb2cadaa8b2ff657001d4713451b4aadf0a095a4c530b3dd47dfc35067b340da3b0d2543950fdf1dec3189c1d8c79c44bc666a5e4392ca49859c7822d40b35456131054b2def643888987ea402aa15c190d210ea3a3adc5288f27963111aa94d35cbeb369677b3e2e485d7e52b5fd5435c6ef2905bf97d6215c28783343b5613f9cd25c944a5303d467322f83db2653b16599c817baaed24715e77ba52ceb8b8e76d1e01371e7a982389fef28110c2f0e3516bb0b83cd9683d396964c5fb1c49b0ebb4b821b1a307a146353ebbb71eb53d4412301f938f183284d9e22809cb8e0ac092443c6c470b5d7148f7165276881f5ac7b59abec8bfa16915ec2830a63b5da47e9e3a3e6fae21eec9a3552b6ee66782e29bec31f14c8d5a9f292f4966f77465fe1db17968f19504971fbf20a2a4eddc5c618ba08a708147f5288573d26804f8b9703263eb4e9706bb7845496d2f96795cbffbe1f1aa2d9908363c61910a2f954642581666b75a7875d98ab2418e1aee5ae60644bd1573a330456144af2312208a875ab1317dc02c12d144044f72bc12a2e2bb8fcfb493ab7e161cb4458b39c4b16ffbc01155a4e8fd033c39d6d634d3659188c2a18c043872324a2c26e0cd5a1e07dd48f59e82a89bac83abe8d40cf38a28c344eaa7aa2b3a803395ca72a8732ffeb8188100a5e2a67c04fece3f680a531913157e0c769ff73c2b0ad80cec2dbbb485b13b28a98f778383f25314a1de5416b0d336b5e8742b3b9fb40efa6f48bd8e068d15bd7c0efac7af0ef6bb3ac0fbd080871cb19d731c4353c5a39e8b9cabe7476aaa6e5a394c5f5df1c67c29ce80deeae445b841ef36931599ab081d03005e374cc812879a41d8f5108cfc41a237de50889d3c2c387fe4ffe40b9d5ab1cc72a29de15b443b535878c0d4a9fd4e7c85abd745a254ed4188fc47d23651eeceb3bcfdb13b9cd38e01b655bdb388963c9b6adcac80f602815a0ce7fdc5347f52d914adb5ef25f6a4d2d942166c0c79e223802229fcb37df862e6dcb0cfb424f744e7995242f846bf672c631f3f55cce96c72ba3486d83cf4296945d282669f573c87c222cfe09dcc18e676c430b19746c6256579154e2d312094164f80b3adf9d5df4eb5aa3ca9afc60e416f7033db3ec687158a8346bec8ccbe8c97817117f0d82cf9351b527e674c14835b9b3f9327889ede81e1cbbcc7e613c50d1f31629b195233a82e3b2326f983100d72f62d3fef6ef69fb258b2670e76e814a9c433f7e6dd613c5387cf44eecd0a27f81fd76e533f952952fd476fd02bccb459b7c493962d9c50e18c4eceae8a3bc3aad534852273fd5505269379b86811b87334916c8b62daadea7d8027c4473e6289e60bc30ba6d5c3e5a9af1fe8d33fba80ee3ff21f668d48607d77cdf4bd0861abb1040832acf827563cc348e13bdfdb52c76644d8d0b3d844569af718300efaa78ef0c63d245d83a0ca953b7cdb5ca4b857f915869d7a443b30535f5231acb96f5859557f31d23c89f0eb39bedc59a491212093229541063ababbdf0fba24f001b208cf41;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf5e96fa9f22c5457b50774c66e1811c634870bbe2755c62be6f0603f95188d69abd00f8de5a749fbcd85f8e25cb986e7a02edff5659ca8a8fb67e613926c5c75cf14d6ee56a57b6c14fa6f4bc13de97801f89faa3132da98b1bb5e921767dfe65ed54b51edafe979ec03b996b962cda6b88b2474f72150ea6dd661cc13bb641ed9215ce27caae093e2a12db488ed145992b2aaf0b5d38cf7d97df93302a2dbb8992ac7a0176b6573fa532dc8d03511e9630d3dca2cec701c6495c79fc890321b5040c58b63c9aedcd5db2712e35b01c85e52d66f7e60a08bc83a848190e57e37ca0f3744e0e8a80686d0914914b3cae4c5c00f98d3c614df988cc39cf4f52c082b88ced2dbdfcd0dc0b4feee4b46770598a0bcea692dd90da16b73e612976d812865149b5c565aaf1de696f554eead606be38fb7d93b117af7bc44a41fe7dd61bef0ce994e75fd8e60eadd2d740e939e98b41c525145356fd3474bde40571373ed60fa4edcce51babc5ca975e597556518f348fdf64c3f0379ad54b6c4bd141a591d5024d4a76988f0c6d21b1cc3a2519531ad2d8d5f2a090ce70b282d74a9f5a5710bea7ae9b20dab4e97f5d7549dd393527032f9f08d8cbfeec017dfe2cdb03471263d3f9486dd837e36ee8edbc59e7ba0b621d576d896c586c31ae7d74aa54c90ea6a8a734b40507922565edfa60afd80f78cbea7cda4b63f3e6e7ba421f223581596f0f0a42d27161d981c5b07822720459cd777c3ce286e0477a8e7c54efe1a119df563df07ca78178ff0c88bc695eec0ef6b0bb5a0d7fbe4b7d311b060c235ae31cc6fa1e5f7c1a3e8b3dfe362174b4fdd1c9fd44d547bc8173ed85b47ed4fd130194b0afeadcafb764ab70dafc5843b70df1442b01ee0f915224d97c5930e59d9ba33500121f59f8ae4960c4371006b1846121e35fd67568af4bae10c17fea15092518cba763d788a7edb8a41ee09f03c6f9315ebc30c1e036a1c4a93cb754e7598db33b9cfc21ce8244012c90dbbe5694e9d693f86686bbf8ee755bffc85808568dd0e9b7d5f04069d510b6a3d2266e60e12fcee11b080f188cfa9cc0c9139a5a4d1fe8eed60a288db9af38f16e4d2db610174a7d85f80aec81e0892f494604e4e74a42e834567c79f00f40bac15040c7976e870dd015d0e343ec36513d2e9a66cb8346215a5e23d7f39dfb91c56f9aa7b477e6b375ab884d631aa0dc6d10b87adef47ad79e2e08a471a43d705ab0ab2921b17d7165790ac867074dd8c1b3d9c224858630abbd7c01176bb010c2fb77f09e192394eaa2b3dc6bb4ed98eb9981a9f4b7d2067d2044886d9bec8692eeea1ef64e2af09826ec302c364178bed47c88d21ac1e83befd01ba9acb96cf08a51028a806e56bfab198c14ddc517d2cb7355ac40cec9b2ff3cdb2b5ead2ed16a3814a9caf4c38a4add35e1e62741248b137787af8bb99df6d72941b81badaecc173832c3f8e8c55711b96baa416cd3b97474974e8ed7beb270eb83e2a086fefb662e0c76e88d76902cd26de4baaab3a9f4d3c4da4bb98d86fcc69cff31c28eadad6c0590c05e42e6b1ab973fc09d18bdf445be7ef3675ac57b7708c9e8c31c2d0094f7168eed6eead1b63cf66874e438914895261af39414b73f186e5d5f8360616566576fac3df3c3df410a7923f70a69cb8ccd717657358da107ad67062dc4e8655c966389a90f15764da89e294922e43ab01a0cf8aef0e30f1b8bc430bb65483cc87c087e44ce981550dc4a9296b871d6c382b8182c545dd82f10586081f087ad9d948e6e9f422b9914d16da2aa4ab396028270cada25054252804a18193cb2603199d06ffc046f5bf6238621a0704b48cf04f1940268997d22ba0c810ae8aa9c0bea313894365afeb8451b88c2fbdf182e4ab12be932f8905a973855ec9f006825b9c48beac95e2f19ac51bf6b187ed3122dd82cfeb99f77ebe4b10ac631ee86f63de448336c3ba9ac99566929622114fba1a080eb7da3c11b0395034b3a0fb578a44b712fa31f059b16e6a34c30ee38f81106a09fe252e38511d3c4699a09ad5bda1214e0df9954fa592d73cc84f131959c537163f8fead2270d0905fbbc6f9bc631ce61f65ace713460077a54fa9405bd2a99089990b534f0b8dcf73bd62e4286c522360d9a71ad1ee99878135f65d7bf1ec80b6a88779e185a773cff0db0437e5a06ad8a72b23902da9415d8edaa6ebae95bbb4a0df821e425c5717f918ae3dd8ac8fd1f11258dbcc6c308a335afb1a6afdc39fbfc54d22ac40ec0f4860b1c9cd141f8f5eacc4021a28041e01f9adc405d3d142d9418a4ae3f482f9847bb1221b9985a051cad204d1a663e204c90cbb83bea64b4863e08afec7ce1feeeb878d5a78cf3574f0a52dcc94e48951b096b05d2a606f97784bfb8b87aaf503f251c8b3078f10779767a8e5079ef698050b6fdc19a12a45c968fe6989c76193353072b55b705f914a1970810f4346957fa6e226f4a9d4cf8b1f9587d741180a6910a445668def72ff37cf2c6941b785348492340d90c85a6c4705f1174c3925f661c0e824fd4041a233f8b660c286480579869401f11eb3d51baa30df0de91d044462620eb39d8e596f0ff3f6902c86e65f82f02ce946b88f7e2586173fcf731e1e863974dea475724519f643e1261f226e20a50ae6617f30519e989849e077d91ef0896a93abbec15cbcd2799eacf4ac70be0e869247baa1d6211ecd5948010bc4214d680afff1b19bf69a959df3abbec4d56ced4b1ab7b799d956499cab33fe5271e8a7b30cf2532b2742373b9bca91fa7d4fb713e6321e41965ce132d29ecf47937dd3e0d80417bdcd2fc266d1de15b3e07ba792563e6922a8800117d544d8807109f5e5b6743ca25ae0369;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb2266c34f3ca757584eeb3de543f35991864dca36b1c00bab9ffeeefcd6c07cccc60021c9b2ec5618007eda128d056241ff0a4062fb24545cfae7c2de421da85aa884e1a2a5522415989a65b9107abd463b95ce512ee6820deaded4232f8ca3c33e28cca502746f7b41ce7d88eb854f6394716c4eb7035a703dda59cec81d35e08ff86c2e3d08545682a62cb8f6f4ff6b90b02cc943d58b11b6c9712ece7902efc97255251a80830b3f26c698e7c957df011ba43e7919dd36e34612a1842cb579d6d266fabcac2d3cd68a65303a4da74604ec2bf729430ff188dd7a87f4a7ce5115bab5b8e681f03305c62ae2ac492eb53c280a6aa4cfeda5fd1d7fe707761c98fe617102dacb56f405a46cfd9f44765434ba1dafbfbe9b3f4f22ce35bc125e0fa89c5842dd3cbf1118fe63f40fd8f4a0d398d721d6bf20630d7ac6c3913c2a69cb8690aa38a602c891decad19603305edc6afd38005a3f1a69d47330de2951f6be4b0ccb851720a179f9ab654f0cf022a50023dc6ac94a0c08ba253f9d1fabfba87baa0661b8a6871e422c434e468114c2cb8e541ef26cb1f9d9509ad3d6c65bc3dc07ea68b7b834d3628fea169d47c9a8ee89a3164c790fb80c762954c845ab09ba71d2fbe18803af0351f9788935d6b125de19f3f1ed490e5765178a85939809b4f8f034d2fc912001169767784e6b6f65358c94c7afc03fe495d29c30dd2aaa381c37f5d42b7fb515a470af998c99a66a499caf858430b9f39540a548cd2e15323504951eedf51f91fa4b34f292701bad9d4f02d2ed9815d9ff04a8822a3335dd7d5789858464b3e18dd44d400feee6efe9d8bb9df1025e8d5010195cdd32e704a37529d154acd1bcf287dee94b2fe8362cfcb54f2aa94d7f39e750bb40e01aeab1baedf9e97622689359e13beb55f5dce495bbe84f13cd433f68eba67fd8c037aecba51e66d2c01fc2c116d5d4d970621cfd053053b0279e04716806786c0ccf424bb3304e614095318ebad26ca489c593e5fad842c2b6c26c5bbbac5774cc97757f9c878e12d966fcf43f6d54e45eda7fe0c03c08031bece288d4c8528953474bd698c73541eb2dfbd4f591633c255ec902b46ae653b101b6322ed1a6b324d90da9484bcec54e1497bde33abd0807591c5ccfc5f9a9fd0b21d17f4d8f5d4e7700e396df1a12d34293f3fe88e92d5d6293b57dfeafc459af0dfa95bda8780749f0c1579c01fa35004a228f17a26c2e4efcdcd4badc317863c896803b99f46b64ead69459b9b561dd1fcc74cd150b82f4d8d6d51175b97bd369ef80895052308968491bc20a0b8aa77317be68c7f8577222008900c1a2fa0b5dd250d28586759942369c786192bf39a136929c7f79a081e7fbe6dbb983b633d6cd57d01f38a2a40b2e9c76f2ff64ba59efdacba7f385941d70f36fcbe913d0b9b84802c500d23d19b6dbfa7bf4d72faf539b87012c75f9cde13cafdfbbc3f7f903338bf475eb26dbe5f93832093a9bdf74ac779506e32dba2ae4063230ce4317f10414650c29a2b5a87dd079bdd31db96b41576984599bfc84ba6f8c2b9dadad246a16c029bd0b239ccae4ff004181dffe06e476ad22b7e0ab4ad5eb0e3302d8af7c02b8e4af9dc4e3fd83271ff3113af79aba729a8f9a8a8fb09a4eca719abcdcb70789203d36ea436465868f7fad4934c14ec3b581ca7727bcf1f694db0d1e4bd8a096caefd0bd4e2ffbb7180db5d68c4f49dbe54d9ed1892ce741753686f1db304d7648ddfe274c2cbd2fef1331dfbfa2d38c6dce971133e48a56b66502b52ee35fd0f72e2ad0584b42c3042a61223be36bee8cf1076f1e583bb96346bfeb7b447a5c6d0555662bbc2cd73d814a921458752876d5b983c11072bfaca88bb1018ec47c763883b12e07d702551ca2bd1995242871f107d1baf06001c29db72f89917d7e9aff146ab4ecbf71871b57a7fa55d022eb90a52b6172046dff1c7f598ea6abb2ee4424c4abeaeb5df5fd25253e111728af95afef74526fb71e6a39b7e31830a0603de5273417eb6d82a226355087da68ea2e12927b11786d32c02c41d5c487af3ef835a1dd10d425977ee2e181b8904d56497d01151e1c740c626a2ee3df3d2bcfc395fb63789652eae46b68c12825b53c7313c339cc3372085365af0728cc7c62c674f47038340290ec75e2b1eaa201abdcdab35a97d302564537b20eb69d4c670c71dc07b6ad0f494d56c6b0728d197f5de5bb29999f9d7edb8dbb74b6e85783205b75727a23e7d143279a49f047f2a541ed1ecd0b69e4891479a960e0083d7a4190273f0818e18b4325d878c32c9b57d0ba5c8e979c34499f6cc2ce49750c3f0bdf7c728b83d45ab99d63654f68eafc6830915fe5b63db9edd65b4b79598ccaa3688f676f73cc957266b3a001571025c0c0e09e40191f27446b96c5a64fb0c380bfbc693e4d12ff36f85e321af9838b7d6ba0c71c37805b5302a6a921c0aa843c95e3511788e7e678774a59e37c39826f6f83384b0cd47b9e1af9431baad828743ecc61e90c544d21ea5a24c2ddfd3452dceec0f6a50803e96ceee9f7caf01b42f8cc94f852607149a5b3afde87cb657473453669101e45a4d088a757c9ac5cf5f2896e0eeec9f07014ed7ccfc73ceca9c76a3a4cefb288df5611b1ce7dbb02255b940e4663561a84a3575cf95f1069a615f43f1a594eec24c98b81dadd82b90c5c4371855df04a8b0940b3b71cbbd3f8f4a80c22ab0af13363348ca283b85c4c66da32392fb95fc02642319ded8a44c669f9c37b31630200cbbcfc508aae9a178f2e555cc9a1b6ec63a7939a3995eaea512ded5ae23e9b74cc4a103ebe4b1fb61b17dcf072fb29e6d853ea26d6086e677b6c546cf0652816b2f25ea230498;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h717a12398835a0906761c8132a4ea7ef442e4247c13629744b305187cd47f1dc52e7c03ab3bc82950be159b9c406d06f02e3d4981ec993e4fb9a972a390df1bd506887df6871ae6fe91bafa80d2b780d4718ec9250cdef626ccf7476fec28bef4fc7455d31ed06626641218a5cc0b9115c4d5c049ae7a6a3e5921d05ec4ad717c12a43aec5e30b5cd3965b1f40731a39fb2bad8047b7daf9eacf9ff984596707796af05edbf452206d8de74a22527c4d85f4f2cf34483129522d1dac93d0c0f90dc83a4d87673ad00fe67a45eb93eb7fa7725750c8a320f058605e4839fb7bd6853e062e1416769f4877fea64d956dccfbebe2f19cf19b1639dedae64c99ab42ed77e27ae5dc5c09008b6a2477b12b328962a703da3aa3bce7a8ee0f87ced3cd02fbc31d193a7e2b25ce83d5ed07c09962b7acf43f3cfb450cf599e6afb97c8a6dc76ba18b579519deb9c49ff1aa2fcc3e960634d2856af1a430c5e8a01fdfb32f85825ca65dc6a53dedbaef2f2e9e29f2339281b951f3d3864fd52c1557d62b0fd991737bd223e46e55c55a408a7b4fa1aa01f9368e3a1bf09b8503614776d775ec86ceb5d4bfaf4f01cf9d443bf83ff1792aa993263775f3203542133bae39d9516fb6768a8c5fb0c3551f7fb51cc936bbb93ab01249d5bd32f0298feb5cf9a35e44feaeb31b497da832e9b0af1cd81ea9f5a7edf5fa87938b4e51871406bc4e2d77d8078d28e04bf40f4659717759ff7ae4b88a7db58faa09bae89c71e6fc5da2acc4539a17b8b002a8f475f9db856029082902d44f7f2059495633fabde6a3f2614ee6fac2db03fdd31573d5aaa3b41d241d7f107587535c1b97d9201c003b4d8d8abdce45323f05b5ed3f0c9d4ae96e96b3cb5218f7a55c276ca90d04ef98fca8df6e1abdbcefb8271a04879678be54cbdb14c021e19ebc66e7a0403ff1e5d2df50c1a218a43946b84e730debf3d53ddb7d423b72cff374273e47b5b436a8e8cc8abcff23dbd3f02298a74ed4dae593e3fd82a2e5b1279984afcb7151565f3e8b9e01f92e4471747b4aef84116a7cda79bf99c53eb42b9b1f0027301f0b7d5baed4b33ea2adbf1f0841b9a7999cffc059c5f07e9f37be6bacb6837c91a6b46c0dd324fad02d03a9a43b9aeb7cd77c4d7f3d53d2ea5991745133fb3aa2c5cc27f50b41d688e8d529a31eff0b537d85debe2cb16b7aba0b500440d769119b3fcb4b1ea282610dfe8138e82037bb7f37b50ef515acb7beb74817885db84a73f2e4da1b67c8ed31976f110919d98c0a81d66eaf8cd8a7231354fa440589c33ea9a11aab92ca5e45c9d8f423fdb26c3ddb4478a86d60adce0a0a133c40e62f53bb6d29c04719db2164ddffb1e8c23878496ed338d3a0b659566445d0d32db59c390c2e384c84b8f58a70d52734a51e8b0d06b3f654ece501f36dbaaebd9ce633bb49916de4a19898331f2ac16ff2892fb9dd84c74e5e6c7145b3284407459e9b6eedc6670f534233dde3c69579320b08d3ad6585807749fb342fa2b96be6e6a6239b2e992a8074fe4fa5a8130f09d733ac71bee1810bd6e4ce17df8c76edaa4243598f8a3f0707f2ca5d0fcf453c9c3804fbc8a9e25b0b4e1ef8fade4870677f726cb0068dfecf975316f9d046845edbb44f815f503e82beeb7701cb5cea2ab0e67009adf3acb7caeeb60ba5cd68c801a4771d294396ad608df9b4a709f8cfe294b2e4a81af628d76e5c4461f7ddd788c67339846c22b32319bc8079d163f943832451247dd0132963785ac9b11314c542f4690e955de21f92c23fa848e746b82bc3710584249b7fb104ce1288a78f71b7d078acd5bb1e1b76ff559adc4b851cb23384e0e218bbd0a863245fa0fd7a4d3fb7cb2b263e3dc70d704463bf0a8287a81325f9077023f401869a14d4bb33128a42f399452944fef01e7971c9e93daa96081cd92ba1852049ae058c660d3eb3d943028b1aa01588dbde7c72f79fcb3c0fd18e307165790a2e1b1195805821e403dc39b9814fc6408deda13fd50b21c22bb87081d1c76368389f63d32dee3d765b61a0ed189013161f6be74f98c76678bd6458351134bf0924a94fa529ecad6bbb636aa3a72020b3774a8d0e76ad9df25adccb853b7ab94a24affbb5f5e626d0b48d5f2ebe0859a583fc50c817d4b5f6b64d9cb9eb592d94cced94092230d8c4846e01b1709c4f3c9383c44633bb467b4e63eb32374361e443551a6d8314f3c0320f4113fe2faf63c0e179419e613ef3a051a14d188cc9cd451aa44f55ff01ff1fd274739d22d2378fb8eed969b9efe010db473825858897dcf24954b98d7afcdf4ad39c168c503f1f0f521c60c67545a769c47751d4caa5b68f3fb2a9209b1da37dcec5cdf79bac43cfe176946c71df13f94fcdbf9675bb6f1fff97781abcff9417e1a713d3243e5e595b037b81af798a55aec3263e49aa291c458299b4ae538d85d37e53940fccebddeaa53613da1c72b501fc9a780939df59c8b28c7f7a0bacce382328fa42c1da5b81645c5ae9be6e7ebaedeaec0724a29b90fed3c517c0027febb601957faa2fd3c85ef122038580f51a280559e1a1eeb1e781c03648223b1c7dc56bd9be8817ed3bf3a3ac9e01df110a03d8295010744c325b8cf4ef693d99582fb275fc537e3acaf23197a8a35d1b1b883ccfcae0c8877629c8be48756c0e5bec8e9210326abc35abde1dc9416ebd1f897bce9ceed853f3f9b1ab3f3015c40fc55452a8fa02dbaab1d1d759485eba316ec30704df52f046a82933443ef115873f67147974e7ca3ad51311fdd0027c4e7d622ed05f6cc2f37b58222d0d1c50366868b20fb7c893e4932d506ee576e0420f7f155d68e965967e01ec0a15a73bc1107f5d3d9891db807657a74e8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h49d1308ca999e9383d7a632c7cb13b9dda1ef51bc66eb1426f7741fc474bea77cbe1eb72f00776ea3da83139601c48fa9fafc4dd1b5c09e839d18c8dd9c507c4a55a32a9f28ac1e72373bcaf2047ee14723d3b7b8d3a1ccb6d6fe4f8cc7af8f745276350e2a2ba390d372476e6ef2e83a163ce0d125758063b634d474ff6fc5a5077676605d23fc8b634f7cda32db89fd3f03a993679565370c26fa3028918f10a357af47ae872a1fa5d77f95fefd4c36670a5e5cdd8e38ddd4f0a2a96d2ea7f700e5a9b37ec2d1ae837bf541e4f26272aa188735d02c4a3864f6350ae90904f85eeab60202dcef84e237901a0b003e987dcf6604d6208b6e34c95b750dd8a1b80eccf08e40d32f12ce17b08fa65bae385c4bd87993be8bb85af20459a07c9b30cac58cba470eeeff91472fcf38dc705338f6779a718a02226657fb25bee5e4cb58a8e4e6377f006b7f6f5fe6f1f5a2eb89156f672d9b38d0a7a3c2b02e8fb0bb27cfb95d4699a3ca4f2d8647d4180438ff20d7710cdb1bbcdc0e0d67ea80d802be666e25a3d740ca38b1432f3c425557bc0405fa01f37a29125a50b501d93a1e89c1924209d04eca155f13a72694e55e70ba6cfdf95325a2f321ff838780aa2d8f03c2f3df019d3a8089d34b506d10115708a7de7382a0b0e4556fa2b5786e58aa3ef5070057a7b5de61138a3ecfae6ab05c70739dab1b5883c3ae68135464bfafec6d125a0695eca48c7a2af8dc1b4908db317991f5c9474666840fe00663faa18df2291ad0aacc111982ae409f2dfce58584b1e4b0fc4edcb65fbadbc5f5f45a44d2f77a2aaca7e30255991dd6bb4a28708442634d8528e96a0c74d4a55fb345ebe66cee3b8908b800483483dcab3e6e5d7a20d6c00cdfd419a2c1226d528fc9fe2e79a2538b2690ce7805f9474a78804dbdfb67a0800cd5e220f9026d86e6155b3d26454dd5af6e04f7ebea5e6b0dbeedf5c5d542e4c839708c9468fe339a58da44bf9d67de2969c5808f7ee555c75ac2fd94d956f3194da6c13ef580908b10bdc476b169ad74c1b3ae0f7c7a3655e3b2de363afa3f7c240a382a2ccc26feb176c16f5e13071a11e760972e81d79d91f60c1466ccfca2680f8fbcb321c879955d04006d625769aa085198a273dd5485f21b28769405daa48228fe8e9e02e91b38b6e5104a089839181366ac5ee88b6bc91d75279b849b872eb33c2728e82fdc3b8a1fb05f91f4b29a4a0bbce50b61662406a4a3d1481c6d0343da43a33c2ae4278be60d63752be3046c04d63caa5e0c12bf9355a4922307015e253e6b62c764527d120e738b59cd46efebb68c36211ec7b6847652b22a3a2bc1251d6902fdda7e758428685c82267bce33f139ce7b6ff4e0181abd67b3a77b5d09896f5fc47e8783e38d48d843a8f45b29416441f3b8617ff31b39f43b6d91a9da8b8f99cd6944388f0827dbe3f5ab846d9c54149a1667e64e25aad12f5c70b7eb71296bee1e4bd46787c87842548a1537aa0b5abd1927e2deda0335c20955006c3e8cdd2c81ad469bc5297c312fa74a4157eb5762f73b781acaeb8cc7d47cd141282da15a52baf5347aef50a5bba5e2a7331a69448f752b8d14fd36b479bdf2c561487e2b009eddc9baaaf767c6d49259098184a93b5ab712dc9ddfe88d6aee1850fa7cf58901e700b34143e3d84d83b301079c7a932a1ea47e321aae9dfd969311725eed2d9754f2ca9a23548030d71b1b30a6f6750fdf022af8a6d8f4da7c926ca5b150fd3eeb03ed412f10d02de21ecf467e76f00ede412e299e6f37de20d255441b83ac99e697650abb32b44ed8e10b88c1e0beb17d00e78137e0bfaf9def24d9287dfa57fe9c51403bd5b778a4cbfdca0808718a066e1c8bcba150b7d40e0657d672d5bceb2279652c048e1c51bc1412ed1e50e7c0deb4fb450668e300cbb62ab1f0b2213d7ade7146d820146d0bc091b4ebf85f3803cb788a3f4ae36684b780a6a63378b9d639f21bd0b53dc6feed0eb97d4d5d4314935b5051771dd15109166245b5077155a4dd508704f797933ad5d84829b472b402f35ef3852fdd709d598d58138420510eb19f6fefb40cf52d41f0066c484d019a62b81dcb99e693b27df1caa4fd1d3bb0856353ee01c27148f491bec693c81d8f5e8b9ab0863f13c5068494628ddb641218a3f8a5fb2b0847d5e2b81569f855d6b066a66e132483f1b5f4e557309a5e8e8d40d42db3cad2c90f28a1a931fdd1bffe1837827fb91df34b3890d3f00b4c43ed32f513f954232af2fe8d1c568842f971d6e5740b7904f088c58ab4bbc74127917d956ae60491c71cbc8e2f85e097af8d619519cd82a6ed4c4582b43b1566cab435900f6390d685028705322c5ed16a818a1c1497c2b9d3ac0f75b892c20198caa715936d08e63afe1c72e6ce2390af914495e7f44a8f6632324434e4fd966a3fcb867e9f99de79401362fdbc59a76aafa67f71fafed2da2720b048181ddc8d102f15c8db0ef0c299d5322581b91bf4b3d7bf9e9a965780fafcacfd9a8ab65bea9c0d0b09842f2600a06fb3b77c3a9881dd8a00fbf26d12187dbc30f9c468f2e6cbde833b4b498a2c783b22d4b3967634099a282e666245c5b3ba4315e0ede73cd80d85a3d1ce5e6f655f61b2a1939b9ce33db8a6ee2428df78d5743d94703f3e23288bea48645341d9bbe5eba821a09e3c01103f4ebf51fdaf6c86e8e849545be42dcb7dfbfbed72adce0c089e5a1fb249c12e3b15a417cd31f57b3d31062cf135fa9cc92824267a660c160f881deca299af0cd34cc631f515a7ee341d1b99e809d8372dac5ef7a81b9d6f678ea3ea38ff2f90109d379652eb4b2a3bf842d0b75cb55bd924bbd627b8d142eeab7e731184d24e9bcc32895e235;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h544b0d91155b4dab0390ad3d04976fc7bfc988e2ac1fc19267541b9fa5528acf500a9be9f28224e7fecc79eee329760dc6efe724244c9221d2d119432ac31efe661acd6c48eb3315c3254f69575cd12c765846dfe4caa3351ff4de7fbc434610811a30a382ff787ef6c71efe65ea5643e4c0d2c83e74d3cc4a2e8490bd0f201fc4af95c1a12f55641f567da6979cabbd98f035730c4dcb12edc0ec4c9cedab05b56785fe8e27472a7bb81d7d688378ac752f5a920963605596bbb60a48cb7c8fa6656e9f54448dc9111dc12afc6f6622c2a79a96c9929aae9c88a71f96234edce095acf5a37a88b95f1064c8144d84f01555b51f3d0ea0780b264849cf4e80f70d16b2d348da341c8e28b7da48b5c9df6f8e78d3dfbba047e8fba11e40916fa2ff4050173f2836e48cd618a8c6ab850e89535ff1957df94943b8642b563f16b6097a7562696c20476abbbb9556fd80b0fe6f38a17489f044d417422bce52f60174d31f43fb6b29017a8a4f90398863e9c3005016aecd3a4fd52dd7d3d0d7711f4038094cb01c7e6dc416b6fe15663c3b6f272454b87470ba181b163a5146b6bd2ade8d70065111cdb0025a467c2b72f7f3828be90045f02c611def2e6eb276578dcb36cb184de24856b225d676dfe950e696edad5f24bb6551b3ae4d68e82595c26d2031d72ae2911a7c2d8652cb48d775b16b12e94ed315cce2cc1d8958c41c4a2787c697d8e2390cafd39e73286e98e656edb5ba32ef648f28be64af17a9d5633728619265240a8d4bc8a55ee9438d35c28642c6706d07789f7c10d0de6274d2ae14c524683776eecffde979b58182c6c8cae4313a7db21a667b3d06850fdfd2b4125d1ed8405c630737c10e3817b414d3c1aac0a0a0066d20234f7fecdf3aeb0eca4a2d63308b45b7b8cf4c59ff9c8c1612a7b5b65b5f8df41bea726d13334a3fa51fd08c1dd6ad5df78ddf2f4d36503ec742a6c6d117cab09fe6d5987cef60fae0a4c662571d12358315adeea1e6e9670e6f0456fa6bbdfdd8b62205c25cae23918533f1cba979900492697fd50354c91a087e627822b104120bafbac3054021cd4a8d95684a06eae6dfb6c74f80150550d45814fe799af9d40bf8ae18bea0324fab76d7ccf67ef681afb35b06c3efe02b7b95eec44ab20b97f080fea3dc152a1f636b4d1c9f4a1ceb75bffe408cabcd716725ee00512f696b5936f333a7f7efbfc4fb1cc7d793c04e30cab7e9be0c66d23e6dea06aaee5d2ecc6dfbcaad8407af1772396978f816fbd405571ecc0a5a6535862178d1a199915ac7a080e35eb946522449f1c1eae7c1807b684344738fcebc1313d8654b7ff3a5f584d89e379fda9b6310b25057e40e96c3b1257b512887e67da9057d9dd9de16c1d788eda76b7336369f52bfcca526c99fad79e2651ff5d0f75dd803c5c82da1fcb4cc2b5ef8ae081d3df1fa2bed940ca6f022522aed418c9d48b7cb04ad9c604850dc38fed100946f2245c6e7a288f9ddcc86e547ad8b15d42b13617d58f04e8c289a6bac72884f5030812ceb0030365777082c38c7b67907d05a79f62bc76eace47a6e5700dc2b7dcd9621e4e32523c2292dbf3b8ae976c3f9d7f16e06c9853844b6b8d17a1ba9de024013666d073a7dc1e6b99fc6095fc75bfe5bbd3445fd352ccc2578b7b41775ce66c388d323d12a31fdd04ff1063d36653a0fb4ccdd1edeada77d109ee732ee36eb3e76d8534822a1a7d4d7929adfd6c42b232288ae208daccfbf190a6e4c83e6085d1ddd4cc32868d1491a2036b67f0d90bb4194aa06365470db38c6102a603cff4c578d7483bb9cc3a20357bab51bb2c35f116b821522244634833aa835fcf4b874fd3d5e08950ea9d37b8f54355af0221b157b2b85d17e40e3a3be03f996c88ca2c9eddd07751c9f3312e3dc855edd92930af04d6137026927430a0dd0b4649bd54247c54d8ebd973383c366c8b75c8bee4801f72346a113f334632bcbd4c544142d846c963ebd39545b4052fb4f47d275044494fedf1ef0137bd4ab052aba4b5f0ff18bed372844c932b23193270b729ed910baa25c0b5df832af243d7a0ce0f213612785b292ff9faeefc5c7e71b3883dc8638c877f1d962495b417fcc5048ee13312170328e90949920b5d6638818bd55480965a3da4d615082b14f99630b3b72ac0039ab0e5e9b22ad05ec4ecc25af13bfa1ce7428c56c21b10e0a34650ba91ff318677f3d703d60cd869504e3efe73d681f97b640ebbfe1e7dcba01edd97a691c391b89f50d025a86d59e19ebc1c454a4be7a699b5d86b08e0522433845c921e808e1da402abe5978e6042440d7857381c405f27f0c88801a2d9dd24e268a2618b88da6ac95af906b66692e25c5190ce4d0471e92a1c9f28ab256d9ff6a9188b721124967663a09dc26ee5cac2e9b123a713990cb224184650f8c1dbace0eb168b49688453698a2dc13cd66a3e9be5ca70a89180a5bf9900bb07927c37e2ffbf73096d9a081c75e1d3c9dd2972f2c40963b03e553227b32e4fe5ba756c11792078736e9cfddadd4c16ab0123a5aada21f73ccca4ad66065a3cf316dc7d16a34cd7bb92e82d202aba61450b43c6e30d11cb35360936d530c1e54800c97342fa191ba95a3128ad9bd0c71c44bd394336b2f1238c65f41a68ea1796ee01da5ac016d3b6776c1bb7822c7e6a9abaa8ae3bc48015f837ff3342e5dea7def3cd59ad385f95c4a96577be352fe7886ae6bf0bca90e6b0e895e249005fc02f56a43a83731ad1437fe97bc9b24c56dd637293c3fa84a8e872f2273336555e75097e9790cc6a15b0eb0e8a6291dd989a4bc9d8eb890c32eea19631d69f1b36b6c811f658c4a63943bd1fbae9d77f302c0fcbe1803ad924c78a69e39;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h24d6054a3061e58a0771a3d8c06cfcf445e6482ea63e21f9e97129188cf1eaee865ed7d08bf776c3267aa5ea386f3b45dd071eb8ac5f135a8e93eb0f70e0c077c3c49341cb2f8bfbba42f2862fabe01acc4b3eb06922c3d5116ea49b7e69e361d58237be87c24b9b9316de0ceafae9c5c0f2d9eef39a3424f778bf22e9ce1e280b38973774fbbb9bbad70710ef3eefc8310d2b170647d76f49fad8fb8d26082c01bd72e99af652153523d7941c01ca53f64985fcc2700e3dc32c8444649e32fd28963e7a67d649d271ff334ca3175dbd3053d53f946af0d7c5726209353b31894b4647fa6c8331805a5dbda1fc1788eff28299567e2d0b4a32f7e527114a143089f9420e01b6f7443a4c1fbab2249d3f8823c695a5980e5c103a06a255ee971b5b776d08dd5cee030e0aec1d0490fac0ec6b40c49469c86f699ca84a3af99deefe2e522cf687b0d3bc5ca734f6627cd3f43fac74f6b862cfbc323080c5b01c99dc0988be31cdb5742294ff1be279c7501cda41480413696fce22dfe371be81f2c3c9457a94d0965f2c77fd3a447fbfeae0c3a16166ff62cc6bb9c295297c2227a2bb140db735ba51b450bd61a39d8664d66765a5b0bfe951235861a2ed497f3d7d16d84a1ef072fa2c7af1e7e0aea4402a3a9b9054d070d1e0e6597b7ba17c6b34e8f252fb1f028e0123b78a7886814bba54d53cf6c7316d6d13db22fafc04d54ae42761bca04e0f074069ef31bde82800a99fd0cc858a47c91ae7257ceb56b7c1781ba4a9e3a3261fc6a69381e19a8dec6383b086c7fce193c2f341d3a23c4d3eb2ba092376392783df83565178aa65784bca9f7bcdd3565601aa5a2e5f3ec5902d5d22c1258de26f2f21d947e13eef12c4e80ba268e998a053d91cc0989018498501ad5321bcf8b4364ac4e0b6f054a7f8534c2fba4c5c9a0fba1eb741925d3c1d5d638aee897ad7f4ca1e091d58380aef22fe8426323a06ff72d36dd1e55ede4a5e40ed226152fad16199a7e4d842d123b584c7aa373261eaff98fcb95b44d2df9da5276ba7341ff8c6898ec20750f3ad4bc4e8ecfb362f1c7e09694130e8143fc58e0d52b9baa7278ca3ce7ab5e9fd45cbc7c7020e0bd5bbed153aee46bd337bbec8199b6233a8cfb6aa9a15fc25b422c89df2df9c442f33b0fa31df87c79b7df7afd4dec0a3ce106b17f1ee1189887a667fafedffbf613b610473c44e9fc1f0d2c9cc3f33dbce5d8395da908d1c81bab8a2da895cbc18df4de3602bd8577dd938ec5da7e5d995d2cc3b5ce74dfb595940b0deaf867a4c26190b297357b630173289488a6b623c78b99a633d1bd891e82653c13c3cee1281fbdad7b0b8903026767fe31656d166bce0c3f2815c8bf26c33470f3fb1f7258905fc8b81ca58c2eac48e596201c1f66f0cdd24452c98d7e59a9a80a3befede3bb535b1886d8b5ca39831187f8dfade883974d225e8e21554b811134124c2eb01e8f1300909b2fd41aad009e1e0d64a89a9708abad2b3ae6c10c5b3da0c1b2a059ca7d1d78ed2842019341e8874e2c1af5a26d1553dc97da7ea2748e8450d1040b841ac524e6e9293f2e58016d64874341653c1db7cd68a1832bb7e41de27d8e11d21c5f59b2f2e9a6a109cde0302207598e57654ae89b3d76a116a608635773b4b3349b28474f2e85b8e45d3510a7432bf530f0e06fb39def244d7a82633b34541df0fd448d04d694c81b5be545ffc2cf306db7181975b17224bd9a9d52147eb9ce6d7ebae73e45ffb2e9785d5e7861ab00473ff821094378a009c74aab0b2f24b13b34721263ab603c5c12d01e8d0edb57e05bd209787f85eeda478fa6d554ffcc9618381486551fc17f6e7f8418e4947ffd5e86c118e0dda9b59526afe9eb264eeb432ad19e5027577008a68050e9de8697464247b6c4e07351601e8bbc348be8b3da5a8df37dda39ea7a4e6f380b79a42369cb6188d20f20df9c589043df478be1e1eb8bbc38ba23830a6c5e988702b2fb7306160e23f7697203ad68f5b2a82c7ec9705e159306021ac000bfcc560d01eaca6a463be018bdb684ffa4e93a7a0d9c996ad74d81364109705d4b21901890fd3389bc2e655306c7b63596b12fb4c9fe5f23f4af8515a8fdfaf952399608a4f7f01d88ca736fa702945e7d3d83ce2d6b73e28f423dbf4bfded2364351c2caf29b1f0687320f804314fb479e6c8ed1cacb077088eeafaea111ce54cac69ae2adc48ba73471d1eadea8b93cb10b95c8b3d6df6a76442de1e2892892a5e74455bc7ef01e6cb802200e35831876241187b6a4372fd1cf5899aa9b6d2aa7e98ff88fc4638152c584a6b850dad995f2149cf423fa732a08c16d93d85b4c319f06f332c478a0c9c7c6a3bd6c5a7ffffeb5dd43e2d10394c8e25204528cf785ab659c5f86f035225f4230ef440e6d54ebca0849f674c59b731a70156d6eb5f29be0e3bdfbc58a7068a7809a793ab8598807d9db12aca87a0400d2a6343ab1749ec15bc716bc15fde285c7222b9937105cda9f6af6f2b15a80982870adfff0403ba5086e378aa9d5adbdce8192554898aead61e15a90eafc2b04e72a796f004e0dab005bcb507ef651fa468d04a428ed3b1667b4884ebfd4a2e80e1c68639f379222d6a810d1315ab18d22d380f68bb175eaac83c5db5091000535840b6104931fab6680521e26cde1ffec45ac993c981ba45fd8b9b4b40f2c7dd188adb5da89ee05478f2f78fb34b89c3c3f5f20a8d5ff05a0d22bf15356837bd0d8fbc906fd578234fb52370bf0e5541c3489a4586f20636c31a05639dcae6a68ac6957757517d15ff54544dfffc90fe341b080b85354a9278e128fdb24cbfb4be5eb4571e3aba684d4c8638bc0dfee614c2aad9b461edde44f210fd373;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h360e3e1b3daa43e45d621f6189a179f9bd33c18b6f47f313ec5347962fcd0999f6b45a2bfb7f2c5faf70ad4e1ce6910d34b391e9fa48ac5cded7ecc8bf445b104462c4204afd796c5f50348d4985494ea2e6f70a45ac1ee0fcaed7a4f935cb3e4e34ca18c0d06ca49295141ca76a2604b847fa049f35b5f37a43d4304d9924d6afe791490ae91287039f3659a184bc17fa2b5f552856e990487546d2e87819e10bd2ef88be80b77400e6cb26bfaa65dfe9e74e8c981622078e025fff0b00a1f6079442de5209dc86e87701034eacd63c0ff619b3b20f71f6357a7a5b36e2f7539d3fd1302cd855813e6a4d32a283f2aa6cf05b103b9a19ffc157a2783eb006df2a9a769859dd2899f9e11662bcdbf67b560f9d29b21d8a7ea1c11aa6ec7ab8fc7edbb7b4e34657f02e2f5a21b4f3aa9eb709a798393a41194e6e62d6e50eca36b92b28631730bfa08500f5d92eb235a3abb335cf695283d80177d97d7c7d84f65596f549f6376031520c16d57f9ba663d3d253b6f54111712ef395b2f3d5f5b17f93d35ce8cd9fc51b46430cc8554b89c8e818d03478e19ff3737c9e8ecf60ac1cc497083eb0086fe2fea69f4c242d3d83bc9e7b906b6bdb756cbfffcc434b1fd7b2b0949aeef74a090463599c862c2582a8982b62c89bc04d3b8932261edba576dca6bdbee5fd8ef000bcb5ec270260a1f2c0f5bd154796472c960a1f0502d6e3f9c2e738f3b3776603786c000437cff4d1f510777b6e28c2855098dc73425c8a3adfd19e57a5d1806118be8338e4785f40b5de471ddef1bf5a945de9d0b96fc72df78c9f002a3609a3cca4a2ff06bd0051b1360910884681fdc10f027a2beac6002174600f6efdef8afe419dc2e0df66dcea7f53a9f09e20126333896fde27acad6d5b79e44a98d08243918890df26ecca8b788fa8e203f8b440c367f2029f42ca83f4b65685cbba0f1960d1be9f9d1a6d670d5ec03bac0486198cb07b71b513e6c918806039cdf5cf0007a5b366af7c6e95ef58bc4d692fb9ca1a0c957fde6eb76b33fafc8c3660699fcddb370809b0eec77cc00317ba1724ad25646695a17a2ed7560bc0b75fe9995f1616cb206ded677decd80f858e0b2b0fb9befb37bacbb97d02c570d749ac930eba80e5f28a52cd04f45c68ed2defa489901ceddbc72fca56b5cc1980b095e34f6733ec2327e1434c7e1fc9155c3e865d6171852e3ddbee6f6e424c0ad7dbe851ac4d0ddb7c832ff421432f6678e54ae975d7fe36cf54c714e8e197b9deda3fcc6600bd5a0d464fc6ea6997c552de1fd27c3f90801f50e28a0f1ea37625c9038ed1dd80e58e4ed7b0b41736a4ebe0f3006cb86dccf6157e55ed7ee7f15031071ea72c1a278de0c956545a1e5b32170bd2f7179616c0f484240044a44adb858b846beace241ecc168a132ac0863dcd74adac3ad307d918ca54363e7fe422a244a589ee0573e04a0cdae5204f2d3fd2cbc4b96cd33632260b4c931b566c552585850c508c5232a4f4aa8933f2133798ed2f526a2922bfbe2e0c8b20b1fbc706d357ca069a2f50fd28aad1c81324b5108dcce5315d75bd5bfa13f7057fb2ca7d447faa7920f6709d73e76dbf75dd47c57eeef577587acba65bae7057b926a161e8a11975e354b9a747e0aa19bdbb55e40b1c8b71f38749a52c6ee60a5e54eeec845ae67eeebcc84c4ad6863faece481902ba5c9690b285fceb5a1d736e6a887359ee65b453b5139531f3354c8f27bad257bb245ec882a4509af35166981f4d13810565a3ad183a2d9b73596bc311641944edf7c4339c427c49f663de7f9e1b33e1dc4c7d7a96b4ac2bf26d455b357a19b7603bd001e32ad0ee678afbce64c1ea9757d16214b1d0f19cde5aa08c1f50cd196d51836d9387033d7ed26d22c48a47cf0c3a19e586a24dc9c2a4da9ca0f2834e2bc612356c226cc6d0eb7bfe16707ecd41396a9271662c21da0377b8231d8367a059b7d7bf3e57414c015ec0b925552ecb05265885fb019b73dad658a1889587f5ec0a2b3a512bec3491a81bed98d348948e88897cb217995ffe133e9e3a74b2435f2f21b5ac4788d919584dd7a0345e74e7bff42427eefc4efd414c7d53864b9322b26aaf537d6043afb97cc08d2f0161749f3b272b30a84145373262af467b0ee6f4ce679273ce708000632300afb40bee78c69ad21dc48703e6028a6633c498539f9613c9baa2dbc6349ed8ee67c344c8254325377b340de797711c16bd8b1bbf75a7f999d5184243fa08d6384191359dbf17c6a1f0f4e441f6f088da74416d892648771aa52cbbca2dfb50f8fda60484589fd0879f81da650d9f2f630e9455977395460461007166bdba0012f09eed33cedf0d6d94be091b755b830b4a15928bc05231e786cf395b82ce434e1fd04bdcdce3fb5a8a0f49125818fec4d05e1f27db8fdbac6a543615080c06bc35d4de1fb3d5deecf95d56da99adc7892c12f4c9360cc84fd1b41f76ecabe7ea0bd525d0b61031156cb050b54d20f67fcafa647d450a4edeb90ed9cce7e5841b5d22d7e4234e782b03a431517d79ee6c593b51bf26425a8e67ef82fd3af3ecd408fe179993ef1ce9c7b32b73394088fc43b334460f7f44298ba8469ae2d5cc4ef7ba79f90263ee42e2d0118af5810722dccb0f596f30c8bac3ad72080915a335bc86864d6637bea3e054cd8546856397d36cd241f048716eefee751a2b97a7b04a51de97d4bda9337e0adff79ed806a4e874234c2eff75be5d6ff1b80cc72b865b010196d06b281247f5a0af784ef1ba935456e949a4375fb14b813f29eb278d3c5e742a58244b25236d4024690357133b81a8643c9400368614b71497101b62eb88ca585ab0bbd8c6ebc602aefbc1405fec0e963149106f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4b290003e83a5566c960f40cc957b9d70df6e7ae445b5b17334248bae19ff183c91b896be30fe0394156ef65fe69ac8a68bccec933692a598a825d21d35ea5b04e9ec2816ecbc7d9a92454b93befb79b95cfc43499b9bf56c78a10523ccfa70395ebf24685a5266eca8589451dfbfe90a8f3c18169a58ad5c66be52c76536eae0bca792ebe8e187ee4b6e8cd320174e6f94b1000ce7719adbb53751287c79d68fb18d7fe1b238e6811be9b84ec7d56f7ebcaf57bdb11d24c6a2d45ca1008d40717b2cedd9019555572b05f0a16f373f7bb2570bd6e18a774ea0a1fd8d58758a8ea3a05cc93659791206bfa1c67102ae6801096974e0bbdec3c329ae7a44e5b51757a7d1e177851f58b0366e1ace6642b40991766b747e06e6340e9da59b76ac2e48ffa54149b3850293d281151c727cf9ec84d48706eb6b982e9cac634c850cf1be8fbf03e667589cd2c5c7b6645c80958858b2e67e9faa2c8a1cfd51a832b0e7c3bcebeb94f47e5e5e52e8e145ccd2c368c7b79788741d78b97881764601e5c754c417c6996ace1fd074bd88c891a4a9328a4a00cbd8478b7ddc7b3e2f69dd209bd1424c836388e20f91dc3d040dfccc55d80235a8c0a8abb46a63417c392206f747443041972cd49b1ed1e1c41dce7149d0abdd4d8f8fe2163fce86dc85506561f90defbc801f86c983d4e83dbf88881f47b84a049ea2ade5a8160a1b597ecce432eb506fedc941e49960ddb1528ecdbb6649e9e7fc445cc292e20ea88b79a992bb63699dc3a5ea2a4251b78315794bcc5464bc63eb4cd88f2abcfd5955270b29245fa86c7c3a619f07e99ea01ea01d98ce8134dbf20e8dd136c32401b47639b484bad64948e03d674615cf8046bd0f4815834e5b34fe772ad16f6697a152e0c990d214247641e19cea6336705917283dc96ab8d02b09079e04d08e31f4e43c49d9dd6e6280b8664cedd0b9ae67dde358a38d1794f72a1e0b78966ec3d3142f80981da067b882cf8ec5321ffabc679b35f83fa1404bde658d36f827974f4a0f276cc294b4c925769383ef57e37e88e8a72e30193a3105269a813b2065a6b0d813ce026e0cceb425219d11e44126a4a7c788692d9b5ca866734bf2e08c1dc8f0513a44c6770a0a97969fe1eb590e5eb8fc93aa6e9664c5cdc54f4b60caba1667df64ad9f1f38039522fbfdc61d2f68152796190de94cdc58752170a0767d0bcfb8f31b668b9c058fc25abca20fafdbeebe8955fafa56aa26d3334de60fe7b28946a949ec392163e41ddbf4af88e54b83e4f28754b15ca2d432b7ab937609d87d004efcb158bc841d008359659bea835a3f89195c75ad3e3a67e7e5480b1b9d0a0e0ea4f42e11b3d7535f9ca1200c6067883f049ac6159edeff3f9b0bbf8d306115d22417ad1d216f79751aed23aaaa77793250abd779fd675e6e1fcdb2fbdec50eb1e140a3d53f75d3d1b2778a578f0f9122cd4a2d6feffc0f633203111f47041caadc33d8c11fd38b2227d224d985aa999ea7cd21c4b5fa20816dc38dfebafdcb62cfba94b7cf7afe114c77a748df711119629fbf2c26209a6935bfdd8169a2bb55d57b31094723b4b5baf930b1d7723d91b8607783eb2ebdc487a6aff6f1dd00ab3150c6143b815296406d805861e7dbfad513c62758941f906c6cef1f74672fbf369a97f76667725c80c23c183346b38504c2c1461dd5e2ea8783c2626910f4e071346e22aee97a25201436980a6f35cf9d2a73ba21974730adada554522f7feccc19138a2e00e0db6ab92700f5533b9e85a2812c3053cc9914361a74cb5d53e5a69fba02df97da49dbf3e3de395807890ad39bef0dca84f72696989df8e0ae33248b03aa094aa632f20e3c9e29030f98a93bfb95399e965cda7f26b3e8caf65fe2f8a86adf8fba81ea35b303881e6f5d2a777e1e36fd84e61f9808f1fc4384bb302aee048f4efe4f7d69bc40d9562d9e9c86d898a98633b3936026c5423b95769d3c089371445c7b7e32bbc9fe23046ec45c51aa40073fcede220533fdd68073a17b9169ddc5baf25001c94c4ca8d198af4fcf4565f700d04e22b2f043cb0f2af6838814b9100f6202e5a2e2ceddbaafc42ef9bbe484ea97bb5ff80e31ce0b797da5af1e53012225d32bbc59b4baf3e6bea8f6a649a5392813ce970a03ee2669c1385c207f7de6967cf836a07607e44da442959fb9612052d0775ffc8d59db89e45f430607191b2d5f0069878b4777b3eeebeab89564d4301f4a1c3e437a37ee9782aaa77b92bcbdd7257eb783ed4daea4a8318f7af0fb1c7510a465c84d34f7894d8010282225ba53ffbdb1cc6fe9dcab05f9f59caf79cdd981d49a7ec9b283f09ff0831d078555c9fff8d71cd312329a0c4ad2fe0be695b3d6317a1996ef8dfdf4c1fb7d1742a5db98cb60dbd44e6720e595e2d21dbbce5d5b628f55c2f94f1c8d25e66eb646a8ed5358091de899ecc4cf1baca881ee989c41984b635b26c3fc7eea4980442dc8f8d6489b0dcf5c944119b7902cc19cbd26b10a3957eb8984e873547abd46f7bcaf9a1a113274a966d98df4402a2a5dd5c8df002c542b73cf4c3df8ac0fa2f8c309f9bab48a3ad7d8ea2e732fc7ce3aa8337336bef3d97f182a8399104a350945b29a4cb0b05e9553d3ca7a335c7b66fbd17717859d99de9ffb0780cddd8b92e49755d07d851d3bda5a9b12347b69965eb76f18d94ea3a15354656a39568b0a0227c7574048a62195a854e38b2129d4038d9e904bd60a8cd585d6847a664bfa5a15d4a7b5a77f5a6e71a5d7d08b554221361b73e758f4120f6a2c61f50aed48c9fca430dd8a9019673d0aa57ca1a7b568d7a350c7aa676c66ed7e0bf20edc09fecf1330f39a8f45a96b653e362b2e1d43b64f2a6cd45;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7f4bfaf6d93e52219a879003d3a26d65f1b7e090fa12a28e50af77ccebd260c887e6c55a7e70cad5fee7c73164992f90031abd92d2a5a292e30745295b0796a717de150c0ce9d26bc56f16c855a12dff0c0db88ac86768b809885f7e8d0f4c22235b6d3e3b73c7a956686f609f155e29f8c17067bca22c6b58cb8661dfe154890d526e3ae38c518d95865836f448c892bbbdf923511762997f48eaa00dd532e3fc9f9ffcc9b97fa56bc8f2d70be2fc829a87af8d9a2f83bab9e615e74a24a84bd8cb42449c22c310925d1fca14e1197d0d3e752cdfd9fa722f686e5ba30fd030aa8caf7b0121db547e08f52ece9a31b8d029db00b457ca2988ebfd0bc7d976cfc6f45cd96f2260048d4453f2d5bdc1ecf21450cf6907672f9bd10178d19932d0d69778bcda88bf89ac16a7695695efc3bf77637d4074b853b22d98f3f714367e550e2a57f41bacfe8ae47c6a1d1ffa3e369913c85f12739413f0597ac4b8b31f403af9a128bd109f459fc391be64fcada2fc6b32191042775eb1ef8b4c90736236bf3ab0dbcc627d400a8c96b7e8a13cd2488be361d3371a1b6808567781ebf79416f7f4943fe8a18143abc0e73fc634da24debb510c8369eab0cf5efe5c5cdf4ec25b4026ecf9f941a8a806b854b12d2addb0118dc7f3ce2caa2b13b8aab402e8212213b2a951593851e657c47985f81c5c382e63601ffae204fbd5aed3234d992304717ec9ec89cd12afcb6a6ee69a305a653441454ec38f76695d4873003924e3b3d8f3ce7f257d1677bbcbe24d49ec110f8eb7c57f8b1024712b279e814c0ad7bbc6e80dacceb0e0d42ad8ea47be04d2c378f709c29d6bd3d4573f28a202726a119179727aa7548cbccbd8c011290d02b59005a896a334ab39a6c047652bc071653012e5e04cf639c9765e40021aac6b224178c91aed96d189e53ed1853c5116b0943186e7d09b2294300083f6fc6087c2f840f28e55287b05a72e9a40a89cbcaf2d73ca3dd41b1746a6dd7e06972798e4a0ef8e24a526b54ec4374223dd6d2df9259869e751bcfb555d02a4d9caad3847acec58b3c513b05ab37c9fb3514023d677b88ca2ecbe23f53c9a143a85d01068804b898d6b6dadf1ffdd694872af6ca8396fe36c582f6e1884d41d44e1726fa352fd15c69b5773d7571c48ff33d38805458b9396eb8b6dbd72a3b4aaa8e764ea72f9aea8a58e37996277d14746591cfbcf93a81962b7b453e388084692af1bc3e6ea936dd49129b05920a22194c6e4bc02aa27187042142975ec6b830c7e43c416eccd0a97f4de8d9f9c868dac0f6d2feaef9fbb4dc52ba8db89db108d438bff9187c3badd213761fef05e8a775fbf706b9ccb2b66f68885913c2e790b18ae9db32d421e580ba3e9639efbc471a0ffd5cac500acecf2fcd6b3599260d0968633011350ab10be76a56c9de50377e694fa2a23f77093571e6497e0e54d6e0cdc69da8087e91038ce2f78227efa61e20fa65f712f4f4856ebfc2f5356917cadaa611a3abc78bc58c1ea59141a63434f19c85fb9bbe27a73051d86e88afe3ad7198a669742b84e95a457e26ce6f833c68ae1f6423cee69e38d28b146ff34968790b5f330d7f9e8b48737391e6553c6eb705cdaeacab39a13071c48eec82bfad627fa234756ca9a0bc98b616334068ac39b20c8455a5d45f147aa1d3b8647ea332dedde0ea8da9c342a962e5487471c3a10e8c2fe1e7b389ba64ec65de45881efc89b8768cdc9dd4455f994c0067deaf157e16b3348a9dbd7a7842420e0aa263a8af68d2ab64adf007c2798e2e64f5f7914eab8665a381bf7a247ecd152ff13da38a2268b50fd92a6359f601ba019f2c4a5747d259a29a4766e5bf5924ad88c7a2d42d7901b5d7cf48be72b7b7e2c4c7df192963647e6f1eb515cb047adaa527f5ebbde670c986df4f650a1cf93e6d5c2e104c35674dfd750225a549e7ab67cb06c2c077f19eae0bf5615623ef28006b6ceb475ff1d0daf43d344578c7baf4bc08672e41107c4356a3d220c47918b45f29bf7bee195bd9176e97eec243c968024ab9d49966a0ea65b5772fc4218a2e91c623236ff16ef104972973baeb7eddc216932c4885e569225e88c4219d98f4709675a2a7d7129fe5e2c14af248c60e6445a51be1defbc0b9571288a52c5800962198222751bcd478e6f3d4da9a5a0a376066fb8e095b4b626cb6b63fb531099030cc060adffa211e5703d52b6298d4215c6567f560bb56e025c879054af180c0a4f98297b0411899f252a714ffc76b2b95ddd202978b93fcd6e8ac39e152b65b5661a99508f87d5f4c52a348ced6609e2552723f459e55ee902b43679b3c92c6a3cf3f7e14663cf6db3b676616508561929fa49763cf55b0ca257033a7131ac898fbd9df32ad59cc9a408237fa46668c323663a46fbe2b7734fd2ab1f492a8f100fb8793e35c715bdebd39bee4d2c05c97acc76a3be1c1c80e71afdfc744d140159b15c3cd0340bd947ca33c0ed6d0e30f27f0bf479e768c4cb376f5b961019500db6c236cb86feae3981c9c41b3ac2b9484d69eeeb953146969a5f7a10302f014e179128d20b913a215e8e5daa682ee3acab3be6a83ab30125875d0985778cbc2af8958bb13b290151d700e30166f189d9287e1bc27c807a2fa69071917035663af209eeaa60421497fdc9f724ddf208168144893a5dc9fd95545dcdb9e4fbf743aa2387a41341c5c5794e3e278d7f9218131acf5d836458918debd77b6bfad1c42cba5591797b9afdaa5fd91c395480e820472ce8bddd45270c26c25d3aba4d0ad30c2448296047a8d14665db294a9469bcbf8ee6503bdc1534d7b6200f427d03fd83eb0caaab084269faf3fb19e90a0b7e31c32b14cd42e0666f58534a84;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdb552d962135fd05d6f4ebe5dc4682c74419845baf5afa7e72e18945444e5fec66a7439c3ff396a97cde6d24abed6652cd8b8235c1d0e4066de048aaa982dc0aa391e770264fd968800bd4a9919b716e96c53934f8410c1ff0f1ba6517316c01cfb8fa44a07d3ca40ef8960fb67b934789d607c176b4d9af50d34ed9d38101d2f1e0bd202007ac8fa5b222d609ea89677d2cba896800ff8ffa6298e0241341c34a4fd5a4bb71230625356a192febca3f6c7c4bd32f819001c064e98d82d2d43ee04b4f21c6b3ed1943efb19683d60db308dcb816994399d1c9e15f7a8242b352b89f8e87bb89a2721d464d4a3249c7239a7e60d17838a265e6c8d20cd8d79376696ccde350a35379886ae334196fce7f4208409035e7d3e2f89714edf8a6a3cea6dc32f57d961d3a65d7a165940a1dc1ddf7aba3ba6b2f9c436bccb4bd80423a62bf4c2e9173eef6887d7310f373a0ad8f47e784af16493920081b6ae888d47708e3b484562ae734a70e15597e9d9f4443b9dcb546f874a2dd947f5930e6d940dfd81238db6b1368e2bad44263ff0ce6f3ed72971eb285f06a512cb07456a1fa8c83bebc7aeb854334eb646db99680f157ffa321b1248f66fa8c5c1f9e57e820e60613a57e1ed44b88d282fded36a0d6baa768b4947180b2512988c20216db1ccff388c2ef5fc404537828e2b21b29168798c9691658284676585950219335cab9972339ccbfd2409f68018579b4ed166cdc179dd7078fd469a406442902283ce17ae73ffde3b970e95223014b9f94595af6bdf6b54abc039b2ab864b4fbd662dd2d201e6e67e67abf2a17898bcc1b020d37ffc3c3c5bfc051758557191cb948320975160b08fcdaad8d3d7da1620ece3844a1ffef68b834a960b0d53b110bacdf1d6dfe5397cf6d973fcd94adc739742e8a07f0b53cf68c7568d52b594daf0ee08c519c6f0b83e068ce88adffb5e2d49b5180c95dd9c2d06667b22d722dc87142110d611c5015a6fc6c57093084045f9a7a937779a68c12446dd5e32c7675489fc11822184252b02c2ba463758a0aee7d4431b48508c16e0262e422ab0a6af16d2abee4e3f0ba453b66713324c1d5c48d8cd54823093124ddda82da6ff555a9c22f2a53c56e641e99bb520aae2f1311db9a09bdd327e8f2cb4e8a5a63ff72e6b14ff7742a3d2d664f31673a6b5d0930ecc0daa90e4d5e3008e990d69b44892fb9686cfb9a168f0508a74cec7588aef58eb3ab56ff493870bc2a6fd8c958301ec51fb57deca4a03f14240fee43ebb8b45bae2d79d37b399315dcee22c291e2055f197fa028c0066bae5ee80e13494fba397b12de38b530e8c0bd0b8cf0d917e7878e4aa2f71b07417f79cc3e00e385019ab6359b392dbbb4b1116c9e7b9cae84c8e9b0a0af85aca5b284ad6f57565ce7ea77eb02993a3063b65dd5f47f166588d241891e6ea5f98b6197a219a545491fa9add327759745d489178b326dca762c25c430d4ae9a1b2cfa28d0b92973b4726392fb7132bf9f3452c72a3e99bef9ee18c5a11f084cf9927f10910937fc5a3e40b339d2b88e22b4ac55216b00af89521cc41ce08e235cc23b24b368d48e6795a55a2515edb3d3fede66313dd3d6f1e6cd08fd55d26a1974bd9fa9f540d0be42e0382bb2a2d13517a2d7e5318fcf2868951375935a185ae3a11d83079a0e961aa74bdb744b2aa1a3e14286c3aff23ca869689c413c887c534b24b5077b4da4aeb2820926be4dc5fb2ad978240629807bf6682bffd23953c01d1fc5c8e57d4b4c1c478cef49ef79f5cb038f2ad51dbfe279f8f8cf16cff7c4ccbd30a890394d036271ecbd986e9bc9290f36b0d8a4810d39fa5e93fd0e8ca1dd4c315c48f310495b7f842b0c28061ea771ab02f611f7b6da5965adb08c1b07630aacf3e1f56a53f078ea3bab122bd9d6cffdefc9e33be249ddaf6536fdc19fd76ab36780865e5c7aa4758e208c450b6a9a86f03f5cbb4aafbdc97b14e3b664fd451b0e96b4fdf0ddb4f19b71fa829c471f901d4ff9d2cdaff421ef95b465899268ba31983fbdaf9e54f77ae7da9b0422acb37a3e2124a73af6eed19d655865d6b4b443a678ed40ac203a0bce184bb4c9c510f7cc80452690b81dad24a41b4c5746e756d9fcc9ba542fa4ec440321fa9de20163566ce2d8f4a4831794aeb8beb34f41b9b2cd055c32aa259a27e9edf3921592be8a4aec62ea2a01893c02fa7247d008ceaaafdb4e2e45577bb74bade3ca62009b73fbb070e3240023b4cceeac54ba2fa317345c7d6b2af682cb03267d6c75da21d11c9572361b092e897613f4418b3cd2956b9a1da4d253ae0c60350eaa44051fb414b512059d2513e0a594aa60471d0d1fb4bffcc6e7a279acf37ee0fbe3dbfdac0f405ab7b17f52c04dd212cd8e7a4e21a192b8938606676c731e8c87edb52c0eb1e69a8b8e22beb128c9baab8c8b6bed44d4d463991835e647fe884ae5cda1011e3562f393b3ec01d1e34c76f5d073c85753d2ea8d3760dc59437fdf271edd19af7176826e9fc575cdfbd8ad9b7e642be1da81206b1f09b77314fd9a7195d089c8ee5b970fe5d944a95e39161cd6c2eba0faf2d76580988c144f4037cd9cceb8e444cc2666b04bea70c544ef80210ed34d1622e414e2c5edc66a35d809607162d1760928ff5df62e32c97f687339d1f6dc63a06ad4986ec4413c8023532addf1167bff4594f3a9957d26bb64302aa6a0fbb0f3e08dc1efb76ef246842153e64dac1d14331737628c50d2005dd41e99d138f0b8bacec72bb40d583645fb524682674a21dc14aa2f6a9561613c250b03adc4ae7dff2221801eee4c5c7c5cd84535471e8660804ae91dda4c5e899f971988a1ffedf4f7308e7641292a6547189833342c6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h489b4e7e4ab94863ae4d6ec70f4f244744883171d709745c73568d60b75e36359aa6dfce04a1a695660403d3ec203605ef3176b93fe992638972883f224d3a8590dd18ed424d871c8c7264faf5fa594af2f38335de25b86899760e9697a9c5d83221676e44dc7c521616195dadc61dbc5b320c1670c5d81e13f1bb4a0713e996d3cc766762d320b55bf7d1b0f417fe073a3cff23cb7873f228ba0f12b765243dbd02fc243cba67bc0995da022932751b5c4b2dcd35793358bbf71a545a71d2987a1948989de4c7196827ba46d627302311ad288ea37b4cf6eff32de0c7ea77073ae4b1bfafa644f3667e8dc90ca48070a7c2e51009e49eafd11b2f685318ee3a9b1a8bdf66a2992ac5a73f6fa63055a5be907b56f31690eae53e8ea92acfdc84b2d779c9bb9b8d99313356d96b9ece8de9d448f60ae36aa9a4286c810e55f2a36b5fb9225659b58dcd6b55351661390e72943e40e0aa8db8e51b1f1da010e7a6452dc1469c03f7c58f4dce3c1764f607a9e10fd7f95750977a4133fe69c709be060cbb43bc84020ba49234fc9f1b005f7a6b76507443f054f0ba469619aaad6e314389119392207b092f60cacd8a29a26108486842baafc91c356792a211ef2febb78f6cd373e38a5ae279304fc0808a5ad6593b6f219364b5cbe8f43007a4a5dc363109e988420fdc358c33f8acd81271cd7a02b2b87ebeb3198e21ef8be066bcca0a1126f1ada4216b50a19ed0250f2686d0680c0863cd039df657311fa6afebc126a5deb3e2142c74da7402c68499a90527616943bbe26db2218e8d7da7eb19331ff666e7f19d336417b3a30209bcf32e9c1fdaf037d738f0129047e37ecc701d307e96c192920cf960c2abb53946ab4ade06dc98d72267dca2b715a5c2f9098d32d2cd907bb738820765ba9a2def67183d568f8a25caad3dcbab6c66408d95e2da77b1677ecfecabdadae1ecf16b9c6c9a9d3d9ca3e8137237bb78b450bd39a09886a2aefa4d440bca29604e01a10cfebc45c5bf8a96b650308d479fb6eab2bb24d602eabc708260aa689302316e2679a169ab4274a11c5ded3b42d5b6f8f8daff038b988e9a8736ba6fbcba440b42c5c33f22aa5184ee029bd951b1a42424e2acfe6f8db02bb134da16b0570d8fc1501d6a932cfac5a0734ea1c79ac4602a64decfd0b02ec0cedaa2f51090d2665ec7bbbf340f9de446dfc7acfb47b9ec51c7acd01aadfdfb663092679bb36d7ea31996e93d14a3ff0c48f63624e4f4055ff7369b0204fe0c051ed9551ec9b19bee6e208dcb9701f459358c4147214f546d7c0b90c7b7641e53628d0f17db76f2c305f3bf25e62c9010ceb4a4a47efa6c25b81be3f9a7caa61b72e6a749771b5bf8ad0e1117694a5df764e35f6c63b7555b69fac9e54b366c6ffc7000fa6f2ba94e95d76316b45591efdbc9bba130652ad3d6094807738603a7b0eef3c8b131c317edca02ffc3ef2988117e73f47578f2546c512d2771168feac31e5edb4e19617a47ae200d0ab281ae5f1dbafbc92193107166396990c04c6adadc653fcbd0611ea35a8c922a2d66e13a8fbb1a553d7bcd8aab95a506cd5699916bb879e6c20e7739dc32ba46f99f548fcebbdfca0ede6071da14e68e6bd700f39daba40f523516a6c89d75db63234f875b03ead2cd239f92ee6f8bde7c8abc37d4c9cb93e30ab8d636f709137cc1367b964abd93512f72be3aec9fa71011d44d3352149346de27e9367d088f8bb587afa0f1d9819f4e4d1aa1a3b3a3b73aad88160bc5dfb65ea34b8d55e5f41ec8302284f9ca43f4efb2863e9b5bb758b7ded3e745dcf88ccae9d1e2a1d2d0cd79179e232a98936b749f518ddccc9a889a35b786c320974a3194b1d053b8a991b8dd111e97c938650804d2d8f7f6d181a4876e3c7e6095a115e2972ef84f9eae2a1a68af89e346aae3392f9f6313db80307206cdd84d2843d2f0030b8884465c913f8b78cedfdcd99e5e2a04ef3d5243faea196a14acfe57df77bcdd4bee4b4a32e06902eab534f7397c6094cd4046b0c36db3072cfa5d6842eee7dc691cdbb73281b2ce0ba863eeea48885e0a151ead8f69b71892a60d00a79b13c350727b03b1a7677f132d8b0591ab866d13faa89e9dc4e8a7439aa3727026f4e2adcbfa404fd3e874e192eb7ec16a130f5d3b2c14d9a42ca8664be45514c9e6d55d3aa287df041bae0b6301b712b734f75eaf090ac7cd810f1a84031110dda8e04e595c03d3da4a8ffd79a97d5be2c1adbc075977cc43151f8f9f6ee131b9e52f151ea2781de7eb81b94aa244761df70ba79095f9b9fcf1fd89805eb1862e3c79bd5f0c836aacf65dd2fa5ec5b8ab8a539bf13adc2ee82c3dc1df0fefe4107ee3382e6bd2a32fa0ee88b2c3d78f60d646dd7c9c0038b20b720dbe65ee9459502a8ebbf437bbb16ebf1e01362759a80a35a438dff35453f8121318bba6b8b8859e724e45e1d84b72569fe0f8183f35ef28e35dfc88114d7274991a7dc100faa0d20e5b2d10c2426929d20c4501293233cec5507b0365fede584c62f5f795289c92f371d97f6b6a154cde84578f8fdeafcf95ca0cbd1e1b2b83e0c1c0eca24e7d46e52b317e22103302a51d331d2078c06c0b57ab5cad3839a3dab989a6a30e6adad74555ca6e9c7d29fe4ca20a155dd3a0d1a15372a660c654b8128e3e4cbd92f7a96b07e2230a77fdba04e11d07d947e507626ed297a8d793c533a7c992051cf012fd73830a72dacae9a184b595cbebd41f23bf160460c9a468ef6739993b64de2c7a59111703e6a6d5f3f40f2d5bb659a2194505dac1f6800d3eaf868b7b3a8a522e1e9d3295d1e3204677d8dabea399b0a8e696400655a2a59d99730d50f0831b97c817fd2fbf6f8a2c3fc5e3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h7b815cb4ae8162824e865bd8ad4c31c5c00a74932dc5d40851100b0ce1c769d27214124b2fd3d04c842588a6dc48a6124da1e63f3f92737a8a40913a119852f337b4ce3b2a275a79d1fe05f615918a02c1b96ca1251ea8e89f7b04b0629aee13238326894078323426f5fd9a4d40f25be89dba27590a121b70dfed280ec5f2ac0fa79112ca7cf8bb5d82b917e7b9b7abfe2d4bb75daaf341dce3fed8164e5039e9746d5a0423c5880fee32605d041a464436c05eb205fa8e697276c9e1b8518d3764bdf07b02944f5c170d403b47e7e018b977f947a73c64a638e9023e953f2ddecf68693d4f4b66ba4eed825d20e549296862e49bc4b3132bfacff1c34ccc81d8067d283f7d9f4edf37d064e6c349924a3797b6d0daa2dc099ac7f07d6d617fc70598136a69ee25d235922f21afba840d727af632800aa689d24ee5b3001584f51d26801cdc6bb67405353aea83d562ba99330710206eb2f7fcc663d17d5ce6e3fe27ba9f602b84cea0795f45510980330bf344cc2e38e947eedf6cbbb002dd3c79765d836b24933baa8d6eaec8f5008225b91e32dcbd9075de85e76bc60751c56fd6a79a760b01bde44c2bc9fd47537f3841df932e8969a16983722c57590020187d88a5bab698fb07dbd2c43b5c2d10a9023ea5fb04d87a3ef359593dd6f8325c5ec9ded12cc11069bda8e6c041e4c8b2fd3b87fd8926034281b94378ce0c9a35d70333ee0d8e546bca425ddc61034895a9b3a35f28715f4a36fb6de4c8226855ad3ed9ec67dbf02b1b4245f0d0f96399143368402c35e84576bb941a4b9fa06231ea7c2de69bfdf4e875dcf27cf46d7fd33762f4738a4d5168ccfaf00d0d96ba9a6b2297c1186e9fb6d36a4d2e00901265597c9923b18fed68dbd83e0083eba871b4451bd8361af96c317fb190f78236c0e85f5efd3c389866174253e2447bf01014ca622be84c9717c080473541e32904b5eaa08da93a5a0b2dbcfadc632b8464afcc9a2b8cbe1b923a361f4eee71ecb53264679585f4592fd17905fbd4efc45ebabfe4d25b4ff332eed91f3ce26ea426761d278aa8de591525ee432f95cdf5a65112b5be88234c3983ed25fee577ae69e2ad9712f167c7c443999810178b17313d50b237be61257ff9b8c370c8033209e9c7aefb2a1aca479fb97a451bdf691a8e01a6176c5044bc25d4a0c0aaee279ca4bd49c7de8e67d313971a904e9e05ab97ae6a6e387ed3251b532e06206f0d2165324caaf9d9f31b556b412fe9681c529ed44aed210e203536fbeec920dcd1d50380d5f2cc12977551ab46eccd0fde1cfaf30fb085c0448ce4da30bb016d433dba6fb7b0407a8f8ad57243ac912777ff5671a220baded84c2b7e7914fbfc61e32ab74b660ae352b4f709f2ee0e158d7c18193dcccca7e7feeb95de090f8d6dec05709d86237f02ad5e968fb557705e87133cc8e5f496b868eaa88c9d29cfdf1689e7ed77d11e7974c95add37bee9a693fcce764a5ec4661cc64fa8b6f20a4d3c89b0feb7d8949b6e79b16f31f653bf03f56e5a386955cd0d92f0a881a3684bc21c05fd8f22e86e36ca69631e6dcfedbadb77173e48bcd014a8b7c76e10854cf8e5e0cb302d507e6ad5032e31c48b0497abf30013c5385e708b216e2301c101a3992429491dc2cac52aded037dabe940c5f7e03d92b14ab2ffb52ac02fc9d88b4523b79e5095a9f1fe47fc3ca6bf0678c01dda1924293b8db9b7608fa53ad8fa5842ecd2e5293ff554a8dd01b8477fe2b97a0d75bee886cfafc29d4a415f490f95c38006794c18d8d53056a64787ef9e0115f01824899cab18d0b6210cc32f0c6ff197a2f381eabed6ed9b0979ae0e4f2bf43565fc26e00d79320ec200a9768a6985d85a0238c0a2acf4cf58550bd1143af3e9e5258ef831328b692bef19cff8b57dda2ce01b0b5ea417e47a445f5a7e39bbbc68b2ceff5d3cb237243cd3d669e62502161546ee795d408c4d40dda1eb3955abd2bf989b463422300718ccc3527019796f2bba7deb42440c0e75bf727f86c2f50be60952310107b3b326fc5f952f16a663a51c59a3afc23186c2c5a2c33febcd165348d5d68d0122ed51fa97979b4bfb8ab784e111b2a335517bbfdc58c713db9cf4a261a13528df50f43d84bd1d1fd6b68fcfa3c243ce28ad208015792d203d54a842a7b3433a616d08dbd72c495d8c0c4eda1dc1731d11876c3f7657c3bfccd65d9b7f5a2dbbfe027aa58ac3e658902a257f7beaa3dc1cedfe2e623083b945c681b39b7027ee64dde115df45a4131848590dcc54062d0521656f02095c67122f05c3ef0b50a82edd90108cf14d3de7fe7c16fe0d66a5234a5b02fb0c233f25ff78cdbee49b587c0d97f5abe236f2354cf2daaddddaec698f6cfb0a51d89d95035e5e900ad7ae824adfc6c8e70ef152922c8dcccd0a2f7e45228d1f155699b3921a91c32e79ae469993f2962c3a24bcbbf5b9832b56a214d8e0fccb52e12639811468c69bb34c36bbeea232a6a89a951c5ff0df42148060d9772359a0f061a51798bcc4bbd62cf656e208c8f8133b393267b99a80bb9bdcd8ad660268f21d5de2fa4479d0d144503eb4d6fd707633e7b33ffdd04492fd273dbd3b0985e8ec7a18b13f055079d072b05d7e5f19f93e1cbe6540cacd2d0f59eb8d549098aa3671209fc007f3cbd9a182bcc6307773176d8da0e762155190aa9869d6811eb63fff50a8b7edc8308a76cfc2c70352832d87980077591ce0ae7e1803926774f6c83e2112cafac39fc24fd3b4f79c2294382d6875a82162d0ff1057527ca9ce26529d770a276b9e052fb0f2d14d57e52149960e01591ef45326cf32f8d20a9298899bbc564d9c50b3f6353273275c99d96dd83b03c70c57b5bdb55b897;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb835241b18dd6d12e0b43438ec738944c775a1211405886405b2593a5b3b9692215457326a289d1969657420806973c3da97552c257cb51a023116df6b996a9ceb496f5b9c360ba17d4bb57664bf124c4d9b6de1f803784cc7ebd141c5ae5a6c894a8ac5f63bb8a241de9c2a248dcb14cf78c4453f67fa382998bac666412df7f16abfbc7628346c806ed1180ac16751a73b63f596b1de18c5b6a16157701075ce6af73621d1a9941d66bdb1b1e21c7229913c87bd6f35a7716cbaff9fa4bb85b8bbd4156a8d77b48473f0ba6a525176a209de0f6b5ee333054f97cc1ec1364d0bba2ff32fa2b035016dea0270bcde2def885970b322857004f68bdc2c08750300a6238236c5bcded3a705e58d4e62d6921a8111d2135eff2b6dbe9e8ad9c4812ef19c8b3767ac6b409541c1e14c8bedd2d84de0a96c9589d083c5b7cc27c059dc978a5eb6e7cbb2d365e934409a75b471ebb84df3bb099ab47bcda5191c5a1494a3eeb0957c216cc472f60e72716a81e72edf76883f288c487f9220af022a5faa14a842a701f10922f067eee2411d283d490c5c1199eac60c2d62f43b0b3cc16b0078daf5a77be66051ac2d6d73358c6272b991f0870b8b0cb889f43925f852f4ab343cd10fd92ba9b61d1c40700f5e6e0ce9e688df8c2276557d94dd327c136bbc861703443169338d9778d876015c2f60ab4a3dfdc9e760df90ced5033db9eb716f79c38c25b8b2060e6e250c9586c82c58a9048fba076b65b1bf55f7690b5a49af107c8f7a9355516f019463c5ef1c241e142bdd5db1f8f45942869d71773ac3dffe619880568985a4285c9efb5e22b05957b537cc887e16918735b7370f4013ba677e84d870b69695266b8578da9b82bef881a3d3258cee4e7ee208388e404ad9f15191c89c22b7062ba747143ebf2bc4006952722f7b69c52008dd56195c9219ab1ee4ccec5546f8ee51c7480b681ebed8016ef7cdfd8d51f38a5e3fcee2f5a0d2fa1716323873ee7d8cddf1613b492b004566f9c0dbf503d67bb62140e4ac8a4df2a1efa1130aaec434e770e4d815b8eb3105b2375ae8ddee9482775fd145bf32141000278b34a2a0e712fea9b6ece16500bc4a36f83af0d43ae8e10f58e6ccbcebfe19df114f86db94bfdbd6d72f8005453f42a067b64b0b30b8a06c6c4033bc09cfbfba7e8d08e3ff465e98f4a8f37ebb06e629f718c66362723c49967fedd87e4cbc485e316579b305baf60db7007bedf922635f361be3580a4b0d373ec944b1860b5faa439712d4aba2a80b7be5b167469bca477191ffbb85fd1d0bd251c00de3dd245ea2bdee788c422f85eb4b728489a6bd6a896cc8456217c1170390afd1872079ad619b0ed558582b1c53a518a48fcf0982dd562e4d18d66d6d67ae665bfe4e0f15f8c7aa9b77f69ee8ada26a898c1d6b3f5b8d3194e51106171104ee3becf8384e7815aba8b5f2578e04ec228536757e1ed9fa9f856695afbefd54a63ab36294f0dab48d6a73d2b54c1232359d2f4648fba97237c6e659a97db24e50b87f081c0410d3aa5b5f017c20bc8a37336f781b09fe246cb50e6f4976f047152d6a01fe20bc54674cf026795a0f6036cc3033682e03993a5662ec38301aae5ff13d155189ffb2f740f0a8c34f1dae46ada1e98a3df16a2cb5803b290b0b64049e36626581e2f0486623c35564f00f04573f064e786b6ebc7572654a6bdffc7ee82955fb02a1b801c748c479d357799c3b2185fa45fb80be29de37a15dbf7c84adbb04d83768a843ef11a74ca33bdecc45d2f6d35a4bc08fc00fdc2f706750afea7dd77278d0bfc246f8daaf62a851c8fc4b93eafb9ca4d4c94468452f162a6daf1825a6453b234276fba761f925974b57abb711cea65728d5f800e4c3f816e1214d365acef45b5a585f349c9bb33d586219dab211248e9b08f613cef9636a29d05888cc3ddb645c3bcd82b8eecdb94cbf6e0fcf518d21c8094de1fb5e7103cb558e366fa3c469d79fdba5e8a015c51e85f22d5f482ba4269d7f3573bc3fbd90d62b7c7588635acb068d03b97d88106b6ed1a19c6438c93150b4777076bc40d5d735e09d846f68806208604a0dd5bb768501ab8b2f26761a6c68e80a4d11e984d5aba11e071b94316d627d50adfa1c6b465d6dd73a4c00895a5ecda08b53c715d286c26990bc301072c0053caa8d31cdada4eae2cd1897df9fe75803579bb6500bb73490ad835869600304a7bac84abdc692508bd2e5b84560de116fdbaaed85b1f396fe147b6cc161bf5aaca9c6aec81999e432584eb287025eea42e01791b18271881b47707ef37e45b23b3c1f10f002a3129a8c36b545f971e4d329995fb27400d3ccf861cc4cd2d04bb664b2674bd53cbc6722a255d04e17dda11fac6a5a88a1e708f631cdc0563befd850b7c23c46a7455c8abfe4324d4ad32f83f73c2280ca0ce8c797cc6d5a3779f09d3d35debba28fbf19491896af1726e794ad3480d9954d685f0c7e251ea90b8f585e4dfe049fe2584efe128a29d14bab590ee24f5075dc5bd5a0e346b50f69278bcdf7bb882ee475188437d56c00580b6e2570315ca4593e25f6de754db9ba6c68c0b9cf2ebf7210b975a0b6ba66bd0a4c290014c2ce62841c6fee2c81549e052d47ac1e218abe3da0d65b2a54572b073d8b51a7a6c6d42e3e26f48d944e8a059ef67c384df27a3a22c2ef29c7b86703d72c419a5849b1bba5663d02c122502f919f0d187ae4a23fb7cf50897ed13414d133b8fc310d201ff0703a68cf86e52f5e5aaf990f8fc791e09e191cc0a02973c69acb3a5bc32c450eb2a9ef6e559e79c5f04aaaf9edf11f6c2c40917b2a0ac4e549a45fe3d53b42f2ecc7d65655011fc3df1a51a46ead2293635121b39ed441;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hba297674bbad2fa248f4adc3e6896af0bd1ab83fe2c6efcbab17df44e6af9041ca150907283243578c02a0c0d6e399837023cf7417ea19421c9ac651c72acd54da25688d4d4d4a616b36e42330199ab08ceee8e8fb7f78bdc2c391bc86fed00caff7c06c293f8562abde449c8befbbcb888afe20815bcb41e7ab3959b30bf3b482fc8d8cbe33b659e810c15b43a39f4f329727b6c2df3defeabae79afe8012d29a4e27ee664ffddac62d5006305846b6384cddf7259693bca9922bf2b5e8d66221f55a2c7117104c041dc61f97b7ddd95153221db00b2adaf8f807c6fe44665845f2c42b726a4abf404e12d4f5dae104edb6e749d97ba6c18158850daf39b10e8f5915737f5e090b728a0de1d4dfbdd76c48b0dbbb5b1e076809cf982f2ea19478a585ba8bba3c7c14411e4583d12e82a352002bde342d23b90d3750699779b3ce4313102e6213f62bd376ca3c171e79f624cd47e231dc9bd7044a0b45574853b9dc22eba3d24be81ed46232c0e2250690f95ba670fa3d4686186737a34909712810c3ae2c5e963709682512f2b5fbad722496ebf94daf7423c884c307a6ab6b84a606c8b78214542ea0383c0adb5d5dc99da27c30f183d25a4eb91c6c4baa1e59d0c0ede22083c74490f96e68fd06d0f52c9321e49f1dc5ad37f73410ebdab97aff5d1d477a244586caaf28a55229a726d70d66d7952113c3491c132042e78714adc83e2ea821b8c2bafb8fa4e49265268a0b54ca07a19d7abe33d7b18ec5cb2615e71de6c7fef1b6a17bacae913f6c233cdf8dc154d79cd41b9ec2a4bddcf4e5f34f2fea335305791356b8498a8e6d69e39a9b8ff02327c77b950275e1c20df4f8224713b3285b76709f28980d631fc5915f89cff8eca59e45d3d5db4b689afcab27f7676b2dccef74d7b605ef4d829cbc4a8c44f1fa140555610e1265557b03b419dc602d62ebff3546070ab99b39e65f51ceb9454137b7ced1789cfbd54f11482ef9c0fca8ff84d9c2302ebc6e93e79ac61292e9b82b0578f73bb2e3b5cadbfff5619468175b2b3e1dc250c613e0577cebf7e0312c4b969f5a629ce2aa10ec53d0c1bc23fcd47ad7c943acc8e73b897a2c5d9d74a343ae3ed5ab639d2bb032e34c6a739009652934b1329c291c5a9ad9bd43339187ccc779bb692f5828b9c6a8cb9c1c30cf4388c22c3b78d9ed8141b24dd847f1f26232788e64e461dc602be8d22d945d7751a2280c5fae8a4f7b5fed9a25eef1e21ba22e67266c0b840d443b3b21a93c1e36d4e4ebbae423101b85cc2abeedf190c0452339e734c228f87db4973631a76cd384e8afd37837b5cf7c6c062fe4cac88e397dd6b8243486354849654ac17685e30dd838a425cc8f4b45fd05385428dd3fc51c0cd50304c3a50f6dcfd2eabf86721485b549ec2e5ca981130cd2953f222c24939b859dbaa64f6528caaf4ca67a54f52bcd569ec3c4fcccc6e3c5a017bf348cd639c344fa1c00ff3678e9109ead2e818aacb2db30a57902c1b40161de940b2006750983527af8728fceee5e6a8b497c0fb9b47f96df1f071a0cc99de2dc517179361654f385b68643e07f81af9cf6f4bcb9527e9f8ec48aca0249047bd0176a1003553acae989ba460cb3259aeb921443819b79b1bb817b78a7a7e41c08facbacf6d9b6d94e0f88d73b0615d13687d20beed12d0f628531559118c17e2b39b33e7e349ba38fdd31f0fd7cca54d571c9ed465fca0022aac571e884839434e32ad0a4d043184c3714862e89efaac286140f5d49890f7d3245b148ea243c008a360294675ace886f85a4366463c1206feb2feb5f68bd163f0df70db50fe4ccae93d06d50606a49d8a666f85abe3c04dd11aff29d6ea6dd937a81f57755e326462b268546e0b80c0f5091a8583b586552123f89048b172e827ee6ebb199d7acba9cf365ccf148f93004855bcb8d63755635b4b623cb3f99bcce2247a49f2918832b14f01836fa98874457ffac0f2e9a0e53437d4832b9620ef522c51f5a5dbb88cca306785ac80ca63c3b02a5d3a91cddbb393cf3c3d0b4298fb43bb17eeffee02557d8acb5cdae5b870f1eebec776cb9b7e652ef880859abba14f0d395dba59fbbb30c0bd8ca988b3a4b2bbd5cb449a9de293b6f6f21472cd2d57ff9789f9016a75d039e7b3a38be06fcc7f9ee4f6646d0836f60f7df434d0a8e06bde230b1794208efbae562c1653521f03c552f301c9a7afd1c1a9f285fac727079547749c3e7285946d58cb657a92c2ecfd7747f4c70eaf779ef0a21fd2cd8526fe3ff6bdc01fa610467fd0e4f30d6d11ba46b94b614e490f39d84d71ebb2ff2a796cd65144be29a942ba64590a128116ac97c9fcf82d5641dce8f49a58b4dc8842f3ffa74c175c2a5aebf24f17f1f7c85d488c8ab25fc6678b88ed6113f1fa4641c8684223103cd4b16f65d8d160b60ee0a1473b34dffdf4aa8281e725b13f4d4da816639f8fc623e998756ae3f3438d204e12aba224dd2de96589c9830e87676318485290a93ac0430f119e4534b05da0c490df7101256b6ead0229b28bc401b284de25fd70076def0c51a4ff1a9d31afb45f6a457f3dc2e2b78f36c60a7f9e3b2d5342428da1e508e5bc7b75cc9c522bec9fea35c99585ddaef93f6bdd0031efab5ba94618acedc89d18a6974b7c4de6a70b543ecb003d0e4d1272b081eeb855c576bf293536f0050d4900a563d9761b845db7432f0588938ce4d402866f2c349bc45078c6d7eff3b0f3e3a11399f1b2ed138cae0af35f9f2c4c4f5b2016d48a40868b239484add39812deae0605229cc6630dba066dc153eefde7b2d3d428e33a1ddb62ec25567b18ed3fa7c2e5cadf5eb164c6271a8137dcb8891c7259b609f3bcaa1834ec287d9141a33;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6d1c1dc209699d3fc8bd96f868731b67bd0032a57dc70916c12764a1b1fc206608ace4b3df42597fea288178ea03bade7a3ea75be28289b3e6ba0b800424d853777b2440a7c63b3578fe9c559bb24774e24473b4e0b44c37e9bc184bbed031f5766de43fa543fe647ade664a3c52d498c80fbfc77486359ac51a7b5b8f8b53331ed9a25452be2ad396f0764d3f81934b05c5146eb048c1827cdeedbdc3f5db6178c49365c2d28b2d62e677bda0cb8c2ea40ab6bb4d8237fe3000d3d017daea6948e8f1f04b54c210e51dc831dc8cf388c8e88423bac99e71c23ef2ea5c65b52dba90c4651786082757fd26c409385e7b2e1e880d46523627e35432383ed380f5d977beaa40c6f0e0113390ec9e13388a288fe76378ff5b15966b6c83c3c10e93514628049a2f4da03c28e76d3cba5a35665483f26d343a74fcc8856c893906ee18239c00ad5a0e9ac2430843d9a281fc50d2b97ff7b905f4a21844586695b6404aa1b129898598facab8dce154c6bada58fa5b9c2863b8aa2a2d358e4d768b25d87b86c6d2889ff2eb2cb4573b00af526417a3ccba60f54ebd148f9869a9f6c76663deb422937be8880cbdb7c07a23837f59d5184c3f0d6b5ecd774df1c2b2e735372e785e7450b24f2e064b5739ceff595fcad5855cb7d68aaff189fcb3f06ed484e1531429879588f80d038ff509e06c6cdafbce784146d1632772b167aa0fc4f67897f5a0ed5a494f210f7e61bde1d746ac76618b0af4983eb79d307308c995bb47a623d1082b0b340d90fcc91594ded0485dc62ac60fdb7efbb7e624cac15df3b189588b932b2a713e51916afc9c5c3cfaa9881930d5b02fe873be729a7f5843c3ac1a03f947d01a1215815ad895ffba4937e3b7edf19c69c7471acd1bfea380636bc2ef36d33a2831c7e26e643a76ed47bbadaeabe0a64bfffb3030c1901b75d40c370146448496ba2f3e10df0713aa9ae5d435091c02b11b4524fe3ab8f2e4c078414cdaecdad207a5892ae0bedbabe1c3ad22919637de145300c494722341f185dcde342a23438c620329f54a19b804110eccb7dace3188df9866d461616781350b70a9281ed7dfc62eb312b76616d354b779c9698c0e53bab9aba6e80a75faed188ac101168b2b8ae1bea751210ee26215aee996387afa4b903097d7c7c9c920117362d4026a782100b8b9213a65f3701ce0421709a96c5d649c2f35791812d020600ccd38810d3dc4ca704394468104e144de9090c867fb4b71fc561a8def188c877728b065eadf2bf01a7ebc7afcb4cfde2d657f1032d871a5b06042d29164c04cfe072cd4789405993582c6e5b097a6bf5b0cd8cd3d29471a1e9686505977c0a241e64a04a96955f5aac3083022c346871001bb3f8b97b6bb6b5b03e97c4eda9bfd303b769c12522b72db1406cee122daa3071816bb60014e2795c669760ca9fc5b43a1aeae57434711d1e6b4a9fca4c5f52998bd9b4931e38019547e97487c70e06ef5f617051eec6d816992e64e1a1bcf370a6ae854df2fc4287191df74ea649e36a4d7088e3a64d338aa6b457b7f78a2cf4b639cb142a73d0ca788231d9a854f9c10271ba9be7e41b3a3d4f542f4396eed3b0cd786f6e672568ad659442f625410042a60785f42e1a28a17072c51f59d484ce0a51f7a05968b91bc1edb84216aebcdbbc70515d37b53f8b0c53ee112546c269675deadcd0e9b906487c19c44ea5b4de75973894883b1d1811f38c7f5a98454a9eb1956742ead99608d4f0fe89dac80d51d16bd922fbe25818ad9cd2549ef1f2ee2a0ab1f471abfe681aa0e4eac2c0c0bc3a7fc804763b07def386b9031aaed7bcf2bce337bc9c4c68bb53e62ec9f751465a7f40387d10b080a7b86afc7b4fd924113fe60f27c9ece1ffb26fb0f66b7e1067cff04a72b8882cb4821e8a12d392c264fa5779a5e589b70ee67629e5cdccb95e7126198346ff0fb87fd546085a1554bdca612b75042b9c7171b525464fe8fac2b461bad9fb80320e770e01581f007a9270c4326975fd69f36a391029589486fdd49430ad1196a3e37b137301d20863ce0d0ba8bf36342614d40086ea13ffcd28fdb3a512b4c716b8cb2fc28c0c6bea0977d140fedd85651298dc1b272375acaa4ae481b9ccab1867498106a8562afd4ace2e13c09bc22fe8e6d92f868f5857b12368eede543dd328961512a36429516ad9727a152243e0030831d91e928f4073c75cb4a87dea894ebc2f9c7ca1fd7d931d956026d7a1d47aefeaffdb6c7638a9b805d5137b7cdf81122a6f56063fd43382ad5ca50a6f318d444c3fd2186e7f04455eb82b686190a4e6f69aa789532c0bc6b5bc1403ea87ea0133fd533821286cf3004a0d0ab1e38e99280111ab8983dcfb76681535739f1ec682727153f288ccbcc3e854dceaf13f9a3727b209e474850484491dc2daf346eb9c11766ca9211b4db940e4dcd1cfae89836e13939372ecd52e0b1d2122716e7fc7f3305779eecd7f944aa5cacbd779beef5d5c8c105e550a3c39f5706eb88e670402abbe4d2d6e884421be5c85c8107649dc996f7e8acf3fc38bfe8c28699d030448e40348d758d900f38abaa0f0bef63f4fea97a6655b3c1c36830a5def2ade64d019f6c9cfb932c52ce902e6b5c8875b15d9854766248a1a00d2212f19a4c9041c8a3d87516ee413ca253e4f8faa2af1ea25470a8c3a0f218867136a0247eec544a171adda51cd0c912517da53288f334b82cc0ddf3e5d190de3e346471dce75f2b530819831adb463c351e9ba3c89102f56f769d79df2532bf1de4a067eb0e1b1deea1de30cc0bbab1d3557dbec8d24fb2c277f43bf6c32777c163e6e37c4ee19a5ef427dc5f402dfc211c04ea2b87174896cfab6fe421bc0dd0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h50a0884e480cb0b9a7a098a7df7404e96fa568e8ea202584e14ec9496a37cd3d08f8e1723591294975e3a8ced49fd2008f72f517297622e0805c3779a9d21f0902207a5cbb995e9fdaf6c047da0a4785f6957104ffc148c2e17063e54a1263b2efeb08e6464f88d8fb33b6a34c6a78456780d51becb8e759d1ca294253d9f9e59be7eb5becc5174b33a9259fd0a99f47758686f33f784f75ea42c271baf530f48bbd68d5b92361e6b408dbc8c328cf1789715625597774a2696bbb0d799d7d572ccefbd8386d6fd527703d6db49934a56936103867fd553af4da6d984ac68d7129de204daccadf249c83f093b1beaa77534846cce68faa29a9e15b0f2722ac029886d200f674fe0471fe6d7b545f342e55f3c659f0a77489c031527adf043a37ee39d7e4258ea6800dbba663c50d8c4c9dbaf5bc06f6846e522ae1a9bafe08bd04ee147810d9d3cdcaf7d654c41ecc55c8def8b642101f3becb3e2a86c2ee4ae562929ca7728381f2c7320b2d19c414acf2bcf25007c7415740fa65c1894df3ddee8b5f17d928b944fcfee0cb2ac4aca5bda9bd2811428236ddb63136a5ad9859864d8349092dc5c89c8744d2ba5ce5e5193b9741194f3761a8a8f027cf28caf32a8164b9d42f697de20f5decad0678acca3aafa07823506c72adf533b56b1072cb81e4e0296fbc2bb42943756f217c1951f3c3a4f1e393c25494051f4a703e44a50c13635a547764014588163c2312ef21e7acdae84badc409416a4b0f48c034457cd594fb67c3a426ef8f4650f8c17ef09a98e0724702fd3f18fbeaeadea26cc5df1c1d7715dc67c1c26bf401daa09b15282d1f7ae441dcf776bca8f8c7a0787bdb22d40ce54e3a287cebb19189ec1c78430ec3e096dcc491fcb0dc15100f8816d957c0c04133f0fe042f7b35f55f09d225f3704452c3b1ccf30cf0eb7f2eb100c17b0880b2e20d4ca2362fbd02a0037e486de8919511e811e4f9ecf37eb58384569a85bfe4e47f67ff8920344b77aab5726c84817defe232bb99621bbb7b0821be40c6fc99ea164459c216b777f51b914af1d822e8a4c75e7e46f3e3f4e59d56f481f741d95fa293f2f5514fb5963bab32d904ff89fb28934fda2743a1ee7b40c023943d3e75827b1e5df19f396c25625d50a2a3da19d11a3ec8fef9311607fc581e43f16bc82393380635563174b846c5f87a5aa67e8107c1ed90394d8376d779d5d23055db036d1a16cd0661f71a113f92baa8c47f977e845e145e59b946acc8f289b0bb41d92cb991fffe8fc0a69b62799dc5a1705af7aa0ee1804e148ed590ea7dda59c1a177089834ff92867688a4bcea6f875a348a7558ec79f408d2e6d6e1931c37df265137e36c2d978b42afc880bae050d0bd545c1299c87c97b6d05d1350e7f3cec82dc324fc2694e2dc640a0aa51c0ed0c63571bf28c9814a736a8b7d2bbf14836102c2815edcaf326764bfe267414aed3a045d8242cf0bbc0922c3cb5e51275702103970d25f1271118a1fcf26a8e20bd15fe2be94eaac625be9c71b81e459a8e48ab4d0cd5bfbb18e354245d3af1097f59df3509b98143533ed2ede0abfb265fe2ede7cc1b6baf213e0bb3aea03a6f5ca653d1021b89a52e1286950c874dda704b3fee8c1e069ad8b14b9781408f2aa3d11862017b0cc8306e339425c791383ca80606515fb81f8ba932da436c0d5d591ac461a536071d8a14f9f64f7004bf7447e80594c80e5cd8a6a9393b7af4374e945e3185353e6d6ae08a0969a63598b75078d4978e9ea9938bf4c54ed93d6fc346b0f764ba38a85d4e526ce0cd7a259f94c3507e04ab6cab17b4f685eb005ab7656a6d2f822416a54808d41940597662955000ee80cdc704fb4ff83a4330c3498ce3c70cae16a5aae3b58c0e79342e097a1a25fd664460b71d19f3bf25031c690618d0242eb8420500d6ff1765043f88fdb5b5dc5e926850502321770603bd3379bf5726189e485718847a455360081f12232742234a4f87168670920c4954b154248457acae84c4c2d3c26e549dc57016967231bde9ec65135e78b19e9211f7fd2ef13dce9ed18d48854a069b5e864ea5a0be08f1f1d8da4699f879a54d647d8f46a1d06257cf658ac845dc37a30841f0c6fe75e9fd6a125ee223cd929632ff0b8a936e30338858846656cb4ea995afeaa85a5742d360d25f2ce731faf2ab68b85127f586e48fa5bee594a6e2f2aa78b507da991bf78031d87dc9954500277ca9dafffa5f055680e99c14e827070fb6fe69f9339a4d363ee98292ee28d93eb2c9b064df45425550c6bd9a7b1f1bfd6ffeaa773f4c04438801c05b263a5a6cc129e3874456e766681de5730df5b5856f90644fec46f6f518c5ba7285da4a609051684f1e36cf81a7be44bc61aff826456f51ed15b3592f604971eb553f25f3f7934f5e61dae218428bc9d3b03163f60395d9f68ada067b9fe773883d864f66fb138f74fc84fd530b638a37118197a2e072c069ca8fa3e977d6ef43201ac10b19dba60bc9dbdcecb17af2e99cb141b5a50ad1089f2118e87747651f3876303b2b96ea477047075f2496a255ce4c23039734c18cb02a40bcd29d908b766e2f2845aa95fef21bf48f448e6f5452b69d10a28de6eb9ee36a8232b3aa50a1994b6a24f9f8f8e9f6adc00cd1b1ce81bccf6f9abd2324b5953d040e3d085e97a240dfdd0942dc31cd45e9014e90f073396353c17b0c3d09ebb63cf14ba14dc53aac0d164f3d1744731f770d117361d35339d26508a38c3da7d2d6c2e8246a577b8826cd146ec84a1ac5036f9ae2d6fadc9fecf905ddb2125d362632556cdc2bd7fb93ffb4a57f66035bc8048b84e36004bbc8d006cb9160acf7c8f910ef5f03311c1b98adfa9eef35f04293;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd9b722e9e0572dcd501b8ef4531583e4993f6dd703efff5b534bb90d2ff7f24ab53d05dc3283584adc5e8a9e9e79c9d76b659e0845ffc3ebb24e6bb75965b58c29d1e9bc71ea4632f24af4c5c89eda055691e1d5515911df018ca2a90b1c8c751afd6424b3f380262fa55bb7e07b9fc03c3a4772e62f711c651461a829ce2f95b32934aff9d2cd25763e2148e7f0082ff4fdf1cfb39d926f1a05c1e699ba34101d1eeaaf6f8edb3727a69076155bb16b9e4c6347a16599bb406ae989b8bd498d52f8e1731fb5dfaa1daf92b14641a0c1212db15f975d077d4c64e767b086f8310140c39c80ef1e58fd6a569c33ecda7a2de6e98551251680cdee4a84e5c177cde6b255ac05f13bdf8eebfceddff6e9b703b166995eb6b84921cd766f95895cd33b7737d308406fc87989b2155e6775a931a680cd4263f7043d4e6bb7bdb486f97c1d39ae93eabfadc3cc2afbda777f00a6a2932af74241c39797c2c8796a2e962cd298a7c3b32e241fdafad657e25e9f1dd010d378666fb21ef7157ece1d46f241c9f080fb8d8d13e224d7f6cd3aadb88277cd69b44fe8c8391b098b8ad18e00601842a9fb8a951603f6b58e5f51908130176858574d4ec824a1b16f963e567fe7279e996c25d60c56a189b920ef239c5c61a175eee1f0208d7363108a0b820e2de8f897dc15a60cfdc119d6af23b57428add3ae34faec96690436fe88cd2367bec13a11a98e3be2f3dab651cad429ca55a419d6613dd5ab072273011483ecdff696968f048a060da2d5b5938f0f8144fcc666efb5eb3164102ac75541508774f4b00d962a7d3b047b53cec1458348b72b18e602e9ab51dd8eca5093bc989333d8c09db906f9f3e432f74ea7ad792d1e62fc179410588619712454d5486cdded51d1958538a94c7cbf403d9f0dc16b326ab65ada69ad219130b44eaca126e38268b4452b11e4975b00e819aaa59354513d87592fede6d25dc9e6aa87d086f8c8f4845289b0f22c2a386be8541742d8d90ee7c18d0173249f03dd7001594384e77c68d613619c385c1a7962dd223c8b5363fe0ffafca4a0842679f9b161a0234290a202b387f75d0eb7645dfe55b9daa5d659fe5f2364c2e5e84dfc17e751e7119ebd223ea5f5667e2f2d520e926eddb7f38eb97e56db78266363c6df6284a088017de8913191061d51773196313414d2270006569c80eaeefd878929a8642a3257d22229ff85b8753e767754e7b10a0ed46b40fb4440dd32c8de0e1e19e8003236c5e8b9f9e7936093366fd0fb982a24e9152730cbd3e1f2f2ebd099668271b218c0514b76b0bd73a25c083e0401ea9fd5829b385f50319a32a3a5ec17f6818597fc3e271cf51d18b44bd752df53c611fa84acce87ff6e19c897d9ff2d997d1b6639b0e026f62e87342c4b1e98f67ce1f0ddef746ebb27849d0ebecc397d3806ec1a1df4477b25430aa5a8e34ae77c8290f020aefa02dcf77caf3dec4cd41caa2d7520e5085f86bf50e81f4dcfdfb99f4a7083492a59f262674f8b1b55451b2f350fd1bafc40cc6a2ff061e788c3b605e62a5fc8685674ca59966fb5a98ad7039b1f89adbec9df7da1df011bbc29f54b2a81d876ca6fa450fe0bafc255b8f752fcb0ab5a0e33aa9e90d0179595c808592482abce4d0630aed7d47796025d86062057df2a7467d42e7ee971ba7a1dd8d90bf515e4472e9a94b3272a712e06290bc5a5057961585a4e6dc733e6bf1d6ef46c76255d21ae04d2800f3f800b28684e32926609ddf1e63e6f2d5a94aaac31c6f90e1c64bf89ecb1d0765e348810d7b23f191d689845ecba3c4825470df3831988bd8688e2babb9ca9ba7b45b78d6ce1583a9c8e5c400a69b8deabbd3526a8c722d2960c351e6c3883baff29636fb912eebc1729ba68718d76e1ec5319a8eea91f14d51da58fbc33b780528c18140eb2b579da1889a76b4aa091647480e68f92f60eda83cce3e32fcd7dc0ec72ee514c2c4431d1fedca80753c5c42288de80f9ad7ffe2d62fbe06671bafa9b1dff0e06769334bfa4753acb11e4a7d2d89228c7c570cd8d3fefb7d47f8de3b2aaf924827d96e7f2a697c4ae98be3b7da517a84303d91124c5fa3c7c100c160d529102ffa73195b7372fac5c02758d464427ccb0743c5a51851378b0c3d60bbd88cf1fb10f9866b40e8c82bf0069356fcd8ff23671831995359cd87ef881de9e7df5e23ed938906d92cfdd9fa7955af6888751980b66a1d63b554996822a182b137f358a15bde732703ea85aa08d7b669e4a6ec660b83e23f007874b1f40919ee361334bdb6e85c78dd710a988552895d7466214b296efa0e72bbd5ee9612833eff86ae227fe7f6b05d7bcc507d59d6a3d84b5458ea3c192c5b4f3b14fec540aaa469ff892ee3833ffaf00aef45ea06db3c7f17d241bb504f07e0efc50008c46e6b7a07155ae2b4e96091e691988eeef63799bc7e9759c72cffff9867fd0f9c7a8993f04a21fea8e0b9d276048c867de01aa3ddfa7dfbf43cf0050668517a9291d3c72a3d6533588dc662ae14b1cd73d6d4c4fc5ef09c0bf99c56ed8080a6c50cab9a5c49586305166926d1ead490921bc9cb710636d9b4f5fae49e9006765f794442e9658e94b7f19360a1286c670d8839fda8f2db7369af79446bf603ae1103ce0cefac875ab83612bf87bc91e9f56b97bf7b7b11fc018a18bf4d0b71aedf0912c1ad7fc2f5ee659c0469573f13ef905838ba628a3e03246bc3c8d946e559d3044021faa7e83f8d07b9d449d321cc64fd8b5cc3a2f9b0f555ca275e194af605c18e3c3d2d51307c32fbe80feea24857ac364bb2ca494497057fea1c3ff2dcd957d6a7bb0b3fffe4d5cd64547d1e90e5ce70b103fa836b93c536ff01eec58b129acaf3c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h115135b1a7f447737d52d320553be64c772eb6a3ac9cdfcd86680b9020b3ee4e0f555f2867cccc533f14f2887bc14e820af6b7665436a708d96bda825d3b66a5a84a7a016ca0a9e5f5ac71bf3d54ae45837a914905fb6d858f9341af14fa5b53e89d6f44dea6d8b566910c852307054a8a188b983301aea4a26762cb9bf8b09b1159d510f8a2c1f1d450ebf29e7f1944d2d36861f85e457f9fce988f097c92d4eaf28824228f3a7d548ba55d42e38ba167bd6ebcbed5bc2386a256129e9d370f170b33c4ff6cf2ad22f0992c05ad5283a834b8e434775e61907695e2a8e6e918ada2f2e772ffc080757cc70e3f0c867096879621d758f2c692dda27a5134e699369c5efd9d53d7c5c2dc0c280cc3f6d72ae27c3e594d08f70fe0a2cf82624f77322a749d83a10f11561d8ebbba1f13fa309c268083e9a0a628e2284eb050325dfee84342524e05074df0553d15d09e8b34010feb7e9b539d0de04b95ae5cdd674eb8c04ca66a66bc74b88331a76073839a0012a8d46a2ea247e86ac7ce5e21a3ca1ba56de3524f17450ba082303a6834f84c86c2740135043a8048d057746e323a9a12f154d97e34f83697676c27da4a44a506bd7279c5436731d8b8244a753e9255c4b905add315888aa34ff391b796123caf1890552cf634dae9d3d26d6675d17dd801b1e37019cdc5f2c9a0cabe627f204ca2af17bdae34f34fffc2f843bdf97fb0567e6bc64273ceca6412a4e2de7dc056bee5b074cf7f3ea13cbd7c96dd5485ab288212713b27369c2e0555707336d8656e1f782c99cd8cd84fb0c2e2b3cdf4f113cdcf734b816109a8e65de89089f875b5e26bdfe948f4e0a55f86351c9034365eb91176dcd19e072976f51f6bd60f7c2710dd183548d281438d508ab2115c31f3bcb2696ee63f8d5c73c59edfd0d8c69041b9136d4397f68d9c938a0e265d82a4cffb83c01b25afdeb07c91641c199b17bbb309a0841d237634d2ec1669241e30f7a9f8aa1fcefe8d403315e50881027d87601bd3c0ba57be0043f553b829afae826c8e8c80d61d764860c4d594f8ff169b917a68c02fa0f54f8aa1b2b0044032ffafd9ace967aeecb320dcd6328a7b1711f6eeb1fe1f152b6295431a7425fc6ea33b22e00f7176ac6395ed1e1f01d1e87f87f5f0a77cdd34d63d6f750e04e8eb083fee6cee1ec01dfb68b8e9fbe4db5e0c63899c084fb7bf53584e2959a8ea04d88a406bb6b15b21cdc27aa027a9da84a2488323b95d6809ed84e19fec31f4fedca1a9822a7e1109436dbf08a5bf0cfe3e29f97076a3928a91c1ab9025d1fcae36f6c0d79ea749955421cf0e27ff1ca6883ac0b711954cc543ecc812445986fc34cd6d5862e8641c9f64daa11360b829e85e0b516b23b3da419da8c70fd2bc6ddd3cb86edd23d607ea0efda9de325fffc5ff2194b33c90a49a037ea1b76ec78f335d44e318d228a7a7a6eac219df14386f6c9c72c2af9a3b021c48faa24e55d6f7b8b4b1122dc12634a722b575b8db1d122aecbaeb11ef9b74b8e63bdce0023c6d9a0d1b2b495604ac59c9fab1039212c5c7fff005351813e72725504fdc0a90b06a56c2b268f8697b8097630f90d91ffc9491d20f52cfe90b5e294b03377a7a9375086bd5b75e946da54350093a0508d4dab4e70efd3a753f5187bb2001ee708a72d6906e04cae67a1279248c1251db3e820c43ba438aae8755256dfa24e4a26e8595f1acbec8983bb42f68321498d636a173340508f12e5bb1493c9f0c8d341e095524a68a1ebb963882d26d56365b931512552510739f892198d2fc2bfdd2d3c837214b9ff8cb46c83ef26456eb91932b1fe37dd1ac8fd48f3b31422c34ee7574ff9677c49061fc265111327beacff58dea7048212b7acc37e6daa18b723906103f62716e0962c478e0ebd311006d14def8802eb4388df37a5ba522e8bad39d04bc040a1b44c171fc49a8d16f7437ff83098f219f44c0463c17338311a2c71bf8626fc5953c8ddf2ab774a263c613963479461dc370b784bcfae8dfc634e3c5f7d464a5ce23512cdea3e35775b711b931bc4b175c91bc6e968344eb4643ec9de41a4fc0c6c37b904b629b27e7bf06278dcb118e2b16f7638881e080ce6e01a8b4b420283ef3da4bdd8a9aa9445234c02eca1d7d0ab8d90dc519f4b400224a32fdd1f866133355a2224b60826b0d243edf4c320f7906b9e2c502592c753db35f464ba7a1532f82a08a2d92f90a6175740153d1badc9d264a55d5e7c8dec37afdbf273342535f75137942abe93cfee91c1b45c466350868a5fa24bd457a9a9c30c2704b466627a9b20ab23569bf5067acbcb39c0cd794d692934e8ccc2c857fde409ba9a90a9ee1cb833f89a9e344f2140df13041dce435b2c383b634a736e3b50f75e4fcfb51d6d387710a48cb5c32992f46c3c260d3e10b42169fdbd1538c1b612b9105c81980dce91d8645109c03c83a50780ce71c5ee12a4fdfc86c6fbd99326ada28c9c1588101cdea1167f2004e45f11727d9bb778cda14012f1780916f56bcd0c0df29a685ad183446a651dcb8aec9894d244cbfae4999c16f3133b7e73af4bd07f9a491719a964c595b961f9b02be5a753ec2593be8adb073aa8f0f5ae466132aa18ef8130d16280c4bd0c68a945c9d38c6cec1f1721ea983381ff936e793a397de0f08ab57b6ed625e4cebc45d94885ef2d6201c6ceaa376b022cf8958fcb773b18d2769e3d6a74467f8cb90eac6894d3c343bd9b5922f194551c83ba2e2ea51687c32263cfcbb5f8d74f40cc2a94c518ceb4392f04016a30f7dae8f27946de6d45d0eba7581d14d3bf5bc524eead69ae91cb9b31d2d389a11623803fae20280fac4f0f6fcadb6d09e7c7715d37807164855724e80095;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd1d43f9201c6d4b9cb70c556aac3b1e7c672e1babaddb7ee0d8f655255932c88e37e8ee5ba82c5e6007437625090a6ec43573d79de59086898768a1b61a7e6754ac28b7d7b96a540b610355e6e37595cc78e52823376805fcb7d17ac25fd2e5dd224f80db92eab29274ebae979526e7c1942b95eca115e5fa441ee9088180ca3ffff9c97348a79e6061124f492a1df9757da9de3184a1410a8613e0dc38ec1963d6fdff39069149653a2269c6fe6befc949f1b8d5c11ee36f0ee48808c51335ea04c58d66032024b50b83cd9a3491a763f5f07410f0b58d4bec9c926fd5a82e4cc0fa9cf7acba0a1975b9956bb1e82a1ff914d329d73206cdd31566ec2c409fe5cf6b822857e7cc0337c03e0b25efad73e1e05c0ac46cf2cdec401d372073a1b2117c83a5cf7556230bb36c17655c0bd51546d960aa178ec2ed9b36e6bc48236e7b0788c2c9c08f4b19cadcb383a841eadab1a9f5ac80fcb387a62c355857f78ccf513c260e5b33f800898401b822d5546c06a6b6b4728c27c9b3811e36a9aecfebc9b1d42f36f5b8fa797af58a59dc046fcaddd07e3bd75a90fe0ea3f25fc85d927233037a8c45d8081f6a4a20022e9e7a1079f1d7aa4dd8607b194e0075ae10dca180f060aaf066b2f0685b73353e2f6d91754f547fff56f320ce9f86f309ee0c25d13ab91d895b76b9b81a54547c4fb2a52f67a0b1b235a2cc225a665f83be2e0fddbd079c161531f7f58aaa0c074b6dbdf1dfde885254f8320c763a3dbf1935b0422a2b0a0109c772564f2b2d4f9a1d1dd42340d06db3aef1563e0418c0b0b3f7251ecf16b346023be53e1bd69de9bf554ee82b1b666c048fb4e32e123bb8ea4e46681f2f9c67c2d67abda431fbc1ec8adb9d489b87b4400df1576b8a88949a89a3d2768dc8961ff455adab91fa6cf1a6f6b3dc796a031013660195b02f7d8c849bb0d5ebfc2547ab317132752168f66fcfb84b3a2714eac66552ed146c3a77d70b2b3948b5bce892b2982c4e401fc7d6f8ab23ca145938ae792a3d8a0dce1f15b5d9e671e831c4c571db250e0b043e8d50d994759869a7235f6194760b12ba6497fc87b8979c3b11b8764b03b6ff2c6260fdb21d15738cf106fb9aa908a9d21f33bc38df3020820dbd8c030091957c1247c7d6dbb7cbc98766811132dbffa3f34554b2b2f9f8ecbfc2135a98c71f060cb712f73989f1c3e12c570aa321ff1bb1905b3e6efddf6b695d633a857b1fedde9dc7c478054d5f781246f24aa03144527c53e6447f24fc5a4dc1e30a1a029b4edc462b25ca7339257a91bc658155b2c1009fa8abd8f65ef6c19b82e87df2f7510c5d8fb202a52711a7ebce8cf123b640ed5ba40c98daa19e0e02aee1c6057b8ea9a1351c27ec9deb2611aa7ba75c828a87bcd3bf83a2ab1522a2e93a05e5bdcdf10425f391460815b0cd131a924146d9ac9fef43c3b08eb098c104a2bea2da39a91a73070667a326c3b2ca94cf9334ea459028b8b096c6a82948eaa2ed6f5dc1f2cb53d1ba09c9381ec06269bb91d276d2d008fe91c5ed5911fa25dab097e2da303c1db7ce52f2fb45de5c7a1014e58a158ee274c083bf37756c5d7c24361cec0c0c1aaa53ad90cfa2d8461af8f492db950d0dbc1b4420976bed8bf58e3150b121ddffe2523aa4ca7f9e122c14d098a71f04a06d2e8338459abb9ac076843f8040be8964e47c3d68ced60e06858d06b1de81e33ce4ce122566bd75a79f1c74cd19b53f977bad7e90891b3224958d4cb538b699855c69d34084b9a45d5bb2d10851625e35af87d41d834bf6eaa6bb814de7940b4a862f3acb9cd927436086d041af88a2f435fb4b2ab6f579a0a18a8caf04e49992c2b89f6f9653c84fe3c4ae69b50f997cc82e2ed3060cc9ec8e461a67badf6d5aebbecc4cd05482bdc05351dded42b3c4e7720261e5274835a178654544665b3d325fa6f1a695c16879695f527baf3c5a50d8f17d2bb562d5406098fbe5b392b9e472543fe6e980e67a5dba5ced141cf3b9abae063aeb9832ae76de4cb0d006cb0529fd44266bb33c079236bcc6abeb23f20310af3a7ff2219bd9d2148298a686c8879950d798565cda48ac6d5b1b70bf78baeea5bc3e88e124d0dc7746bd4229e8f34644aa75321a213ee2ec2fbc7305b86d1ec051434300ae3f79a99834ec9fd1d77743032007ab2eaa8deb7b50b9e1c6a83acb8905fd493b7cbce65b518a86cb8dd55318016c342faa4d5fb04a7410a926c255740489b2b2a975194c5092e6beb78db24bfc8f83cbb7bd2565688fd0ae8af3a9792f22fcc819d361dcfd3663a938ade9e9a929e1001c97979cebf828a54681ec4caa3cf8e0f524e3db0830bc17e92fc49c0cbbb8fd00794eb2e818a5f58d762f3e00fda15dc876873490c5cd8a920b5e979ca62e8e8fd60e24ef48b9065e937dc04c2c124c4b5616705834b2dbdbd89c16d08a11d2d08ca64f3809b8ce3a400c145f17e1ee7c9c51e01db9b0df1b870e2391e00c4b45458a802605ec2cff6050185e9c0057edb8955de1cd7571eb2ac919922e96665c180a7e5135d6121717950054cd9f4f6826cc3df31d74d540c3ee4c6c6120f16a07b8a819084821990e3c236490cc269d54663e2830345a13257a28ec82ae6e33399330e760955f49f8bcc5d876c8809d5c548577b77b1bfc42a8d798fc9f33d80936e8e6f434f0ef7381b5ca5b2b05ad022eb8d003c347cc3e5be48d731dc7413741f5502c5740e3dc698e9a2b8ddcd4807cad609c422b1d8f43a398bcaa413f5144d6fed34c8726e4dc81f249d4cbbf0bd46ca25baf9e5b7225521966ee9cab2c1975b3148bf822ad8d38b82a3c97f670f41cfbbf0dcc73092bf0146c47ad4b5c7ddee28df45e16f568dc099db55bb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h263af91ca93a82a66e0f01a181277f926a136ac4807a9dbc6279aeebfe02ae57f6aaaffcdb69c803c7fc129d2e1463d88bc9f6a26c4e1c36e057c4391f8df9a868ab89b59f9c6d07c1adea7b9cd966f19fae3a1188bbb6555388ae68f1ede55704376087275e9ca0a294eca55d5aa6c017a7bbd641f7981d10e293c907ec143514d40d7533f5eac8b8d688fc7f1d8c91231297b6cf7127495dd27df4210ba1e1cf64543cf4ccee5945e4ea34f4c697d6a186f8ac5b4bbe4f17d93e39c8a1d30defd045a3facbad7471b0598fd1406cd08a93f3445166aac7c9f916c881c63eb2f509ae455bdad712ad3e814d08ba979b2d3cb8ab210ed702bfdb9b7fe69534ec2f4c5c6cbdf0da7bf4ee026a28ea8e8e37223ee9fbbfd9af66eb2bb4f1721a541d5112b7b9bb6ce29776e48bd732608d96bd88576f08c7651c7341c1d4b0157eed877b0884d811039af9d6c8077a0c8cf828f049fb4bc31553e3479ab0d8ddf7400f33e04c691640c8f46e1028e63bea842aea4511ba4ef9d38a74685e3d216ec72ba198aa36f52bc42c9f51932fe9e0498b9b8c55be137d00f59b90493a1fbd127baacba6a0fd5214f606d1f19aaaf24fa1ed77bcb414fc9cec986d53898b41bfe71a560e3bdf66f54e8624f42164fa5bdbd5481907a773d5b8217c390f5ef2c55aa25052699527f042d83eddf2643aaea01e5320eb0121221c77def9b99dba3d059e7d0f5dbe6caaa6aa48f8ec0f7e70db1b610a3a9fd30b5edd2c4d0d56464e65762e51f62532e2c4fde006a6a2ef14e314c70f7cc98ee22e5bfad7732be3a64c2bcc27a3edd0cce4afdc82e9d88b9870d2de6a7b33a56f7c73ee67710ab0dd7911b6bec2f8ac3c7a82dd5776d9a6dce271c75bcda484beeb93390ef14c1279a8ec4ff3919361e0b4353b5ba51ffa202207827e26b9d5dc1db7488a39c63fa6ae65bea42d8cbd79848ddd2dc8c3498f998b5cfeb02cfa90c107687346ca4c9aea82ef7bd2522e559bfe44c9685ea01f61de25d01d6154df21012be2313b245746e9623356e794910ea90b37cceba769ae849601353b4ada31954c3d4e45467d40128abe92a76c1a5454d3c12e1b17884e0eb2b2f7f9b0e35928b5fc409ff7099856e00006bb60c2e0ed960a7aeef53aeb08f089a221b5ec66d75a869a1146991842fdf7964796a3984ae54ced1da50df2127356bdfd5e67d99f34421e10ab707ac23bb1905d91892a1459cf598a3665bd714a49608a6f803ca987868631ba4645075d3227b56a743f76c91a1bce17a006dcd0eee2842d9db10ef5e8d0009a7da7c11566f0d77193207d4d5f3d320221f570a6d9554f66576f6db703803b5d20dbbd193dca1d099220105339630b593de6c5c89ebde7ce9188e2dae14900ee9becf2eee9aaa43ce7f95d7435b049fcdfb4f21f698c73195815cecd81002303ef09f2c890e0d19b20d4ec17988a02c7daa92e528933cc03b0eac221ee68964c9e93d7a9dd6cc012c594b66a437f47942e79fafcaae7e3d3fc6e40e8d5b271f1cce94631785885550ad3517d9aff1aa295715080981b120eec987dcfa278ebe568a7a57a5258c27f37a38b831e14d4dbe948a4ef7d68cadc8092ee9b58b1d68c646078f6589285bc31ee609556e8d033b948d56776c4225f73ea73587a9b744bafd982ee35774710d73625a02a2022d33c3501148d8e3be5e1cfb53fe25569a3f1138ff17d45b3fe6ce4d14027e1cdeddfd38cb1965044e0ae2357e07ba23dde33d4059a57e8b30e721d5b4987ef9836032e62e1e29f673ae430b16fa93cf9e8dcb50470d3538d9839fac34cdbab0ed6accee9e1a0c53786d5251388bd380da9d08943349dedbf22607bac8c9a0327f91562ebf8f36c000bb547461e71048a235b2e7477e9ea56d9698eee6b81a8fba935662c9d3859110b9ac6b6ff800051689936dd692b72255a63099fff6610d664bdbe6de938330c8aff99913f451813c54c633be984a097fdfddec7e0e1d0c3f0e68e29451d8a53cc4ae93531c6331f212f365c742b2a22c217ed8b2bc1f0c5090932d86dcbe686d0a11be6f306d09d8868e37914f39362a6d8befc11211de28e1986a1a4961bd74398eabe480565c889fe7fa8118221dc05948372196a9508d640e2300d94980969d86ea23c709ba2d7cc880fa2d459ac78460edc9ad8eef2334cbb28fa062b75e72005984d4918f6194b5510c6be19518dbf2a69f2cfeec5a5486867945ff1eca7b56b1ee11415aca34d31614870f85fff3937c67851801acb7ead91fa58734c73d9cdc0c8a1784fbd7fe9cccf80e63dfc077b3e187b0afc447c64e99a81b02524b2f847d74e34f75537b942a8897f43ec58d57e91c10d6795306571a82f0064b6a7b59651a7151ab5620e1714bc508a1a0d3a9642eaa15d1249a42a8949aea5109b94855ea6a5aca9926743188f1f496466cbe092731617854bbd46446da71c54afcc488ad1452e4de03509bf6177d2031c3b1781984c5e9ea6aa2a2091f86253ab8e3d6584f86097519844d68ec5b68dff94cf4dfa5db8f64e2d52009bd2d899e98fafbc63c64f735c1c6e55a46bad8a01f5e1c69bf7122512ebd1655be9f41ff14eccfa9b3ef0ed269a3c1c6e6b261cefea64f0d5a5257930e5ffc421d63bfbded80eb87e2db66c09cc5e0899fbc5932404fc0961c3af6e218215b5a0a9ecd325be259b15b563df831566ecdf242159f777c291ea88005351731accd94e1d819ce820560666d5ef9a9623d4a0a628fba9475ae3c862c669167f2a28553cb804ae32bd8d4426ae34d633334b45589b54d8e78248564e01ef5d21d63c8f38ce3c65c8dbf84da8298198b3765e26b2b44d48830a14a00fe7adda456790850208415b2ed45c3250d14a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hac25e3f4498ceb0b69dd5abf5834bfea0616849af94f8df463f5f9ce603e9859175496f94ffdd90825e83a338eaf3a1d0cf7b9ba94ec2c613eb915fe0fe4027b0d1b545ab0ecfbb1c25bae95cfb875e509a670beca206e97bd12a55f17e242613ea15696b62df9c8d48d33a665da233850ea0184f408afcf823f26ad7e70ea1aca3c001120b0bcb74f7d6fc6f1d70f8eeeca13a43274021e3c2c780b93f90aa5e152366253fc10cb20ea1c349e45c48061d5b16e2f2ca4cde914a733c1c12144df4deabd5da139fe4862c95bcf6519454a9f1259e057baf8a9bdaa56f110d0b3c0f1a0ef45a9db76f2982b84a8bbebe9ec7b3e45cddcb495ece4216c8587b508f95a37f8b9ecea13a7f7059cd852908e6ca4cc16859cff6505e066e3b9cd75d9b96ef56d4439ea95e32b3192b0c8c1ccabf6f154e208c94c109f51b22f7fc90caaf0e33ebfe908686ad06f9ea5e0ce0e87f2e613b1decf4ee5595368d30a967937ddf328b1202cc51b7dc78fc08539e14c42200632182cee754d4a69527af98bb6d5c250ae6700b0496d058c81cfe4faad0e07366d98da517c4354be07a8cd461db3acbfadab903418bd49178f178c2407e872ea9530ae1cb246549e11b4b00e6dbad3e379ac46444cc34ce5e3211ab2b4fbbb86913024209f2e9717d105204fbdc613bd3b6e32987421995a481059fbeab64a1a71f145d6f30173489f7fb2faf7ca558e34bcd5f37530041bca90634ddbd50293ac70558da89d4e048d63442d9da41c24b64535df6df83f20bfdb6e9e3704510d3cfa07338252ac66a8320726187addbc9da47e85954471ad9b2094725f22096a9dfaff9e2bd529a84a18b49f8e8e0e1070393e7f12df78216c655ab49ffe29326265d3af11508ed904faa6462eb92b04d65e6f4c4f33060d7f1fe4000234f2e39d250b674426988f9ca1f70a1f8cd4ffbbedd883b6e89727f96e65498b9ea4732a7be94ddb7ae314f749f45aa18f6ab45f1c44a8e6ae3b28b0192aa778bdf1f60e7e7dd93532d188d45456260daf02bc3358fb9a24145c22556d7965e6474a8a4c248433f130f9c6311409960e9c14fa9c61096a8c7fca6d072b0ec23ced2ef814efb4a8368139349460824cdb71c8b2024525ca9e8151f504038878fc11c215b3714a7b7d865d05d3af34b5e2d13183fcc0a93970a5f85a314437408104694745cd042f9cf011e4841275532840fb13f11b3130f3b48972dcb5dbefdcc5d1a8955f64a46e1d7b5946c2acf7c0597b0f1235eb909238d5dad03cf6d9a99d8157e0587e80d5a34afbf2d14c99e83159d2f9dd531b85593d19fbc4a354d6ce5b5ccd3bdd4d7a015fe105b815372e53afa41a8d5ace55d821f06f1b0736c2ba96873ef41420a558fd4003752a3a474f242e7daa631a7c406367c6d85bb51935c485b45d01c03ff85cd70aac01fd16b297421d3401194b77637a3638a7a1e741fadd040e49f53bb2c30bc4bb4e0a44b11abea654147462851beea27debb8e3d2393fcb6e8da11a0e1e555022ab3277e63d4ba4075f81fd52ca9b49f21193122d310354084b5af5395419a615bf392fd36950cd56d4298cae89f2de1183f94aa126acb148383a7b67b50cd83bc2c263c902847576ffd5d29afce478a907612a4575bebe37648681ca414c4504ae268dd922c0704fca369410758e869e7920788ed925125e7f56375e3080364415d5824c623e4758c33481b61efd8d6f9e701b56f4440499d328a23bbb9c3b1624c04a596448edd44f5becd8124bdc297924f7dea180e147278b643c353f8d4937530d58b8820d6f128d6906a3fa7e9b63eb4505cf51ca9d1bede8c2ff40981dcefab40e9bb2096b20b3547fe4c2600740334c2da14319b4da4e35eac721b33eb55feb11c02d589bf37b18ec06ca5abefae6c0a49182a1d8cdc5706f6f19ec0f69d8233c3de28eb1fd588bf32c7877a724e03dead2a76fdab8d3a77314057e82d7dca84eb01ff68dda86270499f45feedab1b5c4707adaa49ca909a1667c83a91a218051bc4526f00487e582532ce8fb9b66f0414049a32b43debe7ee1151f90c9ed5e99ccaa3a534956153d95113f72081a0be3ff3cee251e39d59760877aafafd1011ed395dab7a58cda625666648ab21518c5d2627ca06fb1e6f373f563d2e137ef122b975e83e8553e7b14d320784b8d7f326219c407fe85c4d622da8672ff1f35524f7d7bbb5886dd2c7d6da4f0c11441bdfb6aa245396535cdf01ca12880621d04d8bdebd9ad22f9bcfca49f8edae28bd36c8267ff520b975bdbf20f3e36a8e88db3a87a2e07dcf0d2ec39732f97047031923f8bd6e75efcca1223bfdab8d2db6a810d2c3c6dc9632830da85d8a18d308112008e735e7436c2dd2fb92e83bdc13246951444482e01ca1fd5e265b58a93595d9602a7dec2e9eadd7891e9de45110def4220c973c33fc03069dbb3432a4f0fa5d9047ddccbee4e8d24fe075c9e1a00578b175b66e7f217aac9d3fa46dd7bee1b3ee5a572fd73eadd1de22c20db4b5d7a9181b9caa983dd629145a64b5ea7d795598b9d1aa4fd3bc309c1eae14e7749b32caea935db227d4735c124df798cc52ee94fe6ee6d391130ebbae03bc09131d5bf9da0b383b7c74c22bf069d942a615774f24f802d794e4c89e68ae6000f88d1f4b7791d7270cee04ab3cc1f42be8f188cc96729b26358b398e442ddf9f288178feec32dc9b7ef5cf97b37b3708c736656aa0076f82ebccb6866766746ad0553dac2f0fff90b2795cfd5226e63647f615f7d6bb65293e9cd9260800b7ecfe7ec3326e22c341c3d9fd28c20606977537d25022ccb04ddbda1b7848416658458c803e4d3b8890816c286f5f086fe422865503a5001849d5f0cef86a83ab2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h76e3ca31bed82421626fd00e734ead4413f3bece4e94769c1c27e9a61ed85e3dab47209c02187280ba0b13f7a433cfa1be94a949f9bc524cd572fd2496dd111e29a91f22af4e14fbca1e739c26cd492c16084a47db3ddee973d0ec244fd1450e21ae3de698e73752cd20f1a5a7964220295eef77ac7f9919a4d10d48ad9888ea90f52158cf540f3c09198bb5bd8fc057c1681055677f83f7e8c5be2a363a8c251ae7d56285d7af4dc4e3c82fdf1d5904bfb21d970851df044223dce779bb66551931b58ba57ebc7de99b8f8e11588e4f9bd06dddf147de6ac4037415f00eb484d5671b47188179bed424f3f37893271afb8dab429ebfb1ede97eb026717975031373b6f1b2abf1d4567f5eeab7c7a436158b9fa71681e78ac6e405eec36580ed9bec1d773b29c34323089ca8ab3163e7ecc2f949d337a8f847cba8ef2b968a74765eaee3ef2a7b89505b321fb077573d1f73b7a8c9e5f52311d8673fafa1586068d13d8bbaed579d81364da61e6fddac70e7e6c77e13f72f619ce9a1865c80a65ef13516f3d7c00b8d942bd54db583241116ca89714069d6acac818d0a49a419d6c32fd79e87fc9b6fc1b14056cb7aea8b278e1e118578d5045e9ef75a1d6de4bfa35df7e976e129ffab07cae1a1f261c25399335dbb5f9b59d2358f6c1420e2fc306db910e6e361bd5fcef2243189b2198f91f79c252dc065106ca8bf35f3232d8be43748ea36f348801b1e53660538ea19c603e01fcecdf58cd7c99510fc936071c3ce14cfb9ca95aac58e5f38de01662fff282a7920976a0d1b2a4569da664f7979825031d27096433e04e7eff8c82734f73852ace16ac356af91003739b1e8db4807d5109d201be29b684387fdff8020f53b436ff7fdf668dc5a6ef06276eb3ea3ef69e7572201c137d66fc6f813dd19732d09732888703541a4a89bc61ce644dab1478872f214c11622477c05feac98382cf7b055df9e57dab338ae7e76040ca281d14b1aa31f0a1f7b1301aff4526ee4327d67467b639aa8c911780e32e328d433c528f08b64e4c277a50caa99c76775a199475eb52e10305867e8d34a4476967c994f9d06c9370b28566d85a54211eba6fc0b6ca212985ae27240817fc64c1d7a306814a2a52efc3abc3a86abe4f821bcbc8c2c7addec2a628c9ece4c4ac480c574800931a6300d81fea58412cebb22e5542e40de47a78d132e7ec3c012d299028766c6cb3097dc2811de9b277865100249baf44e7fb0329d8c2c4bddc6d0d72b71df065c6f417dd2cbf9bee2ce30574dc6ae40aed2aad6895aae8dc42b41ff687de2a1bc06030c7a3f623f7e3b786b4b96ea212237e1c61a9acf25590c8497d5ccc47a2b42f8ec08cd8dd7c7e108c4c91c32c710c509dab26d2e812b9002a3d09070162ba36e694e874f4fce5269132705b72a2d1ed86fba2ebc5bb5d7dd870ec66822ac2dcab17c334bae241bc3d799a6c1bb8286e7b2632d497b34c9645eb44ab79fe7b69496559358fbd1503751e1a6e118332f77f7a660b7ee92c9f09096409391caf656c57f93fe3c14b6048658153a64e2308703b6066745d64d10e2a3c1a132c279c48f4ec2451f2115097eee2e4a2857fb240332c1456bac7b3ec92226d561e47a47aab7e08c55906b671b4b1d151913d303dd84c0d4f986c2b4df387efc24a434a6cc0327d1e1f5d4e1edd4419b722efa4af65b704ff8a0e235211832d78ef025373dbb2c0f12400224231b8ff38eab8157550db6de237f59f41685ba034cfd1cddae0d32bad86737adfc2a26be7109463209d771fa57228f4a33ebf31ba7c2e05df166d5183599a4d2287af83ef3375834096e95edd89c78b6045b302b960f3b1de51ced1af2da0aed6ebda0e8d55de205df1a3c4cb3aa61c5e5f73d87acc5fcc5f91dc47b0d635ff0b99a1e7fcc2b7e733043d1211c112f3596a83150ebbec9225dd0555659c714ac37487b70f738f8ed96462992ea960e4ffa483fbe1065d41605b173837a148b5fcf29f0340ea4523699ddf4c83934780d3dc2ac36c1c4f5efac7ddfc9d917d186229e327dafdfd4fc75cd8a9050069c0333b059dca027595dbc449b7185a509b4194c6135bc48c51d26f8d3958564dd16349712127c4358579f6312bc90c270388cd7cea0d3ef86cfc37382fc40fc566be412c99bd02e115711ead3dc7da438abe1a5c1a8e269cab5779a7bd8abd4386629dfdd7c4fa10b792f064534c1bf0632fdc98daba02f820cea17828819d3ed02bf645be1c25781c290bd27b07cf87b7092e4e19094260ee0c1189d27445067af372f2bf25718c19d05890576bcaf478ce28018f3cb1f983b465bac8f4a7edf468e24126a06040a41841f5e435fd39a0369778a5ae7b2d6c01966d13e56f729e851402c5a7336b792bb34e836bfde7c2a4c84b18b96f2c3f129cac872461ea693385067e35df0e705e12095e900d8f9d5c25333ee04d7e8d923fbdec4d8d880576e9dd47e4bea6ac9f695319a35cdfe38f81720d2b39e20a616fb5eaef332b0429396cf7769042aecae1627ba56ba10427c152dbd9ab1618a6f894d305063b3f4e5bb05a19023f9840f51d34c7c441bc1160ad46a44c0d7c68d9443c3241afd42d04cdcfd99f0643b0bb8139627d481b6218b785dcdf7761bc71c70fa4dff3fe451374f5a1ad2a31f16eaf3ed97af4e63fb205b68851ce8b3a8a64e31526900467a5485308010a8f55ba643b9a510d36d577ed95380d5937d5fa5fba75e5cac42f70964dda19fd1257e50677c0062537cc3204d72395c9565d228c9cdec762b44cf32d7424b77fb1ed9118d6a245bfba4a99101f95de502d3a8c55a476f6d0201f15ddfc61e8be9e62e35b1dbc909f80b9da0bbbde81eb6070050ede48a95;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hda9cbce15624d6b24d224b89cc40ef5f77b0fdf1ad16ca6b388593f9c90f3b819975643205dbe27fa2c676e4c53f4cf3661e3b8745195a1878004851099e8d5c583b88509b8722e6c0c9f00917479ba49bb5d563d1246ddc96f25406dbddb868999470e052d771ae5ff3e8c5b1c09e8a87deed532e27d3eb365949eb41a089b7027cde25e023ca8d1e41a8f4bcdc7f5b145ccb74abcfb1c9f7ae6721f60044338796a8799b0d22182d479ee9c0f090c290443677db70cfebbbe380eb6224ccf09c6c9bd66d8ab659984bca086241ffc4e149aea34a44f0c2224bc237321a5642ebeb197c9c6fa928c565b6defd89d201a8985c5a13c8ae7de410a16e414df9aa2f7aef2a559dbf8076dcdfbeedd2f01dec910f9fb54b14a467835a950599c5f92bda40f0ede5d90985325da04b14e315e74b61c5b854df09eb28018779bb002a34caa935174b7edd8e260f2b3b48698e07ec0bb91a6c2202ddd7f4fd7bc68e551b006bbd0c789a74c44b8a83970b48bc99a32078c2a7b09aa468d06e5eceb7aa48fe40df9a678d8e106efe926abdc5e6693d7f6e622f786e9dd0be26d5062a9d4edc1e6024f44b6ef122333d15e9737113276df89377b174e760b349ead0e187d184058e6592d3c564799dbc39f098f5cffa428e32ca6a7330fd8a3fea45169882a2575e3814e493260cd789921a997d908d4f4dc4f8fba348c89bc34b549cd2659975d33f0cb373ba6d940d1f65f0627aa3c4438f9b705ad3227bc6cb685e03429340eb5b7599efea45d80b251383feb052e4f7b9f273fe89d8bb33fb8247566d27ecbb424b761290ca35f96f2780ff6c5530fdb6a64d84ca48c54be3644df2d657414e74621968e34cf74a47a39358e5b8f168365259d6abc2af0dc7f41d052dd05fd5f0ffb32419c4aacf643a78ebf8739e97839ca3d3644bb618729991405f9b342d5f49d5ba23c4ddde08de60ac312b0d591f120694d7e50ad09db660ef643d039033dc7936ee3d8f46d40afb9a0647b5b446b65c87baf8116d09d0b936135f7834fb288d5aa15ffebe94d82f5b35457ee7387e3684bf69fcb87896768905799110021a31bf4e3bc754f9e8d5ca5ac963c354bd5f5427e42bbf929fa8ea3b4de24a49ce1df3a48fe5f6ec154658a7712f5a512281d7e05f84723a7c730a5a6cc3359f753f1ab5753932fb98243b14210e5f67f1195e32fa78f1b7069e8bd31579cbaf474ba1ecfa2d9270b3296528891608831c2decce6016f6591354d8f5b80e26d16c6e832bb9bef208b66ad28d60251231a11d2fd244d864f9789f1acde41713f6673d5212fa610feaefe0a03d257d3a1ee37df7556f9a02ffb7713638cb7dfa39c523a3a431e65ab10d24a20d56d0a567a35b398e0d6a9be12d57936fa8c786907a7fef11859452ee1830d60b978b9ce81a891ffe294f4c77154d5a91771c51cc9e8ccb3419f4d4c75227fa24a053333dea003089f18c2e0455f2f5bbd4399698b4cb94ba467d82dc9ea019e0a1cd2d91ae248b97cc1d76c2b4dd4a3bd39185b30051c390fd9f1c1158b87b5207209635e130bbc7ebd18ac9d856d40a6fe9b96f109eddcb8b1d058854324e2c43aaf7a7e842a46651817f68237434236e8004d31ce5a8e7dbc8d64caa40cde1d84ab6f1151a4486d161e50925e3a76b7b6efbeebbdd869ff807702b79e4467d52e1124c2fd0924390d1943a426aa068190b3ebe907f9cdb2c78b413fdc8164d2ef45593ad33b9ffcf250c43e4ff499ba812a5ff329c1c5df4934031c08a66d91bb81be64f8c363196940e0807c7a05fa65f016df91b82960b253e2b89e787a9c28f12d4be4ed52e7e2fd749a391461ca4239829c2be0e10ac645db6d1d29e44bbd7db210bf12507399585e75a4ce8a536a74cb29bd0b392b5848ecf4a68c5a7e3e2b226d32ed06c52fd014a9d051f8319850957ddb1d7ce0c93010988f90cbeb8f14f4ca05bfed1e732a92b729bcf53b8efa013de2fc5859d892c7bb43a601a9343611dad1fce5a5181223c0f537a1ac35b17956bc198d6c43c664311c9735dd7183e664719aab77e93beeec74391494508d4bd56adc7a34c418c6c58d9e2c7417bddc5b730d382c92ad626537efb29de86a1ea095dafdcff52c4f9f8f7c81a087608d4cdd59c758ddcbf48ecfbc52402864897e7aebb857300e8071a42d34a716b187a64dbd2c13d3d946c0d2a348189b7e376d86659af322ab50fa0376110b355a3a115dc5981e93e7dffb41ba1a89105e57742f62fd2a5e6c0d45eb8fce841bf6fb93ba831bbf9b547d81a84f96619fbfce8b7e1b7f582c9c075f21174af14b04c948d1409ae6f8df29dee7cd858232f9ab385ffbc8bc3eb7822ceecd9df7e2d36f599f57f3932159e61381f8dee608d82231d8a811c06fd6ee1e5ef056784f44cc441c1b99a0e02e99671bb07c5e7dec21a911261e3c050b675abf029cb175aaca34c18e0dd21745ef0b67acb9418300be3cdc8d206304d1357552faa97e2e2bb24f9da606d1dc24c2ec663ff951629a0014d92bed493a582aaeeaefe064c0957df87c9f7937321b80ba43bfc7d9c78176edfb9f1fe57c342d43ad34bdce9979ded5be915450fc02d331a2d799c318ac3a2fe535e4f9b8586291d45b85757a1b794c0424b5f20706c8677127ea45830f406f2169281175e89168a1e2f46c89c891aa3573bc70e8afefe16eab652e549924c077578279c0d91a0650cecff2144bc9633af4fc20fbcccaaef5420c56e93eded31f0cec361e533ad3ffa334e7e66a6d1aec758ecf354e8f06d5025ec5e9dc8b4d4499c0b1a7b8b2f3455dc353e70ad86480275e225658042de36f64adeaa548bfaa1c047fbe9d464e7e809d20376c136414014c91af6abf35eaa95;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h285205de9c22968f08971280928c52f8ae476c389a3fdae7c20ee40fe1707145ba42b62eaeec6f052b61eea7b607a542306c688fd6c204900bb285fb6b6415bd926357a7da0088063449fd9dfc4c842c37a28094516f410a78567938c05cd7a70b124d7024dde1a3885e38331d86a2ada20c3931fcb5790f9557f507feef5b6d8e1432eee53b2b051314eb323f05afba771640da058deba5363583aaae37a4d6f50e6cf09c07ecef912310635be47884a0358150a0171ea0fd12e2ee4b621d34e3bb6bc40fff0505608501f0e50c2121349dcf8c02b5288c71effdb68fee4da22057f7e3471e5c4b49386d39d135f5a04a5fde6ba8554650378374f021f76bb8f968d73ffb5e144b974b2ff9aff3ee4ecea2b62234d3bac6c5c6128bb036e638d8c9b7e2a21f221847a9b9069749ae2c88fdd2822ab1e00f91bc49301cc17e07c37f5a5572aa680a1b402d583f3023903a4683d43ff0c2c73958b0ebb25616e68381da4b8dcf0be8f8625384d1fc431c41d79c2ca226f862fdf423a42cff5866a0d01f2a5675118cb0c1275e9f41e3dede83c0ca02d219ce9b817f2124155fe8ab110df0309d0a95148e748b96617ba6262d367e2764035ec6d009f59fad6a7d44e060e2eea37135c74cf3dbe29a0a92032eb9976202d9c22a57b765840890616fbdbefbf71c00938d5ebeae685bb8d9a8d78d8bb5a941fe2c1dfb3ad85711b1f5e34c81281e1063d7e017e4b1b9d6791a202a9f332eeb8918f4c31db18ac347071ad2e730783fccec4dcfb40beea28fd6d0cad55e2e067fc5d6c64d0e9056b75faf453c4220f4858aeb5d3251a7c203a3f8ccda03d43f3c56bd0599531a8289f6cfcf8201e37598aaf0925437bc6337320826f991714f9f1bdc0b4f03673cecb993c03f18b9baeeeb82c20261b98c3c717f35994527f551859dfdd748df7c3dc546bf6fae548ac87f8f22c7a1a790fbd1106bf566d53325523bd7d5344a7feffd425f99b418140db0ae4480835be9d3c4afd27c4bb85f566b7f1843ebf495394be20a743a6ce54f02101a31881ae233ca73ffa388cbb5d93fda42e408169f211a2094e9f54a550134083cf6656d495dcc7e5cf553755c3ac794a7810a5086fc758c42644116b89adfc3d796b5e04eaea7c2796763427ad975d289fe83b08875c6b8caa94549fccbf2ba995ab0cfce6e3198ab50e88cd9e49c2316f01a900ed3af3dce893670fca4ecb6f216dcff2ed83dddaa77601ec343bfd270f04e69fbf07839591934d88aa5ce4a7218f71b135b585aab3e6b9fb72230d1e1f323937fcc0ba14c0dbe7c8ce5a5ecba2726c5dc249e3f00461972bdcccb8f747cd1bb1ca4b9d2393548b939db1154506c52d3b5681f750f6f623838f9bde9321cd4315d7f438ec55d88a599f37733f3b2a3065e14147abf00fbc2999e472b9ea53ffba4ff42b14b1b9d6101c144b669bca417477f43c67bdef71ec2b33762ad345786e21ffef5f64728f90165a7925622d12092ad8f145215f7112b0bde48aa137bf7b14bd159fa0ebdc5f07ce78baed4d3b547a916d07331a1590113374ce61fdb35e43478f23067a3077ad4d30dd7843d5e37156b826efc5b5de7ae046eb295298eccefc6ea7b5701ecccc32c412060eb0f556b7268e59b5f3277fbd6277195127b664218a26c9f60da746e1cbb36cdf53e027d018462cfccc270b1919e083f525f92bdb9bcbfd7790d277185d0ccab5952454c8f1cc7fa0e964fb4337289a506cae017ba63b1e0af9387caa0a54029e8d22db1eb947fa5f9e8147b86f44d4ef53fd2480417a6b28588ba3123e219c9477ad6972b79679131cd3808ccf4f28444f2dd81909026ac6c7f0c0ea7a89531bc3bb4f81201ce4cedda9af27ce44ab53302b4c4fbbd63f7396dcf5904357cca8c787ad0400ebc059f3ffb5a8f1f7df1a3f66ea55108070b788db46cdf27b05287ff8b35d66612150e216cb249980790408cb4d5f2afbcf7f2dba4eed7768dbb9f4883415e842d317c1fbd114c4b7fba853cef57e0924603940d4aac801d18d65524247a19851ca5cdb42dad8de1dbec9fdef6935200a3c02f74bbd2bbdbae8c33013d1360108e92604bea4b8aa920bf374685f98d3b92e783b07539ab95550fbd5dd374953239ab2de8fb66e0cb732adc4548c680603183b7601a22c9f5b6d80cebc155876e64f31a52769e41894a971c6b5fe3eefcb0ef65a0847758a9da5f2244172e473161595d1b42d809fcca79e7f9a0c0c0a08158667c69c33245e5046a43eef094caaf637ae0c23f2238567f218c2f4e253991775fc800dc78fb3288645fee5a51b6436fbc03df58b420c435fcd3d8954d7e1434359ead98f200ddb25842a3f89cf2a1e63eef8f619777516964bc22e659808f571e51796267667dc02f78b941e2e2e245afa59ca7482255f3d750de7372006aa9a8e5cb3fbb7ef3528caf2e1765143e796cfdb8632c0329a44dee863b7057fbdeaeabdda6e3cdbbed51d9de8df8d082c43a8fb381be02d0c57ebcf49b7212aab36cf3285ba41c15031007288925640ced8dc3325c2da40d0434dc6b934203529a300f66520f11dcf64e1720bf4b096849f922b4aa34704fd45db6980fd03afc25c3d2ca829a79d0f48e414946cd93b5db9dd007521de7f01ee4f542eccd3ff9d227276dcd47dcd4307fe29939c961eb0d85cb1e3e95a249695ed8b8ff7bbccf6922c460c2b8c5537cb1476be64b6ceb0837adb30de5aa1c3643a4a2e9df9c0b8c49312530037e878a281ece3a0eb924b4548504159331f590850efd369c783aa18272a7509e7b1e72d869a2157470c31bd579c9348a3e5620ccb6fa42552dc29bf0ae90bd5e5a3f6c00c9e23aee3e6e4eae00e45f0e82bcde2a790842;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hfecaabe3c8c4680ec8297cc579d8f381cf8f0988aeb67e7e4f1928941a08e65bc41d6cf3163febfd467347d7391aa97726aa4d56e46828629d73e3bd51c0a41ea0d420b69b147a9a5b4b3f0911bd03c9b9781dae1012464f79d31f9ee8f65ee90a96ca84402219e2495782041a17b2b43b08bdafd97c1ee844a7c47abb6bfc950fc3cbdf54246ed3ed8923eeaa665e327d1c4cc8d7843fd3c09c887bc09336b3b44b2d5b6a414e23b391bcdd3c503140a945a6f574457b79a98167e5bed49eeaed6fd0fcab90519a4bab4a776c6f32bb68904407cca85fb520cd1f6bf2b59a7e871ea57ac645ac92c3520ae12f2736b0ddec02d484d8748528ba2bb26518b915873a9b658b0fd93346c1445b4e21b0771a33e2466eeff9e69c9516d4dbe35fb599068d40bbdb24d49b895f659079b8e172879f73b7aad88a5e022fe7e06f930d7ff74b75c3d6327490e6ec618f8c4704d271fbfde0da67cef1cb02cc38e7619c83dd14c21ac682d2cc1c5f0ea9e8cedb4b1ee6ceb5830c5b929d442f4e87f66cd60ab42a6a66adf9668ca28e2b5d879aead14061ac8785156a71912cd83e8553db3e864b9f00667bd2bc4c46c8ad64063577a4ddb81ec8e8c97aa6a05d08cce03725255617718143e7396922f95f27a1a76bb43af4da941fa99ffa02887fb48b8d8ba3ebbdd97b849cbbb2653ed332106da4e30fdf04d326d00b1f388bef88a95cb944f706b7c23eb0499b6ab38f7d93a3c1b8a05feea85ba604242e7aa82c4092878b3d9e9927552ae4ef45761d79bd9563f7be7022dfb772c5d4873356c3ad5bad59eb3bfcbe80bcd545c89e854a90525f8d174c1d7418e2b9663ee6ba3304ae0f15aca8d79557f2467fa59db4224d9a4985c48d7f5e09566ce4754e16410f073ede98571503f51d3927e5404911313d08111ade3ce80c62bbc6d73abdd3200f977ef1f6d8cb031526555eecb5a161de4f47b75230021afd3c9198f1984077ee616d5b6732120154c3a56ac7e170e50f812466c3be7a00b5d27859e1ae6172f16dcdd403c6cb82b90a592efa2b7545c2050d14468ba6476ff5cb10974191275cc4a55238c07482ceceb4d52b6bbb5e46ce35d6047d16773463ba85d3f1d892ac7a0bbf49634a09021eb34fcbf02a8a96765155fae79a87171b4fd98ba5f27ca7954eb3bb38afe126010af3c51c85994756d3b96339a7ea52dd12a4a23d516e217367dae09eaefb9eabaed5f637cba81f60e86b2fd3e7d35b47ee66fbc244995535936c693538cd83cda8729f131763c60bf73764b22571bf3d26746b3a2f5e20cad0e91645f04f9392bcdf21ea4d4a2d26061d8c524bda6fa583abd9ee6fb208e2212cb559fa69d125ccb1da5b9f527abdb946e15cea9284c4c9bd788b701d048ef795cd405882460abddbc965505e5532f6a3fecb9dd92f67fdbf4fbb0157b5a8d63b3c5680e59084670ea29a9d4d8a301a5a7d10a8439ece7f47e97be238105e72c78f4dd05f9711cd22f28a1fc6c3013b768a9fa48a61cb944cb4f2bc123b7d2132a7c473c7a8b6885b0b4683b69477c158e8f69f7808c0900b84687d531670a60fd44fbb519ebd38f34fac6f2a0b465f5dedc0d676301214d66fa1c5d2f4e775a41624ae261d89b9c46f9979ec532e75972ad9f4f51de16c53fd567b925f47e888195e2bab1539b42ba9680f73a4f74d89412e9122f65a0ab3f6f72d114bda863250eb8232e1e07a4232bac5dcf98dda17fdf0d63c64b02347eb36be7fcf4bd775726894db7ef8295d43f724a843b17a2e6b598e3c90dcf77beea0c22faf5712c21a2a8454cc4827ca7298803e772f2bea4fdda39b13fb45e405b466dc6738376b6199331e5c95b79f2113fcfa07703a06b59dc3d0c58a3bd8d054e61aaff1e8471942dbae33519a3d73ef7fed4ca6c613ae8851e513131865a3f8dcd0fde0b6fd933e566a4473c06608806467d259b0941ae95228603c30f25b80c741a9488f64a43bdc7e96f0f2abb7c2d6edffc11dc3ddc11c7f9e034cebd853e4dccffaf1f64a214eae5a72de6e1cd9e77c2de5cbeca7fe9db3143d9ba3d240e1a8a8cf53e99d8d515be10338435eaadd57224fd8aeea973ece84070d2753e17b7241a41bb9248abcfc08e797b73a0a65ab5217e7ab93ba9d0ac77bb23d28408d9227595042a13b5be496d2aaec0b6e1d27881cb9f2c112fea42be85a06af35c06141424c9e30b28075154bdac9029f881a8058e313b1251ea9b4dd3704c86c6e5dffb98c1a6d50054c19268ca4041e8577c124a2ad7ae6aaff8a92949127b178c2ad176381dc06044bb6d047db81ee36e19fc778ce87d4904e491032ecdb9e85960c0eda16db82ade3e6f219b0dfb4cb977ee558a1ef4291253bcad18ec98ca453ea6e0b9db41650107bc8e3bc295957de1ea7b60f6f9a9b0f7b9cc0cb6844850f289cc36c1220e5983826802903aa241086e1b1b8fc94e34c3ceeb4de435c33d31673868aea442b0b6d4f36295658a2ac06f80027f09a402c7273569c6641116688c633fa35ea897f339db093b6d5a9f1bae52aff491dcdcbf72db66a797e4d3c3441597926d0470f8c6f965b43e2d1bac27642914f72e518aa70618154bb81e26b3c992a06ee5e39e5da693f74470f94b128bbaaa681f41008e10d09dce7f566d60c77270f6f93e4cde450f76c813929086a47f8d024a22c4ab46b9202aeaa8e11b3fd23a031e9039227d78c1783b24d56163dbae7ef88c6cdf568956946ccb530305d835fee0fb62e3dec1d5d13f876ab5e290e03a233cb4d8d116ad05e5d3bfd3fd2dec1f5ba0bcc3258e48dd41287af89b2e4d030b6680fd93612baed4d80d4e4d289093053aa0ccec929ef50b25ababadabeb76d5929807ace3c65d5bbe4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h41febcd9c5d2e2dc7abf68c3a11b13844074f7e4a8439f6bc894ee4c472e08681a05ee833b9f786ff95a9f49201759f1df0ef8bb1fd548c1a081ffe69207fced2bbac34a7abbea116cc3e17a9acb6b4436f5f103c792c9bbc59a66ed4a82c1753b45058533a647f6a21cb2090c79c17b7fb371643b4170a9b340b644320a8f26c3632c77e53e546dab7132f84295471dafb7c6a81476f354520a27287513d91331635db5590525f77897d40061bbc5a8132a044d740efc3f6768975855e279c6bfe1184c85d87143695558f04244f4ca5d2c66d361766925808ed137bcf8986c27227dbfeed51b79bb8218864129278ade38c10a7f602ce80f9cb5e8392bbe10d85eff2a015ca8328474f114f2a44589c32859b6b7ed1d6d52bd65836e3123ecd3c32f7bfd966af629b3f981a5f5fad86731e671f315d96dc4ebc8ee9c1c9f8fcb5d79a25ecec0e455dfa7a614fe3b4b12158a2fc1212b65cd0beb190bc83b2872db240c36bb186dc57035c7107ee50bb169f319835c9abf36b0796c89316f70bbea908f2475c61208ba19261df6e663cce219cf01212e658fe53519ca26acb4d9299ba6e5538f1541c66070e5ede83e94320cc1ab25d04fde41499bda19ef53f790c3a2c04fe105dd54a9f46a87bcff002cd7ce2539fa319dc0a562bc02a3b5d1a157129004f1f51c353a9b6d68c3d1f100ed0f43976b5801f90b4dfaf9126820ca798ff6b5689c989593e0fad4f552a4096184e0510fa9fdb9fccaf117cfe7011690f5661beb7914b549a4ac7bb1c7b3d9fb00230001040b283248c2de9b4417e139f48b97d4cc6755ed0ee923d913951889e5cfd65d7414ad9a131a117480d42f382c6d1ecc7cbcecabce2a399305b53bf3c565099ed03e161705bd2e0d40b21091943bcd1ce9013d19dc02b3c8f92c875e13cd339124b005641367cb8c48bd6428513e4231ceeb87d10d8409a034476d1c5a3385d8f5b6b9ae96c3bc960bc309fb79a7b3420493d2ff346d659d48a5b57f121fee29936a33097e17603a3273aa8c079bd3a26c48bdc81e281e7298cedb5276a17579982a8f979d292a63f127651e51f0d89e789ce588d8f22d6ed49a3abf1669cfdb4dab6b328e332413006104d97bd33b6dd0a727b3fd80ba4a0982fae384df3b2a57359a8870ec78ed34ecc7bf91ad7b18cba8a4ae53fef8ddd32dcd93e9c856ca010436e2b0d5d473b9d4292dc18a78b576444c1fb139d97cb31d5a98849dbc583457cd9bd126c5ff5ef578c9d89e513ff7ca6bc5f6e896e17c881cf4fe84d5139f93790dda86568253028491e8ca248d597b66eee7effcd7c6f83da6cd68177b1ea29fefaa0634a1d997984849b8b749113ed4bc6a57eed00b2baa3ffc6da31c8eba44c66e2162a613e7c93515b2c9725831703d1025bb9864271db664d4c81d729959788a9ecc46c55a1bd662a13862292bc6a54afa7ecbab112352d60e2a29674b16208264e25c43673a355fa128626995c7e2200319da633eaa11c9244375e2013a5ab9710ba516ddd49cd9a0bef7cff182bbf5a6961f665ea49b1014255dc72ac269f34ad0fbb9310a956bea9b05d7092b4f50ced194bfec4f61917e49073758cf82a03ff121fa7c8e257c11b5d6397ed1546c08185cd9e6968b8813abba0b8709d90dc6324114f718c89e179b53c03882dfbe28a352757acf03ec53c38b533667120c8c2dbe009a64e25fe759cec18dd8194c5a29798029bccfca2ec5d891ed6fc1bff6047c513c0dadecfbf5cdd409613d7f7ff06c81d938cc3ae57af09c07d6adc03a612d76bdeb84a9af23556c5230536664a8279024ba2b2ba82dd728df842ae18929208dcb6da650dc688c85ea06e767a1132261a8e8ad82520b6789b1a0560a31989cd43708f05fecaf7e397c8ccc6c04ec0ee643bb11c58e698322b9b2ec3b83c83337b6594f7afc58531e4accb568c3c64edfa5ba571b928e6198d20f6367fa378f1fcf69f3b6037a8d0e16a4f9d167e561ac23f0216918fe3239c51d7cffcf9dbb1dd070730ab4ef652ba63f774664e80985c099580625a8c67107220f315062a182caf3abbb0668192fec4b7914bf34243bbde65c4c4aa7ef9a610115aad18405dc695376e044c2a7e3b077b113f978f74a1258261ee367b344519e152af9f82d06bccde0132ae1fa63064f1c87101a7289eecafdf6f9a8e94f1706ed0f793907c7736987c13f9f8497a2099edaee7059490ae3f7cbb06c07b7f4cc6ba419ab040caafe05c23e2e163c9c27b6ee02f6f3ef3c8a521efa16444ba7ab66a5b0228ca4b37ab333f7314b90f9f91b3ce98fa292c21e52f53c2f8b9f3d99c94ed8e1234308d92927e5593b325b9a92e022d16dee4b1a11def199e8e5356f41491109650eb5fb0130c090c74a68ee21521706e10ecde3d1f626c4bd5f9823ed064171059eeb558826d12034bfd28c107cb60744ce0befd924f9479629d4af76e084d587c3e30caa9b4aa6970d1a845412469f38286196f015546cd0e2d18c5a5395d39332bc6f52d64e9421a388cbfb0f0543dc0b30125ca09258abaee46724766223c80cea682972c3de3feec0599f336038da1eea362383a495dc996dd2c75fcb67cb6f82899613634cc816192428d48e3e925771675bf5aa8a532f714f7f1bc0b70b702472c37d1df0525a0d468c149e02e612456096d6ebaabfeb6f67f809a975184e274b147ea62147172705f6d84716377711bbbddc36d0bf2b28a448015bed35ed117f83c5de94c0bc65e633be116d62100a2d4aa48f239571181e2684dc00822405cc2055d4c8dfd28b45be772c3eecdb54cee9922f9e90f1e7740b02eb63a5cd86baded76854bca565dbaf0b7dd39323d20a97250dfe84cbd836e36ad034c582;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h450093545f748f9f0246e4ff932bea470bf37398ad82f767a32367b1947ebfa8252186cbd31f9546eee18882a0d0ce6b5aab912a26f1cc36c8140521131615fbba7ee9fc09fa509de54adbf9d966c865e9540e5287d5b31f0b5f6f46a66ad8fe99bd1fcb4336fcd61186e8f72de6f13345af68f8398f524091f34057f4475f1cc6d337afe27c57cba76dd2279cbd785962e68cacf0d838a41cbf268efdb486101369e31612028f1df6695e2df9e97a4a53cf2532cf54cbbf218d871e4bb2bd66b3214308b5573d916f72ef6be11ec9bc6be5435e879b663b6a8f0748a65a9b34068d9b0b12f614269d02dd35ed8d1b135808e0c30d5203e1e09b5dd714f4b2790554ade0f116ce24e473a48b3f3b9cef0d8bb1a471c28c406b00a49d724dca690422c02201ff72ed6285948a931426947bd619110658fc0e18227d63a00cdcd71d97e417aa4293ccb7a3269d6adec181674a37fc25b978cf886f29141f0896bbe042fd74121da44379aed275d986c64f19a61def7492689d544b409f806ac26a1aabea53e0f2bae5ae28c0ea0dc4e370683ebf38866d52ed8dab2dd3c01414a4f6dd1e8e9f959e98fb381bd28b279bf8f7ae7cb35358c549ff3f2a5e4f30c69f72f1bad6237f9aa20adda102adf8eaaa2dc457de47181c7284347dfa0e26352c633948f94ae6ef4e0ce63bc6a11552dece5579b1caa7fe29f303fd13ee3084ecf8bcf55dffa8ccabf80d5598b91f01847b473aeb9968ffa29f2143883682551e6b5e209a7eb8b77db1c9da49352526c7221ab4b7a2dd978b8a4be377e0fa802b0ec5307d7503e6a5103bdb7f4a078691662c9e936d2fd417cdb188bcb0238d79766090df5b1d38d9576b1c42ea6104ebd927b9b2235d32058f58e6ab3682fcbd33255f2f51366cd4f84d9a129701e9cc64a874a3082da04ddfb7067ea2b09f7a23b2cc53cac56a4b7fa7c44af687380ceff9f376ec29d0d4b49eeaf6144bbc7555d483a246c1d0b71562c2ec4ff5a796cfc84756167ea9c61250656019d8a16cf0f6ac94b6add16d1eb89e31b17015e3d7c172f061ecb525e845f0a96f3c40a6cbcdcb45ce10458a682f7a675fe7261844399794963a8fe70ead4a9558cab277aa4a7e3dfb7af388f58ea24fbe1ba14fccc913bedd719ee24f3f0ec776a4a8c51588dd6e2190364607d55f9ef94942fb0b0e33c307dd6a0fd19cd480edebf52b53e3b8c77d20e4bb422c1c59794cb1668a231dfa548ade9e7ebfcaededca4f233442e3939b026a34753a1a749efdef27e3f0cc5d54624a9c6a66ac56a5531f20da2c2c238a245752c910f9c587323e8fa2061753b36d72dc79403abc68c666fa4017b90af562c65263f52c147343e7a30f66279836054ffd2fa7e644d6178a20c4ec9fe2de30dfde43f0e24ffdf75b426ceab339780e43849f3e393a745817c8a13cad407052ee4498fc31d0e5a8d2f9a5dd4f1a3696695fbf4176bbbb8f8112cd3a67f875eeb70242e59ec44686a0b8411b23d97ca593cd011d9663f82385ba949d8401c55584e437f5d077ba906d249b87d2a9e1c30306d4239c37a3826c07596d80ec4f10e83643636b4ef646d2f984c797f78d274ff1e66b1345ce4849a5ed3bb6e0e5079a309c037f4efd241e60bb46638b993ec78c4e404d45857f5b30d44442699908dba9a830f3c2b550cc4e94aae584c0d9ed2b5d69f3470baec457a337399349efa9f0f118e47997a890ceaab63ea58621c1397f4c510b8b3a8350b87d1618b7e40e3af785d4ce2a7856d08a3208a53d58ef55f853f27c320502542d0c6229885d8fcee7cec446a48bc2d0eb210ecddbd337c4cb4bdb10b008d788b830150c62842b9cac80768bdc5328b3ad5e804c77d97106e503b385ab6591192512a5b064d3e285b2a0b2964d757aa65ad3b3372c20f37ec51d912bd1df1f27cefd27e7482639c2443c967f118e81d6e814e7915903c312f0116d778784cb130ce040ad974f18e19a6898fe25c5958cbf9f998ce12df98e5dd1c629baf7d3e14913d544e0390345043d768b272b5a38846c3b640b466b5988bc4b1d33342c1311e03341591895fb99949a50a2d1545fe7a77a7e0b28d18083d0a8179e01bb85c33a1d41ba52cec2d9024e4e6aad6a4640a0604b47c7df28afb7184fbc6837099b552d5c1fdff57b8dda85dbc0d88622f48b1958c3237d56e9dce18baeec40b88c868ac61b74a81b63c132c15213915a3d199733c190cf13625cfec2252df687b6317517acccb46a6c4c2766c4e0bc2fc47a669a2cf2e4679e1a6fc7f4114d05e6927a1b5335d0263910bb274dbebb28628f2d605200a3b3e864a13550da8b306d3a2f7e546af184a31ff4bfb0591f2a2974d216b8541d9ac6269e235a9381a33fe387dd3f626d74540fc59f70e959aed5cb79853bc959696fc904ef0fbd0079c18cdd234c03bb7b414c6417b44b5b0d1bd9d0a3fce6e07be77bd325b3e193c4e9f7625833c7091d079759e5e4bc0ed9e3d553a5994d354dbd37987797eb0dfb0390670a89d7d8eb039078b9875f3fac6d05e6257e3ef672dd7619cc9b401f5f3b3b03e4d4f4beee2973c074268f92a95d76ef6dc31d73307304358619bbebd8df555f45fa1a18106ddafca9b82680bd4b3a80c4f7e7256f25ff15ada995b951bf6731861570b97bf93e4f204144745466a80905f70a7c33231eccf00cd8c158358080311cff709392e22d2b809c6b5d75b7d170f4e952dfa3bbc2672bb6194a517308dd8a372f3c603225a447c0bb33e709c6255574d5339abc0d56eecb872aa12e8525870186a06e1f20bb28540f9c7a3a2bca8da15172c02b4a6eaa27154b643f18fe17600b8c13e89786d72de69bb931cc73723e1b1d3db0acf596ef5c51;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h59e98adc99cdc8136b6f620c3b5d3c1a2de5791e5682ed0dc978c61636b62f8228b0067935eaa6a7ea4bba3b2415226a93cdd35e8e288090402632d6b4324fe3778ea6a5145b7ed06d0bafbb88033b8818bafa6362737a47b836994db1636b1e1d3f6d3ad2c9405e4e6614872cd61217eb5bf2b01941a5df6cd369344cc7582ea4f8451b4e39a110151903be328d59284b28ad474ed52fdd220536d2b3ea525ed9402983c96e09291006f7555def07f2d6bcda7170e04edbe056e306dd306ebf4ab097672055b8143b386fb39648ba390aa07ab741e7478124500ba5750da9aee1562168dcce966bf2db99214b596bc412e5f4590cafe3407f6f52cb070114d304285c42ec1fb6e87ca6189c1d49dffb078cb567ad34d671c1a25bc215ca442acbeabf96d2d0b0c01a97dea48109b25d405a00d6dee75d546a9d1aa1b6afdadff18e3871fa5b54de4ad1357989719c76c0d9fda53cd6761930ee314931bd4da8dc144dcae5cb439c51ae5216de1125bee9860637bd66c8c45efc6f009cc7c65786a161d8f84efc9d43d4b4a70296af58be284b41c5fcd42326bf451c188c77a1e208a124383e56baff9f6582acb60a47f46188e5042ffdb4b3c2dfe3e9ea1190059a349fee4f30e5d1c46d859b6a5f45ba1ed9db3cc365bc643ec4f773177ab37ea0059ec07b0781a56ed9c6d6aab8746baeda20d35357fce6971e7be4eff6409c9497ef8a11b89dd87373772a55d5a5785ac126edca17be5f1f7aff61850582e0f26c097f0fbc2da4f26a32c03800203ffa74670ef56da7c08228e360880910f4b1e44d26d4bff786a35ab5d1f01d8c70e54d99fde6cfaf3c36b9e2af8cf3362d754ac7a12a57e32a85f61a87d5a43f69eec3e9f849411eba07c551ca798ccc0ec06c3b7ca9f4db732977a9a8f20b9a815906c8f8df71ba9d1d3a79c84de950555f86399ef8b15b8dec176ea4fe1941eb4f05cab02cbec92428bd22edd3f5df81d57830a4a99bb03b1cc364619e68e6916be567759e2929091f32576d589e44d6cda7c7cce53238203536702ff595fde72f499a314765ace704eebe7a472dcdb43a57e59806a2eb0c50a5ea23ca1aee1df024fe30cd07e7bf06c3772c723b0332c37a17354dcd34333f95e0e312768c9297e781072706284661021078be444263b3d4abdf4854f2e45429241b9b35b3760414d4dcc7ab4c3ac76af2d8cf6984563d7c2a9292c07f2dba32cb3158da4d6fc42d0b3b53f199748aafc505844b84c628e9b02dc4ea26b5b1de7919712c721b2e3e4828dc965d9e79542cdc1004216d77a76d250b05bb9e70678f4ac02f3bba4eee8c7b3f909625cfaa572c038c83ed34b45eff006696225439b92624e786288ac3cbc9ba9bf564e681b7e2dec4801cbe82e8a5a94bdc72591984b788c84b4b69110845b10c95f9e485d574e02b83626571d44575c98ea471691fb579af92fecf7f6bfbfbde4d7f81353bda2ed90e0c3d5082c05e2ac0a61622a124ac6e5428694fb84f77002356de53eae6f4c94ba49852d717f34f2eecd67c87150ce9cd7f741648d425a957a21d92be1ba8560a1b9d143a40e84075752ff051843c2e41523e9ab3d039146cab6ef163218f781e020e36eaeec2c896d651f84831cdb9b72be7861db9252f357708d03aa0ecf05d59850527860804dec71fd999b180beed2d185295245bb76f172c35add45b5872452a6ab948c453d752e4b7e622244f60c0eb4793a003d77ff7e262ff55ed61f27c076e1024477267dd4ce47ef80ae04a8e5467faf1d7e21138e3909d9582d31a77fce5400dd5feb1d522c2d6e4b997f47f7958f182f51719211d81c6a6a53364e274dbb7c9cd7f3abc26fa0976bb673aa42aceb2420d0c24ce7b26e1574f1b6daa0824345c4e10a31353e1f8b357746c5c0e6be202147b035840d1bff48ec744112552e963353b68ee8aa421bdd9267e0bd462e76323d1b1a99a44be056db5882cce25dbfb8adce61e0aa40fdeada6b6a1e06c388adcf7ea1ac049524f7233abf0ce190be483a2901609ee1d92395ff8e639c804a7678c04c038626fe9040d7ef98575b6eb03ece382cc7621ec8f4e719fc758da859cffbfb7005e404e9d8eb29cb15a3fcdf6ac77686c5da99aa717e4e8bf16805abdf3d0b1d3054b10bb43068686e6b2751689f7bcd8f410bbccf66454c61c7dff3ae94d64aba7f88b6089cacf33ced7dc6364a46f1e0da7f6578ece08e1b665cd475fb39d8915c0737794781d16b26b64f020d866570b583d55b727ace9adb58580e988759aa05b53dcfb9aa3c8ad6d6d2872360e10bd8c08a4d7f46fd3e8675771f9c586313fa7146c100cd909ade0b917c97d2067146bd41c99cdd64275c395d85dd6ced774766a078dcca16d7d14824a851fb55bbc990b85f90bf231b90136d3f8f3e9c133d1dc82b4c058fa5bec080d269df3706592c9de9da9fa72667d8fab386ffa5372b229f8189cc23f630590cadf146591398aa51a35b014d1c3f8bc428679e01d79829cab80f48f7e6d15e789a8568b354a7409640557a2af2dbdaec0d4b911525a836bc8103426868426fd6f92a22a37562327c475281d48e49d9750ec3993b38f556bbde97e1f3de458bd17041a0dd6b3728b8b4ae7b9b4e496190e761598e585c2cf93d02ec91b9bcd987374cf0e3fd4a1295242041391655adf8483f672a6ffec04367337fcf2988dd6a5d9a6456d64e21c250676444d5232d684b1d888ffab974de66c42e2b9746649a65cb1dafe26fc086a5a02432430a5765481114adcd5df3ef134147c2ef4880bb2215d4b0b30d5db27c2394277649c789772541bf019b9f70b2efa491b96b2e5170a023dcddf25f24f9ec36043236e6eedb01b0350e5fb172a3d06;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd4b3f30498c12dae9a6751754ca55f26bcb042a1d30fc9f8eb4a893334cdafae300c648c7af8c0eea44b25ae0c5dbd6a7e8e3982327c4ad77b257d24483647946396eb34783d80c3df5072dc98453e7ffdf3086b91684c25abda338f69d54013a40e61bc5a939a235e5290533d5926ca539f591dc0f91b9590b5d989371a2c6fa00c901a340c0f0c38eb025160b0353b234b3663598fb46ba483dadc84b0212f83ecb3c2ecd9e98b302e0253149cfd68d9bc6ae48955664378e53fd0654aad946c4235bb5fb9678fb60fc46ea281cc328cb4a119b4dfdc1783783dfc472db7724ca9f5dd6f7891ada784d8bb334ef8604af8982c7d61d3e1b4cbfc683056c1cde26a2298aa567c270e04a93c748d2e3cbe632369c146bb263957735b23f526b13b3f8d2a8fc4582314a95918d5460697d857e8a82b91d6c82be4251b6a78aa3c753c033ec5fa0d606a47cbced09ee5073aedd5b1129dfc96ef7b3c12dd6a01f89e361916aecc28121348ad62ff2e099b89d5bedf155f2d52e639282e581ff51a2c39bc24563a428ce077667cc4e0b602a4b12fcd3b3b6baa527e440d6697cc408bd5c6e423e04d4eaff0692fd34c05d3e1b8f10933cfc3c1e6c9f2c2a9ffcb63d02553d160059e9ef69cabd06043c34d07792388f57e3ef464bb485e00f67422a2ce973d53117b986dc8f655f5f6da2e10d0b0a4fc642a7c5e49377cd16ec7b845b141e4ba71bff45f68e089dcb1bad65a363b8d024fd6213bd7213b060695497f82a563dc6c13989c0ef37c499257f25184c7eb4a60da6a987658c34ed21303e19177105f70cbaf83c359aea5d662c36a5a4b8c9f79e8584e7813dc0f4e8031812a805f93488747fc4b1efecffa6213b4ffcc612e91da3daf176ef4193476b19b6b8870154f6d99c5e1e73ae23b7fc813749949f62e9b82af2a8eb62d0c9a6b73d22c3de5a527a16c15bca0aa41c6b1364a0939acc7eafc9463eeb6ae1e34f2cf1076b54cebcd38647ac2de4bae990670684a8666dc8959f7c8af1a1f49afd2b6f956530e1e99b9c3c6479661b166cb5bac2b52fd90f014becccaf1f7350de6cd8be5bd577b94e0d98756ff0315c4d461d79bfb97233fdcad22da57a9e130a2b8c0a7fd9764c9982a6ec0dfb7bedf3f529955f58a2d9ddde1aafd3109b885861cbfc3daf884e51ef73c135800638fc3ecaebc3701c534aec999668107d65e3c8c7f4c7871c4647d17849e47da79bfc73886766ff990e7f5d9db780b1204be50fdecc760334ac57b6684be4ee5bee20ef6598e34e90e0b13c545a565d0eadd0464459d25c4f8ac71c898d1b46f95619612a6744226c3d0de3d12ba7fcc3bbd6825f67c5a002a1342b0905560d8bff6d89f33f7347dd5e7d11d7bf67cba02c3e2e274f37ab24116716714b18c8e8044ca2cac84d4a8aeaab60c9857849ea0df1c2ba430d5b1fea8577b3e8cebe53848bf200c4e153b99967dde258476dc9dd158eed6240cedd9085aef867609493ec3c10b977c3b54f0df29902c7e993d377412e6e7cfca0043fcf93175461d57c7bab269eba1b28d1dbdaf41548836006a4f5fce5fbbe48aa989478cf963019dffd7de9dabe5314d5da7730ca470e11713b01cc5442d1e806ddfc4cf8752913b5e46c1ce658abe7e72fd0a83123b5f7d20e8e13c39bc791647f541d9f31397b43c32e2f39394769c7d7a5ec62ce28dcf524f176a4109bcb5685b99076458c5064cdcd4b2cb094b0c3f22ac3cda71aa3998bb936e6a3aec8df355f1d7a426e88d7a461ea1281624ec4ff5792ce1e49b77b9241306dbcbde1ccbbe00a42c11a6a83174e271ee5f0fcc45ba93f9cb1591c18f12da6afc4678476330a069d4e9a71376622dff78987316426f981dd150d932514528a807aafe935fc85a686aa0a9bca9084152637b7cbb610d7b91c4fa471f136c11278d96df8f51bb6ccff21156119e6eb06f97d12245dd2e480742a9f699a49630b76666b9c78354c1614f18dc946838499cb035458b84f6fb64f138a48d8a8abdcc3eb37a3d97c956608a49aef4bd3f221b73a4cd6d98dc3a2bbc06ebe273f85638b4fc4b51be9fd86cbb1c6ccae79c5210f31a9b2d6d62aadf3a84d17c2aced10ed43c552db39f42d6f09f8e961bd1772e5b4bc81e6ccef1e532700affe0477db01566aa0f438cb0907aa09dbc8997e63178216f0c0461b208bb01c814f3d7f1f7e3cc36f6bfd959f0eea3f5efe2fa6d9ccefcc27ff624764374e51bcbb451023b0d4c60404444e8c24aa75611b69589f636b3b81d722aa16aa9741d1fd017cf1b2b3dc6523fac5cabd65f4ba77348cd901bcb8b0445ae5587b018e553431d8f32598be03da1474a4b3914d0c154e739dcc559bde07becf09c1eba653ed0a855ac094aa24870c5de0f0f9b665a6d045c9b3da5c31376c718c342223b9e1666005405003a68c1c49cfde04ea2c54d33b4e5b985ec95957a6dca15e7f5d1657843e7cfeec113649a69eb9597fe10643ab7c72200ab32597b6cef02b134152557874d6a52811edd835f1bf6eef6e30c37a7e18d8e5ce0ffb50bec2d8fb26edec6cae31ba98a17676294fb8b8b9f81a35b02ac5cf2abffb58a66652ebbaa2ab6a00e0a2d1f610d3357b7850437db31957a2e3f47077919d2850d3fc3bf056bbfda91ca29b2a97b0c08885141e6dc6ee15a67052d16519f6804460f5fc565b568c7e32a7abf716c5302ba1501af13eb2fc4ce11be2351131cb381fec658d87606545e3e027932829b91451555b846a5e1ba4828a092ce18909185182fd8808ccd12b445ade7d1870f318f5c9b364f3c46d5743d8e181e7b4d8693c0072cd290f4bbe686a4d6ca52b4d968fb2f1a0fefd4586f307fb6fb1786df93846b156521acd900;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hd0d24d56c39406bc03705c1c8090c9601f266fbeb9e0741e4ff06db62d9f9ddbb00250d5342e356378dec6a7b0005368ed1dbbd7a318493ff49622dea6b5c175a7cc1064877fb55cc46e52860cda81045a2ceb332f8c95944285283fab02b941c7d2f71377919718b9031f2f39d6796768b98b02fbd962220e795b4c58fdf609a7d6755907d8444d4c674c8d88d493ff6488a8c57faf2d47069c102bdada9bda24204e1f2a766fa894abae41cd332c2d827b0e3b098f8e1143a949ae587d0f64e2b70c1cade2362e1f7fa960cba03a5cbe56c9a236382e55c7a1582a74481cdbff429af28b7d523ba8fe86a88baa6a1ec5d3fd7de8014d966f54e031b4238dfb15e342289d6edca25a0bdb152827e75de5c6643686348b1cbbf8ba101c30591507c62b2d84adc1995c4472f603e805320e1e599ab1ae767d5fc3ac6ddd4ca5c7a4f4cff2425eeafd76c95e844b17412329de15812c115cbaaa947d87a7ad34cb8b62da14593f971459b96f8b7abcb519e13dab890cf95388a59d64d20c6c51dc30dd7e04ec446a3d542aa7c9e34f5574f2f8130c40e73bf46d82472c4f2067f512db4502da00da80c2f77cdf6665bf0c4c688055338cf8d16dea4aa84a23cc19ab5c6eb41a6d0654ab388a08e7bad01b2cab00f485eb13cc066d82ce41d74fe999433a5c50a68edba752ce231f44236a195b0ae10c9761518828b9787f9d505443c1ce2e405f9c67ecda1885742cbe576f55e51050d8a5ccc4eefe779bd2c5cafa0a695ac8293ed6d38b98150dec573755cb39c6ce3c463c43b277a6b25c64ed806b3fade6da8ec9141c28b08aecdd62fc157695980ba0fe901e90ba93ba67103f8d23e828c66f275699e5f69248e394761317e2a9ec92d8d55434caa374b9abba4ddb184868b75a7a178da2d7a3947ad6cc190508047d1a588844a2f089d4098e5eaff623513624a337b12cffde30eb4a9ebd170e84177099c438b4abbe7206feab9236e8e5ffdc24d03e2e72b7546396fd26a8e9fd568c0f333be89a392b4b28dbb07df7bb2e3a1fa29864aa4f5a04469ff86c6aba7b0f88505b881b7508c335932abf0edd1bf2dbb971c5fd6a97f5623f1ae4558e7bd2767f485ca48405d02c2d84840efaf9ac9adc2d3464e77d139573b815020f8b7a4bf0e6fdaabc910697b39f607dca22412fb61f0e4b97c8ecc3ea98ffd25805b9335b5f21f0d96f7b36504a15c50da8578d8740946709f3d09ef04070c7690c18e44b6d8befb6360d2b70892f73a85d41f5c4e9514c80d3fa014156ce77d95393a2d7077e5382df251ff1103de296170d4d5719b57ecb97dfbc980881bef51c2395006dcf0805488bba0f481374e27c8ba596b24fcd91a304e687595a5b0128501255c35a57f4e72cb98a0a687983a5373fe15ba00555f49c509531f4239fb140221fb85d44cc02a9876aef0cfa6cba451e1c6a01c495b22f1ecb9adbbf2f5fac169d33ddc5b669a5e7349673aef28374dcbac94823c38a0f04095d46621433ed120dda21d9e7f12a6f54335883b409cfaa299f7dfe2f10ab9dcaea1360879c02e8726304ec49f3cd79fccf87d493a2653f78a81a8b728840bfd35f846c286af02642fe0088d874ad08947eaa0b0e26fb604edc0f938e3aada6f6a0befb1878e04ba8103f90eeb1d5e0f75b53d4e1af98610f37adb73a7666502320ba750b9c133f979ffb0e3c1be176922468f1ac0023e025446c267d18384f038c369bd99b6f2dd000c4b56f722bc42075b7fea6c8cc932c64a85a892668fb2ed334edda5735cbbb0a717ab1f948ae35e31a8e0a6f17518a19c7c37381cbef178454d5e078816c6276e0eb96d2952e18b366bf78751cf53013973c6efd1c22599b32da9c61ff9194bff677f1aae0181197939ce58e05a96a090af3a937be79fe82d16037354fca8df7c2a9a02b814d9e3421931916c2d2d42781565b1bc95224b7643ec2f214fbdcf062afc4e746ad13c8c9c5838aa78407db85c82b0fc0153682c757e06518ddb9cd963a91488a335240953e6cc1e2c7a4d2cce0d00ab4d84dc1b79ce2b7fc91e6f505e373700cfe24210fd03c9c33b28621d5fed0f79ba28dce86b056c4f57c2c7f8f462b18088eabc1ee914db665a2a7769366d2b180ea7a443e86549259e53afb97ae727f0e132560649578ae2ef4bc395af435c14f233465e28e88777cc7107662826cb90d2d8a0651727036b16d1d04180c112edd3670b0c72071bc4d341e5be48faf0184657c28d7f06222796cae459964462820ac679559e7bee45b01dee29680aacf8534854059eaed62853bc557ffe7231fc7203b284e1f5ce969f0e080c7b711db73b518cf18ea47b3c447d6144267f41625fa8e0847250f5bb78d39750904926ac1405cb48c722952bc1b7bf23e52705414263bf426e5b3aa9d03380baba3260909dcb50b3da3b80f11d16970463a910b398cae0aef6461f0cfb81c6417b040444a8a238550daaeccaf0c362148af5fa1677b661ad1608a4474cbabc10ddf5e5d725f7625678869b95cec0d03e7ae3e9fa3e0306530f90a37dd1abc3173fcb2382b764a6dcb02da34c65ecdd02e556c6001f43f274401295d7d45eaac0294993b540c5ac56a90874d44ed2b56d6224d3390869bf93090b7c2b7ee4fa46a2e5e3fa210fc958fef8a1810064a9dcee4c6e9f7f5165274ecd4c75eb0edc362bfe696a72547c5f9311249d64f3d36fbaa283617969d719c973f28fa6012465c465e5fdf5d96a8b7db078628e136883dddc371c87b338a2905754d82f0fb7d56f6173858ed85f631366ab3de7ba3e58ede81bf47a3773cfd8bc7eed8062cb11b2da851c3efd852b7f147cad8e33fcd89ffc7c3333fe4b5d7f34812710977b273d0e0af66;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h50815e36e090e46e5ad5f59f3153b3292418de68a6a160888acb381cc30eb2fffbc91c563d7bf06fdd3902e8d0276cec4e59eecd99aaeec6c503eebd166d99b53e2f01dcce83585eeab6a9d0e3629b7c1ba8e1277e452350aaeb8bb35d6489c35b8ae1c9498eccf5f2bbfa3f1b7135f75d260263cba761b80500643e9e41ced47e7d5ff2afd5caac6df29a22488bad8a0bf6bb0e17adaf714fe25fa90e729eb19c7ed4772258f9db3f4794e6610d9788f5941029c1ef1027611e6782abe8d4091c11132f12e12cdd2d95d786db885887d4f15efe594303c0c7a638bb54fac92a0e0e38af87e05b9a6166dbbced02cb37d01eadcf1cef2ac462d0b7965bc6186a2415af78d9bbaa80a7ea7850016fdd5572cdad45e386c9ef9832567152561149e3b4b8d0c687c1b61c62b0e20eae93bfd04301c38e146b65270d0c06cc30d28b1817705660e93879247cfb16f6596461302fd9d82f3f289d25e3ab2da4a2d591d35d38b9e9bf7fbc7f2facf712cab74324899c20a2d4640f98f449f3bc5d9d44f2c61a62c569924ca1fdbedbe968bfbf6122cee75445a77f979cba20d81c1b50193b02056fd96f7f225c9b348f259cf6df9128eacc161949c6e547f96740f1125061d0a5eafd88ff6a95800a9f765c3d38cd5dc83a999832fe784eafb502a61e33f66f3f347d64d71d19123828df8f56be337f175519f2527797ec52a5ce230ccc98a48b24aacbcf65ef2d6bbb5e6490351b3f2cac0d0d683ee5919617cac07f45e494310230585ea7ebf008bfcf3a8fe7ba3b5d3f2365b67e6d83fa87f3654d55afe871261dec723ee44b7c9f9cfb50d55a0894c99324e1dd41c87fc9e1de6d3af01983ffdb2a1ffde4d8bdfcb92f02f6b06cd55de381b00761d1baec04ebaf0135a2735820ac57fb3d570e3d7890eb038770c7cd68dce051cc8902eb3507b33f87bd1287f72aa31967d79c13a37ab5d70e087f3c4c0e0c904fa4b89911107253afd2817f62534fc9eb45de65599c81925faeed89a09c2c6be81bb09872017f5c8c81b35cccc41ef9a532b33bbad71e896bae4438548e1fa7fd01850354f13d9ba977375729e41ea60710942c20120a2a147f602d276f52c65e72158a90202fec1a0ef2f386bad92c46ab9e3c02e38b4ebab3141ea98aa44a6284e51588c7cec69e83d193183a4e82583c1698a78f2ad73c591a6dba87716c89c35218428342a42e2bc11350896dcc64007a1d29778e0d328b24d0a98d0c405b0cab33ea3403f2dc80796389549c48c70fee98983059fe88dda9423be955cc9bc8b5d9425594cc7486cee469d3dbc90e04a4c1caa63c52a0f41e0713bb6422aa21b6d7ba33c760fb1b460e4957f445bb217aadc2e1576da44ec7ed86a7bad9e34fe479b671f0e47e01704f5a5cfd5054aef29646e41c570d2203da8d7a9727528991d9b33db43bd7b3cb5ac51ddcd423aa55ae7c08d779adc78f8c28604f0a139b53c50806e321c5894757c699686375aec748fcb6497eff67c46bdb3704642c34824ce4d25d9025f31f6b432ceff55c97352a498effc6a1d9bfb67c9e30b303954cf29c227ff6d94926d820d1c8a9b6ad34d8f5d118e3ce9e44406478c5410b96040798d9d7168f6ad2f901aaba45a001db66dca1e8394973c1a428cb6ef49b8ed3677e226d17366124a611bdb2b4de82529339e4a88e2fd177226a87cc3151b5e3ed012055be590fb4dd0743e8d1ddad605a87ec75be148d494d59267257b324309624ee4659496897e6bbf7477a440c79ab0d09c5d144aef3e0e5d84b1e49cdea8b85f2e220e82b5c526010fb7c4be1b4d91e4ad491aa47a170bf76cd14c427c4eb19fed8222c77a1d3450b1d8a617e9806fc2486fabc92c0f3db199cb113cfb8f8e7cd8d987b289238b43a8b9b19f52c8f679c21679cd55769f648a207da12037988fac0e90a2d72afbdd411bd7aef3bc377943a0eb08b8fc6562a02a226d23cecb5038f0858cd3d51babfca96c1d380bcf4485e61ca5f520bdb74e7c74cd2c438adec1d86e5d7e2095a30c4237476184e00f1a60249e021f0e6f74ee6f984a94fc97a24750e08d0a103728996602173ace3ef86660f913bde09f4e56ef7b0e5303f668e8fb1b46c9609b910fb20866731fa9cfc52aa1d277321c15315cda472f589dfe17b5881e8e6e983b3809b68750a7967711b3f2bf9c5bc4da828771cf0e6d6cea8a46acc79881474cd62111a62ef20e1b72984f0901d95c25ce9c52a852aab15f449f5b66537adfc3174feba3df802e7a252e5a2ea3c45927bee52a05f98521e29733b6964b6f6ddff75a71099217d8ae5ba6acec0119035c0ea4fd37a481f706e056bc4846b8f51092bfa9ab7008f9c71a5eb18502ff55f0e2f63c9b74a05e016e3e748b8de08c67be97aa259655b903381af55eb0b238dd8c86f092b60f3753e180af6a0eab552a69e38368a873bdf7ef6de7c846982322220825760f4cdcb3df4fe1c6b591380f5ca8ccd4d18269b76c8ba02e6087a550d2560b1341b5358588777c038336eb0b460b85f7b30cf6cbd5fcb104bf082acf46fcd9412e02e4ae1ac7fd7278d286a4777046d6d6a85e0cbcf998193080076c4c04f3e5fb6505cf18a7eff993db12ec60bc7c643890a433089f41d803aab8e38465782d8652c90a7f9694ce45d3f98dfc2665f74caa4cbba814bc5ee7ae067767cc9508ab561d703e0dd4d4330751e8ad95b44ece30665088a456cdd7d4aaeccb3d283ebb6f67aaa4bb4c93638eb98f6f13692d56e655ea443297812f6996b9e6fa0ae4c46ed1f14811554ad702cf39b69dff3f52b2ca8f1a89612d372f70dc91bdb9b230d7d017ba08ba0651dd2e1af802af4748da7c8e305d61ab798a5cb2901410e6afa1f625f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h2e2908d0d11fb4566a17c28fbe10c389349a4d4f97cbfaff164eaba6246e103dfc7436aa3b5bcd58dbe715c48fc60ae1bc87f6d65b9e95e1e00400ab6257252281ef49c1361f9b677659dcea59397aa20bf051a765afb9a74a1e4e43cb4fcc104baa3f8482cb01c50fac784242dfa002b908bfef3af2b1bc69a625e551841c4721d073ee621c8d20cfb620ef8c9aeb5a10df1c0502d722eae96c16631dcf01af25992a9cea44cfee62418f55597216be5a4eea0af01b04164a7a0e054a3d270789f4d2516a923d7a0b9117c07a4ce285b639acf276df2cae492202e18cf36111aa86bcb001600f8d298df46344f63f752954e161fc54e32be266fb5cca2a83eed3dc392f330646bcebe24720ef81d526006fbbcd20a462c82acf6ffcdfd756d90b95f2cdb98760150342cb22103ebb6a234175589e5808a73920325e560df0eda2d041bd170cdc5acbbb5e3afb26941d400354ace526be6783158cd7999df8a9517022f00ef9dfcf57e726b554f215c4130037961d07f44b973ec5f2240c67268139686f51ad8ca726c3037ed96ba62fd74dee7f4eaa9635bcbb7948f0d3ea542a0fc8b66f49a1003e7c26bf7ec5fc2b637a1e83db24f33708b1be3be7ec6e984d123774683b90c310d6f3482dd4447a94272c6781049fa2bfd18fb376cb0b02db7c32a6f7e416263880eb27d85d4479926b64ec5fd55f97a5c43d1f0d1a68e37ff447281cc74788d1615548f783999959c94aef2e659d1f6d0f20bfa40007e87edcf8185876daa98a7f2befdecf44227d04e39f178c1db0f23147769e0dbef083ef2b0946c5d7d5e200fccbb782be177a69dce8b90fee94baa146e05410e9c93569f7e4675d56c5707239c3bb19ca75787810d05927fc848f537d12339bb244b7fe0f94d0fa060a3a81d06171f38f1379742796c82bc1759a3215234bcf3d4088a60747397d34cca919c9897068a62664f22a10f928b5aaed6a510481b0a12559463657b7d3e6b8e8ceb1bc6559a9cbdf9d534d563488e6eaa76a6404d30a8a7cf082f1b143a88a3893b36e0b78e015e9ec322486b280b33961d35cc995d248266be7e1d1925d49ce241a1b49c1bdfc622e2e8791964706767604012689044a987fdb3c8564a4283da3d1c5df574af20472540b5c7fcdfa6f363a4243573c35f05e01b13f7b562dff40513c6ba21f4360a70f697ef372a79e74ea1b13c3d7cef2f9e0079f264ffede70f81b3a3860ef12948ee832e91457630dc06adeca7ddce00c1816b90c7cc39b5cb239f0d44106896a33e3adadc936e4d1c950ae0c7a34524d5b27ccc3bd7155a0374d2f4456beb5aa2b82b3f44ea158452eacdb46381976492464bae1ba9f30e6870411f1d8dd85b85a382714ca2f07fd1521dc1c2f1d085c6371d353e9a5a786a99e3f3c113f0428d6b26fe1a7bccaa19af46da4cff4a30f953408973030245d7cc7ba4b76310fceed05640065463c8168e6280bf45b37d9997b18a49139afafa7359dcd47977b0cedbfc86cc38177a81af511bdfa144946ab5734b990002f5cc53bb8a3fbfc2646bad1c766f862922bb073d70a8557496c21d8d1309576aa9ea69ec4c940922d2212eb618223d9bccad155e4e9bee5a1027e10b0569c0e2459dd3da1ac386f75cbc1945acd90dec7cffcbe9e3b4e8a80d208b77c06a3f362b3e2eb3bb67ba9c36615dc448f60d0dc7188afc0edff5eea0b054be97ac5c7e0d848942660e82ca6a6f0c4e952ab2e4820e07fbb9f93816aeb04dc7326d3696b55879f45b76680ded9ea422fc88a0de9957581b7759a45b54b7d9455205ce173a42082fbbd00b024f70ceec4697f6f80d59f0469c43ad4ea030b5ea98d8a6604f9bc91ffead8bee71b4074080ccf8f5763fcde34186a2aef06a2143a153bef9e4430a8ad908c4a756097a9127c494c7cd03ecd19a3d4297a8242f5e56a1d91cb9f5933ac704325abec41c601613e3ff973a91261055a845846d19d7a46826d53098a3738b9d23c0815bca1e40750e4c061f29b7591dcf3c5f83e62c5239caa3592ac68d01ddf2f758d7610110cfd8da73fc042956d9d3612a9e836161840d5dbcbd1d248f768ad94a212a0c40c66575b64ac91bcc757ada6a67d932874f7a756926cc27730ab10bbf1327e6f6a66575774b362af392fc490ab54154f7d18ad1b178757845d80b1a326f60607ee71315b8f335353b8609444361904a20dcae7c02fdae66fb483451b05073ec8594f9102e76c2ca40af88bfe732eae6dd7faf98c3a7660f322ce6d6139935a55075536381a9d2fab294af98cba02e34975b899c2fe5333723005fb549d35edf1b8ab10da1d13d7b9afdd8f97577d79446cdd28a147da57918c5b03020d8164f3d758bf2bfa176646205b863852a51dc7f29d4f84b32a1ff884fba55dba7371403c60809a0771dbf560593b62b0124ab959bf41c8ce27237544d9cb134640aaa5eadaec5cc2286a3bd61a2fa21daa5c7151b0f7eb7e6410832125023fd7804d4eab7e710a3e574154b631600f8b65d3db288194ec786e0c27977047baf2e8e6eb45dd300b689973d13961cbf317a82dd5118f787c95a774479adfa186d0206d01a965d7d9dde967e3be67752f197760d86f6277588a50e11752997194c905c46a374bac40bff05c3a7b5799da2ebe10e9179042137d838d469f648a507835f4a49866b4f16d1f6283a1d9721290c073ef46ba5dc3af2944d59be693a4830f1769362194deef0775f1011d4aa7b49a745810999ec1f1831f330c19e2309efb7e24f0fb6b8197aa48a0485bb050418d4b12c99362b6ecac84389807e0002d6ca4e697f556ed7ac687fbc51d58c9b4c5a84be488520f3049b36f616f24caf68d499c43a158f07c8392b8c45a28;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h412e3fd70214ab6a824a260557f1e56be395ec7d6313198616da05e9cb20747e6974218f796279255974cb3a04edc4452c38393bbb822dc6548f319d4f3e9a5ab7b6976c592b8a1d1aad3d6228873f86e5890c3d72600df1eec4466e076a5b0e2c1c6d092789b910f9622efcd10b73a13dc54da1147490c85c18c7c54a01e88856c642e15ee7d9c2c5cbe46a909116dc61035b706318c869192f540b87b66451e4a697bdec7102dad04a25fc919f603b017a53453c7a0263ee4607cbc5fba2bf68a2c68b1965d7af454625d9ad8d0e117f3efe6dfdd109416f879dad5ddf1f8261466da029d2806116b66091e45ab3f95d0d0d5c00e6ef8ea7f6cc67e5d56afc345947cf527925a9bbb582002e0d2e126b7729df3f89b63b037f08b138ce0be4a2499e3db6d8c246b5a705033fef7a392f3571620b6b08bceff023954ed1744e381e6eba747f8a0487a9c65a7f0e21c0b21d0b0148ba6b29d77dae690d4bcb0de7529a15f00766e128631d3d9b312aaa6b5d6839eced2929ea9610a50d267237cd6cc1d96cba59962c45382b5ed9391681651bad7b848d7bed040bc2c013b4617250e32bd5fc5a528d9f25a4a81f08dc515c8d4e6a1432e6075c7c6b06ff7b42d2360c06ba744b0565a6a65a5f1957eb21d77a288542613dd50e80ebcde81aaaac7b8ee61752e9392dcf0004bae0606b15954614c4c3dc0427ba639f0d31edf98aa6612f4b07e75390f424a85aca1d0d0924e938410b3594b0c5fe6521de42fab6ff764b2ba9eaabc7524970c630ec58703078eb981de4b3ff2c363cde4d6abfc9870dd71e41e041a3d00c63205b1d051ba68b2be1295ee8d74ec671acdf647efd696811daa67847fe6ecb83bb30289b005a4fe7c5075fa94db3f23fea23a09cc8b024800aac449a4ac691b5dfc625e7109813414442ac98c01cd32dc0855ef056d96e266c17bf0306059b595e2fb17dce30b1daf3e40e056f80e64b670b5a39d717c4ad25a79075344100b2a0dc94fd5c8c8f382e93cfae53ff3c41ec71998db94a922517aa06ee342868d1e791005a0d216f37d7b3bdd288706062f7eb8f8d38940186bbe22be49fa20ebdfde06d8bfc8ecd84aac985afac01d19ad854577dc520ad58a56290d72eb94ec1ece70025e1ac3c2aa1ef6eca3815392448b37d0d9b36538c95d5ae5df9c3fd98bc2d57ce876e45c7b69e36ef13b4e26c1bad24bfc6a5eba0ab5f95e33e41ae3c57cfd5d9320a857b76ca04133e8911ad35b003ba63f091ddb36745a5bd63e092beb63e5ce74149cad303bb4544b71b87804110ae09172472e520d10cb73ea4c7f7447e32e0f89a1ffa5daef3519d69ae43224875bc8e4e5122e5cbc64663451978098a3640e0b861c9a0ab66ae934405d575d87350c0de1cd48fef283b97ef7d230f454a876e1ecaf6614edee8e2c45a21b00705d451b77409492bdc4a89353fb9bc6896d77da4dba44eb146d32dbfb31b224160a0df4cf4ea87211e29a9b32cb26f1a95249dc51c91e2d0839ef0322fb8d91638b2ccfaaee24faeb2b4b30892be931aea6500975d37e5e97fd2b1a0ddae2b5e3d76c25cbc6a3a871b2a61e48d6684d550365f1e48b18f71fced996cc484c0035d36674498dd6ea87f870c79da169a3ef82e6e2956e4c6fd35868a2b28aa79edac5e111fa895e228d7bbb0f41a8a2473fda679a341841ca03461cc723a688363a5b094298f81f692f67089d3f683086abdb5bf88f0c6ff937edb9a6856f77c04670d5b08f0b62b9a70458e190cdc1aa8e29f55ff658e33b2857b309ce739fbc3a61e2b73062ce953ef42b7cec0eb4174410a6fdb1216c59e4f6043ac674d8a97ceec3d388651c16970c0cf743f1f67d26362bb1c84220b48d1eadfe53ae0451d8f8ad342e1901bf91e7ef14bc2e103d63ddb31eb3d2ba88c6940550bd4d5e7f8a3bd91a0c5bc6dc76d0d1bda664f0f0981a0dabb60cca04c507bd7c58e7a3da253adf1e39b0abe7dc801b253c9503bb487244f291fd0241c3846d32078b5a0f4e6ec1d9165fa2f8e107d00da620f27af76d43adf154dfa4af942a99a426b3d9c919a34e52b82637c71602c2361cab6fafbe97a39bcd4c87317b516071535cc0fc61a5b3453ac1b3f8d610ef8751f19387b660a1e005e1bd554d87d7c3b8e4c961bbfef6b32fedef7d84a9e92dda3101d5b04e5553e4b7faddfd9f942e439eb23e570c195398fba164b935d13f9c8f8c536eb0330379d0c3b061ff9b8525ade941e3f983f9ba6f2d1046e95cc484fb00ef7430760f46793dcff54033da992f4e665dc549a55c2aa77549113a2a00fab0284058efa3686565a1cb10dca31a375bd9371a0bc502f2ce859cba6d3dad2b06aaa9d9298571ee03a1f4f700b6bbc3bcb777aa8db40aee57687f58457f3ec1805431243d23cc76887707e766089e865644c8ddd8c457cddd107a63ce8e387a2f0f67ef7de79b054d6bbe578500604f33a6f2fdaee9f919ecf16dc00a4f370dfdff5668f56458d2a6c2ad50ac75acbdb0b064a2bf5b583e5239de5405f9ecba983ace45276fc017bb74613604dcf81d85a50c244483e21fa489307a6aef3331f36fc8541d700570b387bd915b6246ef39415650e52b5ba55a31986b41be9489f958a9b11024ce42d89db415a7ed781afff7a1b9a5ea730860ae7a542f49c20b783d58dad0e078ff4ee6919ad527c87bbf070c3421a56e5575a8672d1672c62572545aac6b7c9f4b8bda2c3a93f6a706f10ff8187a9b13bf89e62acbc8a8926f767615ca2394659d676728f49d8d5ff0a545dba00ee824ac8c6df5e1d47aeba141fa3ab24a042c306710d316766e6e113bdaa4ecd07722b8c35acdff958f3b5c8fb7469a35d633abba48e180728e186a48;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha0ae730d74862b2f2ec0938ef50734193019e724707d5171e55c9a946428dd5322224b9d3d281e4e28bd0a89afee175e56df5178737357f100bbde1e779fed8a6499e24d68ff145ad1f71835b7cd39dc69fc260e085b10cff39958d218091740ef08793c4fe34b53387d2642cf6c53433a5219dd25c77deea57afbe3fd0b7abad18ef7febf2abd8fcfa9e2c60fd90746797bb81d8d5a3e54066de3a5a1d5997d94193d703337833213335b94f757288a669c8585a07b683e9961dbfb34c947c77e4bf8df9101048b3141e0ca848ceb225330be71558f499213b8e8ccab348678040f06d3ff415cbb5c6afb9a124dad3d9afeee8d5bd2e1fb2936cd682794797c4f93dac5168bcc7926d3dc006eece5330f60911f6181049fde84f4f6f877288b918cc03bc639aedf6bdf92b575c3cfd600a005211d10fd96b63a3b8d2e36e51e91bdaeb2fdfcefe9b2e36e69dd75b3be29b287ac4ca15d8f41eb271676fb350307140773a64e03cd9ef1bcee5184ef99ac8e8942e896b278286da1bbb6327a13889fc4bae3e6275ace195e7e6f526e1c92b6e97bbf277ce777a01dd6d0203abfdbd7a5f17baeb85d98f204e83ea908dfea4f2371f510455e10efb08fddb98ab8a04e10d88076da4b4308c1c7e7cb8b5677829db03e11293c49bfc624e2124f7a071a8f0dab4e7ad1db10cbb756bd80d6b758404c46f3aeb479feae58e05534e45f03cb2c8a6258d97e2f4f986e7fc0054fe0a328701064fce6fe79746f7e2f8cae58770755a49d6cd89f7f017c46e8c3313bf19803c06c4f3a6e8e5311fa56cba872954340b3616b642455b6d6118c0c529c51e823cec99f3c82abe8b49261528ba29adbd2f92ead1a906c8c068d8d3a81f07ab2efb1aa2494df2cb4f69a3bfee7fb72c79cda9cdae154f34755e3b4b83c440cf9376d28f6a8a91081501f5f9e7bcdf3b761d72e51dce038eb974035a513a21094d62c6e24a8ff23bc315cfcefa30b0250890b3c5565a1080a8f577b8535cbca253e76ceea91e0de37426574e81faa29a52f5b1df0f0fc9e53ef06b3c0fb63c348ae659c89fc8b98c1db3354cb87661314e855538e7d4ca53e46a846e398abdd1ed9de177df8034be1dab514befcf3e85c525363272f28e96d7f5fa43fdc66955dac246b4ac05384c56d782bee0d2328f89051b6584ecd841c56b5cbf8bd71f28c7bf6aa22828fa00ffbe1fe5f136cf90f66dec2c8d92a50590a7bd89025a74772c3c7e5f96718f5e09d503696edde4852b21b5d9a8f0be9b7c946b6d10b902f07b98409aad448772ceaf7d76083a8a4fac1e18616b84ff508a989e6b8779afebc7a81f946b32e4ffc383ee683eef1a29bc9cd7c3fb7ff3b6ccbc05489dd7d0f0bcf29314243689b1d926190ef99a43ef9b00ad2c2548f0ac869a1219916d1866e88b24876bf7ea757f0e9913fa4706fa586787390387386dc6aa02833ba78bec02c8957c0b58645b948227e815b41e9c5366a359acfdb442a581cd816d006dde6586dd3b54d6c1e5de5e0cf2ae65a2379d61e7e898402f1c993d200bd467d7576b5062c6a379faa84035f20234036bce6520087a50275e17f6027bac7af57724f4832b52ee92342deffe9eca2625f6dd7f4d5b46ec291b468b954a3b9cf7eaac82ef4e34dd336ff6330604d3dc3ce4b4d60de8ef716a4d998aa29cbbe3ac3ef6e92e8a53e946196ed9106c0574158f26f4b9f30dbaaa91ecb7e00dc7b4225134682b8318c0dee578442d21b2d504561c797f1287820939815422ea0e50af1a0f51e20e664361e625380221344d5e36f17b7cd9e79697f9aa73c38086efa08ca3b1a09dc13e2b16999686e80201f3fa37a032494d16eaab7232cdb34cb2639fb4063360e090b5234dcd30c6423be7c21ca370086db05e9714a7ad71a190027ecccd1fc50c3eb7185304b275acdc2268ae56d0445304f40aba6a4be589f93be95637138d858645409468c918152facfb35eada9d06c1021876b5c52ab7cf9a29e6e127cec957d728b4a08462a5ec2569f53b4304a2eebecc767a4a43e6f2545a738af37840b6a0e811ec930adbcc9ab1855374aec3fd26aa57069708a68167fbca5f9119f7d14d3a89de72647f7b89d64d7339b97e732fe2a4b24a45afab57bc93960c5beeb43a099e1c4c33c4f5f91f68439de5630f8be5dd1ddc4eb8efc5e2fac2597a46820994bcfd6a227748d1e9f1797584aad3fb16829b8185d702b75c99170a78d92ca171e1c560a950e31d176e748caafa973b429ff5cd8be9f0471640296d2c1566981a0349333a747424bb309ef4c3ad42245157abf1932b32a26c178ac960a99e6fdf4b79cf7f78cbf1f3dc827fd832a8b1c57a6d6020cc6674b25e608d44eb24314fbaec80eccdc346566bdfea8660570fac1f975382540bc87225671be4097f9898cbe72fcce6ba2c90b34495a58ad804776b720a7ba176cca576e270994f3a58a42785db41dd457c976ee578b92f20fe2925e61534f8a2dd3e9910240e5beef8d8a63beb9ed6604b0f26dfc86cf19bdc01ee00240ede071af9ce39315e3b5185c2bcb925740c9b1c38ce940acdfa116246b2337cf8ed98bc1b04152d55764d4646ba6f64f4dc43e0e29d83917e4adc861e8970dcd710a3ae9178effd6564e6a586eeafa26319fc61c90c0bab0b79c3e4df0322a8fbd53a7e3f6c784df9234527f85198d7690e870ec671800972a1643c84506dfbf2ce84cfd38593ddf0f3398d009a38cbd1e7bd900d49f196df4ec07d3c547a72b35c0186ebb51f5a98f233714b6ea150c1a0011a41824b22e502b36ed7a3749e5e0d49b3cfb5b47ccc33f7bfc93241c30cde80cabf7b32741ff6fd7dd24422f8a6bbc4f56d7a8b9e72f5dfe889b0f71fb1b12;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf35f3df8078caf2def8e7ee1d2aef8541b0ec2a213f8a14f46ef1c5522c0d2ca9c35d50bbdd6dd0ea5c2528747dc2796a6b79872fe602b1c0d30fbc0046e8cf35768044eb27e1461d4710ac591e37d086a93237e8b64934125aeed7141205c7d2bdd8a35e93abeb93a5bb04a069bb1d7801a5141f961f13c550bf1c24961075e6ad9093ec5da45ee0da06846b2fa08e3977175e91aee17963f70535d46d4501a5c495d3ecf467e74155855f12a6ed3dfcb351a64b00b179109f4aac1d8a6a58c46cab47877adfb3919fdc9ed5ac5eb3f9b0a560fe292a90aaafa7721df0b7a4aa22a9c430f53361f73caa4bd3a7da95aec5bf4d17ddbd003aac0fd8664599cdc64a8aa5af63076d84cbbb34580602ca61ffc4c2d6e2843abfeffc59649230734592dffcee5d686194240c972a25acdf4e6b5feaa43a49a39c6f411274147c86b21403616264e0a978a9df3ee9be04e7c594e227813bb41b315ae104f2070b73c9d2fdec0d97c5dee1f988582d27f038e9d5b47c76e847b52b61913157cb7f6230e7fbdeb9bd2489eeeb64e21148822e9b9e5e4a99c4cb9648fd7a0dde4105d8fc9118f43ebf909bf585b0de3dd6ff16a3baba0ae1d5c174cdd1c2e02a2c50d1c130948b4f4f014688ba8028e4f7091db32907fc1ee5ec47e9f08706d70dd4d2fc07a1bcb6fe5df9fa9ea94d61dfd6b98e1dea27107b38a6268efb6f43384acb974377ba7024118e806a3fde9d53ab408c7b5271485786097d91e538e386ad76cce6b5b4ea9dbe1383900372b251b4819d9bf53db06cf4dd409a574ce5bb72a8de4a2c495c82c67c0023f1fc1d26918d051c10bf4f0ccefa5a3fa9438ff072f6721c697fae12c2f69ed68b1ed49b8c937c395b078472cefaf8d213beba2c022667ba01a15697b9b8d91f3226a3939c81540a58398d38a5a2ea5571c7f9aac66019e5760730b36bae9c35ea477251d6b9b45df26c2ddd1fb237fb1b7cceb5a9d94f28409ad43c47b919ad0b927d4b38402a74b80e143ac385e62bf840800f6b3ee2b3c880254e336cebc7a6904c50ea4f754283ad81ba03ffaa03ff3e04beec973d11c57c8d423e15b340dbbcf6a26a60da5b7af03c8d8e95f2bb29994911ad5ab799df881e8024fca5f17ef3726929d3e7c8aeabf6d14eb043de50ed7277d32fdfe6e2502eae27215692e58185603e0ee18e56f670688e54e94b4e0a1f57853a5cef8882ab9b6810a06f12de6bea16a41fa5f39b4b3e8e543f5e97777c8a1a6826092c2bbfbb693b6354b4a3e72eb769904ccb1af29a5564883d6b0c0a5c55370e6dc7e067378a4e4f0b7adfd0c43a40007fc7d8f9f7400c0de4617904a646127a498454373c25580c265dfd81bc17d14a68a2f9bb5b912765d77560bf3664e1a3b1be4e9911f3c31a4719ffaee6105229d4e8640a3b1dba774be0a84caeea8a6b8fc380eb8a49bff9d5f51dd0f0d06afa71c50290cad03048478c1a962b2b1cf49b1351b2ba06a16001377081a2223da383f1e5e64ff5e1d6d608ff10ea3f584cf266d969c3fa4bd6854c283647af2dfc1e7110953561ca095d88ca88aad3492b19eb1c8052d3b7644c25c554ff18ce6321e324f26cc4e5c6e83e08d884b71681dc0d5e61e4463d3f5d485cd5caebaa8d92f396c6e303d26d272899e253a90d90fef4215b37c4c114d916b62986078e48a602c6b8d806e4d56e4f555ab12794c4f1f9daa7060eac27c6ad8c9137e8c41a5959813bc1b5e5af3f33a83b5627f4e3612ef9bbf733571a8672e7763a7088e1f673e65706b018479591ddbf87f99247deb2c359d0c12fa8ff9b78bca1697b907eea07e9d243978fc92aa3cfacbb8bfde78506a82d0a1fd9743eeaa018928de915d6c0bbdb4f420138e876ab941c1690ea2429ee85d57a0b92df21018256e6d68bc6daeea10ceeeefc71ea72c45ccd45050d164bba4a84447300e24dbe22af1ffc40798b007bd044a0ada1ba7dc9ed41ca97e9c972a6e21c11d1361132d138c0fc178d97727acede4d92f6d1c5140b2ec0655ae0b91a13976421bb61c155d685b5f57ec43ffcbf857caf16f12315b25ad869ad575eaa1ba14eedfcb915be316d2af3494acefe1f6348d43e881d5a3af11dd0d7a889039412fb3806518229943cd4200425f50a3a14de714486f3bef8675848f1ef77e133e2632c12c3b27dc8a6554c675658927a9cb186fd1a47f68a7198771e4c79848a6d2a29a4ae5cd2cf05ae1c2fe6ad83bdc1c5d80fcac1d2d94ea83fd207fea74868752f7d72cc958edbd36cc21aa9cd67e0ba3457f4432e16e299ad5c169f1f412abb3cb5da1782c062a20764340a4ec1bb11614ff07a206623a4f2863d76aae8f15195e741b3e0507e4ab8678d02204a9eb9bf59563ca4d65988ea6de06a15abc91d81cd0112369199eb72b29abfabb4991c7478c3434929b0ed7856d46cb307dd3573e41990f63e1e37c75bca90c30d1b57016ef9b6aeb1d68538704421cc66e688990f79144050a7029465829077a67b19e3d45757e61545a0536ee3efa76a0c8b3dec48b782562bc3ae2fdd336a3a93b64459eda1bf220e096776d6df0c41d4e3d597ba3cb393981a4f2cf425858e3a603d4d0396de5989fbe1e37956f96471188916a807807f66e709330396980d45e8b2fc52a97971454b86a68d8979d6a6b306bc98ba52edad36dc6c3b6754a43018b956da98c4e6630e25ff0700e8b3477daeeff55c0f583d4c9d250c9d59066a11450342cb19c0e6a9eb97d0286a833611dceda18b375e00eab06f49cbf8a74feb07e2ffe3341a0b7ddbaab70211fb1856dad7744ee5e3fa6ffbae5c860bbf3db9758f2f2190871ea93c12203786a5d82d7fd5c67a78eaadefc6f95d5efaf4b8e56f8be8bc1efd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h4ac6fa1a5685d206367b58d202ee11d2a905dc41d38e167ea0304cc99ab149e7efadbcb94112a50e547eb3b5ceee295deac382efcbe4c8b776ca00e25247f5c78285d5945a9e6ec809c6eed6407aead3db440da8bca5c23b23be2a3098b7ed38ffa93e7478efbe6207a181dca3d0519bc9a60a8997bdfaea267d80232546ef0f8507a5bff7b342851655755a9941619c18b589680635364061fa54adaaa5e91cd423524d7666af1f845652ec16cc75ae8abfe3aa897f70031c26a063bb3d5df82e41259f3dcf865e33b9209f8c39c66889191491f696d4a1d04528a98e3e116855c44048be5c491673a4a9ca236d1c670ce35c6c16ff7895dd31e0af2c81ed97d94bf0c531a26c8e6b477c7c4e4903c37980f4bb88e612a635d2739dfe9b1420f45cce96bca73e76895a3da85778b62507ef891e1212b59611a1d1e58e8555b98754d30e9fccd3294a6a6ee2013b34216b09b32f65e172512bdd6b654fa754acb353a82cc0ee4917bd9ade45ce6119549227bfc271f38fe807f28194b495893af59f4080111288a5b3512192c36abf4d67f40bd2076243d63f8c10f4f928d6adad25e1c4f5a26c94f3988117707ff27a444790136ceab4b43f963514fb814c337a3b743176f7f175d52f097da5e706662113338d284c0f87e8e8ab7e13b00feb3a989188ad5f80095e3a7087b69f135d880d7962203048231c9e1671979c1e4e137d67f44876031853e716fa7c6446b63723e83867d78d7081c2d4dc95ed0ef8d1f487042da56a7145b8baf52177327b14a8adf00bec4f71a488fac33887d85012e1fccaa9700e215f85a63f58117a4f5303aa891412939776b280f106c1a5e77b3a746739bd5efc8905ed206b6b2064bb47be39af5248d3c583ed6f7480b8084881145d3736be85f6f74604e37e30e5229dc6ad3278052d4921c75fd7d6e51640d21a17c64895e8fbc570ee358eddce73b5aeccd7ae99f667c5a92e5eda7875ca37df7ec8a9ba1fa8daccce6e952a1bbecb067cc8b103238daf6fbdce1fbdbd447da8465e319a0d81045b34d665a1af039dab639a977d17d5db83abdbf4b4d07034757c1ba627fa9750018956f63757e0995e8a74b7447708b7fd5673739daa51cafa8b18a9c5088aaf8b5d45d04fbe50aba05316be17a7116a64913bcc2a70cf02de7c87927a85cf520e499686b77863752530f728075c16cc2eba78280068ed82768f95a73ba5e5a2e7e51ababf2b18f2ae6ecc90db500e739e401c73dac6e550cd6108731913a7130edfd0725eb7e5a25c2adbe834b3d4f7ad509d4a5de73542dc0d55ea08fcefb05d043fcf37c2bf38231a1892a5cc782f8e93d17a55b2b7a24293ea09914af311de7878f52e37d59a9525a7c4c49f6c9fdaac1b92d3d80c40efc4b345bdbbbc3cfcf6a508d5b44989c2227f3e24c870e36c1c41977ad8c6c787429f6f82b6f3df4ae4a72a410db2e56373688c51a4107368996f780839a79f71c5161083b89b911816f5427cb2fd14f561c90ebd5db3b6b2364467038b8d5263e42320f8fce338a1af81f8ab7bcdad859cc0cee444fbe7800a96eaae659ae8e01519d419d629235c63fdc1dcee9411af186a3a704005f83fe3acaafc1c65fbf5162f2969f3a5e1d935dce5dadca62ca8d99c80455c1042f3870b720eff8f14f721511d8e2de06764fc7e5f856d3bcd2a07bc407451eb417f7f7aef3d9f34208ffc096eba98b0837ceeba034997ae243c3be60acbd8c43b091b1b247fdc75661c163c5c46f726f0fbc6bc035cceee4c4a9537131645337747a8018ee4f18cc5faa535abd32028e728cb9666afd028376ac79bc553a1de55473cda430c4aabc7211dc2de0a11b237d268aa6d63abd47ddc06e99930bf5b7fad0dbec82c38a04ae8624fa004becef2cb0ee34f044aee48def8b8a7e6c43b324be39d34ae1b6f0eb1221f09f8ba05b0359dc2c470ca0407d30fc1da8b88357cbc9d5265f4dc3f43ac60d76ecc67becbf87787a0f5755af561e149caf92e2d05113279e44bd031392b5dd5d0f133b3f0f4edcd7a07d9cb8e5fd01e21a6f60ac759c441dce9739c148d65ada913569673373c152e08669c6183d832b03a0f113c2b80839e82db8aa0f32531fdc12bfecdfd3f534bd47ddb365337c4f770f496f3d3ae48b2118eb9ff2c81413613670b27504e801ac4f03230a778b80bded79c81f1ea3c79b11dcab09e7179d25b4d9b06b65da98c9d5090954ffde93efd0d731a34f3e6d58b2533428098713a0cc1205607f3f47ef1d05f2470a2900307cfe25fc0fd0ea9d73d0945a293913e3983cb4d5738cb4cf9de2794f049feab86fe26ddf5973df78cad6f785271393b865cd7cb94ac49275f074603990d62e1627d3040ffeffcc12aa9b5e6d846fd79ed09acce50a2b8ea86fc22b6e5aab3402d694cc385623720df18cee1990736d38d5d0a5971287f686b81b9ef2a984835c44b183b70a27dca5ae5dda7c6dcd577b0ba7dab829334f94b98083dee2d9914bfae77e69d2c298f3b0d7eac13b5ea243c9271682e38785347a21174d9ad28fdfff12c059cb664e63535f48981eb03ba449c9c10994e19c5a230c7a4bc31bf25a32a86f946ea6d56e1264474e5d720da927150f9de5fe6ecb27c4a11c3fa040fee44fbf2f5b51e6f78acb35002177bce797dcedda1d2bfda90056dac2c0996c8faacafa0d3070bf1da30a41c2af2c5c31479f40a6fe7a53c9642386cc17c349cf1ea9aeb0da9a7dd89b7824dac02496fa472e88c96575895a4fb5f96bda5aaa35da528800a669bfdb39d51d18e82e4e2ddc9de2b6a7bd75d6c28ca5fd38c4bb4f98b6835d72a5d3d6f7e68eab819defdc94823652cfa3b9cc9842891d33a48899e2337579c000ff62134;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf973fe5bfac7268cb56daa1e35ca8c31ab33ccae55a830ee4cabfacc8c3103ebc00e45d659a62e86bf0caae0cc08d893b87b438ed9014df772086ba5035052add9db608e5e90db84c4fcfa5904768e3124ca2e4652c2372e3b6f3b4a33f379ab73f4c64d73a1a1b931b73a0ccf494a679da1b14e748a00ff6feef9e48f7df851a4f5fcc0b199443fa2fee87fdfff7faabe137b23a98a08dfc2e5750999dece5d3e0c784bb5469571457b5fe9eab9c800152fbce4732c7e835651f7174cb1998e15fb4f282d78b3a6f02b04f8e6411b7a8c77e4fb311a429b4548213bc01b78d45b6993eb88e279ef0188af33af75996e5dd0b4749c3f2a0ff2edf4830a6ed1f133c23f0c78e0b6e64007779def8bcbd67f1325d5910346494ceed678deaf431bf4f82b7d87fd1d0745c25c0c18c1b51ace7e57e956521df1cec0c857f72eaafcc8bed19a38e214d7f37c9d5c2e2cbb5a82110b917bc8464501f12dc940a212f354d995a5b567951ffa040349d4930f8802204f4fd4528597673ce517785540cbc991fd38b5aa722e995bf0d001e07d35460b0229aeba4264f6d2385def127790fc7983b5a92b082dd385677b99d29dc5fc45cc0f7719791f21a06c90c47f6d7daa765fba8846a57543ea6155d5929ee2d8a1f9cae02836a7ca9c533caad65fe844a17284fcde4222825f39aeb0166274048ab401cf57038a86309607c8bc6eac6bf3baccf70702e708b176f4293fe9158659bfbdba33bc1398bd376eabb48a9e858b6232138206819f1ec4c54d9fe7f100ddeb5ef4b5b2509ca3e34811668d4df4e7c08f88821ed72a3261ff0297e491d70f6949595f339e6eb72624ffadd7e29a7ef15d6c4680704d9fff06ea449901dfe3176fef197f52594d67e70123e093a1925fffa477bc327dfc0affaf4b00088232bcfab8b1ed053174b4db0148af7a68fe94b396c6b5be470212f58c1372ec6e4747855c3bf7946e93f5918d574a60bd6ef498cddef02fc770d74103c7d4fe71f02f951b054461136ef319c4214b216a65ab7ceab4d809771c671b8c8131b4b3c492810013f2f29e4ee0f28ac57c32973f4e9c23ab829e23bc76b3d607c14b2de862bb1f0184b969adee75697632173262ad88b9e528caa65ef037271661d15c8f1316c7d924ba30bca2f8921627ec77c211146f85d28d6ac6942197e96da7c24c5c09165d5b26038c3ec73225d5edc86b3b4a205d2d76093ffded181721d16ed7fc791a667d34e7d1b5342cc0504b266dc9e04678650d4af3b92b0a8916d4077bb44ab818c49565a48b07b7f48d4d421312061417f40ebd2a6867f6c4848f752541e5fab468d0ab48416cd279df8353b8cca4480cb0d47e969142b85925c554e359c525021b7313dce21918e1808d998360e93eed619bbd0e445fee9cb24157357d9d2b791943a387a5d83dac5d093cf2867231ec8e894376585fdca9d3674ce979522cf02b459e5a40bd5f1b3b4751c0b02829dea0a3831387672de2475e205357df8ec3855ab5137363ab870cbe70f91be0436a022db3d1f615e1d1bde5fc189d6a27e95a3fdb7a1d908cba1554136b429af9e33cdd3a490e59b10bf3714446ef3e0cac54e225aa202d1de2f3fec0695c0cfc90d3056c0ebb27baf205a6a07fe7e03f5517394ce80a5478fa6b5326a34bb70beff796af3973703ec08a18dd8b154eaa551a4cbc44cff23cfb2bb2509a0e91b51562609c83714edf49cf0003297273ff68d6a1b2bc3d7e1eac0bd0564b64d08203422a39b021d323640b37caa4c29dc07766e9acb7b890f1a8dad6924f5ebcf442f2fd738a4b38e84300a059bb8ee29255e9cd3fab27570d054b64fd7d0bb9264bcbcd8bf15663f2922082e0e2d8a7b520d4ac0cba06f9b69865f77950b246ba3f0adecd97d3743f4714514426d9497b67382c19e794f19e63ca7e16eb36828895219f183a423789f661eeafc466fef15b38818587d51a8aed49a532b959e0049385c58dfa83407be787ccea134c54e3a6074cae216d364c4b842e6296c7f68e1f876e1b25898d151ce61269fe3f8034a6780852c2a55a76dfc362e776f55be0570455c22ac5dd3e98964b1f69567a74026483399941a42124cb0a73aec9c8f43802abd3076d820bfc623f8f043ddaf615a03c6469f494c15db3396f5007314b6bda357edc282a9b10dfbb07b0390aebf92326a0e676f91c9cafa1b1e11eda02ef7e86eccac3e197cb68c7717c9c7f25b8b585249b1fdf95892fea9d9e53b21c23fc7a7aa1737ab1b5eda02b76ef9ef13734e431c0906ae421c387036cedc9e91cd9ac1f7c51c8200652a6c24029ac4300ec2711f216141b4c0f91cc7de55d409d783c4170c676ab797fd31dc280df5b2ec1a4527aacf5c4d7145a8252a0eff3547adb4d8756865be00ea2c8706d65a03480cabf85ce4c761ca94640ae1849d054368840a20b8878611f4fdc117de8663ccb9c6f51796553c3d593fe43c10c6de070f0a444cb94c5ee5d76b31575000df8d5630d1cc509c9c8e6c5e946a9645a56dfd0bebd30b1979b99bdfa6c2b4d6efd195981146a18c15b0052061971198d674e4b5eab9f65d6dca92b0e7d36f620b0d77833e9c331a1d172e0539a5e66bfb2acd568dc041c6c56eb3e20176bb00dab305594feea7b8d800076e7c744cc2424d40058b3b0378157d72508b8dbd3f35975cac81de802317cf90e3fb2d2bb3c86d84157d1caa92981869db939913eb5c1fd8bf8e59e234768dae287fc6e50147a80551a2b399ad4a2021ea2b4de67e15ab6735923e9c44d348cc0c828a83e82f3e5af8bd321464deb3e642f54a53aa5d34f6a278ac5667a7a14715bb6df9af77d3e6b962afeda2cf443d1c032182173898a4ea866bbf663cf5edb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8d983e44dd49e807fa88d225f6fac7faad0e3d035e9adf5f29979987743d83100f3c3b216e1ead65002c5e60ca85bd990281219f6cf3447e2ffa3772df6f1e23531f85b7e43f7244e50f0895cc9e8039f01a50be61aa6efc0696ee09aaf2e6fa223d3138206d0951242f86f073a7755e24cebb89ff8681118f9df15610d595932f7db39d980c4452c8d05fee5d15b953d27d00f92d4330a389750a831e4032b5202a2c27cae7eb87d98663733d1afa15e7536127b143bb30f6d996a3b8345c2fccc2f56c14173dc652ad21f3345939cbddfb6dc1ef05df106c020542e4c6954a27dc9331467ae69cea86c087e70d7af618fc7116302f8b0b577b8647b1ae3a0d25d6d67be46275b4867ceb009287bc4db532cc094488875d56d4d346d0d192be02cbdc8a9f97d31c07925048c75ba11594f61c69fd76ccfe5e903b19dae6515716f2acb39c467cef59064fa7aa1aa3564d85f55c223e9d387f006258221e5b4b243907ea39b9b5903f5bfec95149629bb9b1ed3cb2c3ad6705d96c6b954c924ed5ccdd7c9573e34dbc2a4e41ed5b3b89930d9da0a92921ca8d96b46a880d36bb84fc1d11464b0c6c6c5116c0dd415306ccdf019b3db4dd8de509f69aa2c13847e829ba4f33ecd88ded75cc873a45ff31addd81dca1d549e9060855db79b7e572b186c418e48e6757f98d530d9a5a0ca51523e2370853e23744b58eb60ed28961367a41703318c3957e70ad8f60424d7d0a8c7a4828c11c70e32c535d80ff3d4bf3e74fb117f6ddac1049813eb63b79063ce0d600bbf06c5707c1705881d4856cc501acc328082ea5e38dc2be23cb68fbc986c62d0b2c1a706718f5cf9a4fa74f49f30e4802287c48b68778a898817d65276aaa8b57e6f7ae9250a4ec28b551f58f5905b11c9754d415b8e510094c58f201cae058408dbb3d04469d7fe3d6a46d3644ba5e7708d08e1cff0888671e5eb99d3780feac8893ab0a097a45114ffcf534be9f47dc64179c962ecc136da4623c7375f7464ed1f920c1bc2056ec2752f8a3155013b83e5d80b7df20de3e23a82c87356ad1c136115714923cf3c886285883ad9a1a8ffc1a1d5d15da4a14374b0bf75985db845a3ef2e6346fb128cbc0f7a4ff16eb1fbbb7e0a3903483b3f8e55e667ee90243970309bb25940b3469957fc93ed67604c4cfc01a6c6735de701676540fbcafd52c62c1b6ae0f905638e8b5a90a4b63b5ce4ddd6411f4614ad38b9c518d693644956c5e1d6ac398e2664ccfa65eb772bf9e7670373aaf9a58b462a981e15c78f75c27769328ba8a284ac6fa9d9c03d3587755a82188a33f34088cbcdcc4387d559424183e462e27e1dd4cfad70ff0ca717de402176bf038e9ab53234a89eb1389be2db5e079f36584b2cb1001596830ed9ecf880297845855b3271458f6e20f9f161b955313106b8acd03e88170034cf9863f4a679b8c99418accc508a96dae98b4aa93c07e7f18de274feac2ae1a55a1f1fd764eba4e136536e362cba7d1488be557f203faf9050a047fa2be798b1e5cb3d21ed766759bf230ca8aa1174740d78de013bf9513338a6b54f6565711337f208acb188138decbedc6ec6335b8c1f6c7a885c310dd23e548ba6175f65868485eebcc69ec375965d68950f399d5bfe7f0d9472bb3bfaccb578bcce61f1c354dc50e8852d545ebb10e9784a1533c9885df39bb67a0b74e2ef63d8108148d985b1fce958431823e9f1c3273bdabe602ff362dd1b2f40a950f0cb92e5b7a4ff27fdf0dd75037a6f9c9a52216a0d5180942e891c5405777e4cf1615a6dc1c635a22af2f571a198ef8157dd7cc990c9959fb84421a0ed6635f02377a5bc8621598e79f34fbe129ed50093bbd9f2526d6ee6ca2c1489cf8fd733b27c582b255f8a1dcfe209fe0cf87d37a4fa3cbbedec7436886773dc01715ddd55c3519a1e4126363408a1b903e9a22f45f26ed3e30f25bba93f182e02b7fd37fb783eeb5d23a1aa0f3df1499e84ccb8eded9c15217f81ed33c82379c46b74ee17283dfed160b9b267228c1169bae9f4a21164078ba5a8b354e37a27a1ae50f0aa8cab534c2429b058b2695c73f30ad76c3fb6769f79639884cf8f36f131aa8f980bb529dc3728c5d30a0f29b425f6d645fef6cbd6833730da3a9402189a4d38bef241717a39cb780f7b938be5cbc9b803be85f7c0690549e8714b4d899ed1f5164d0c0aab343c45be9f1ec801f5dd6865eee27510231cc03a85ff805a697cdbf6f62052eff48ddab0b7f75dc8064036f5cf29014853004dfe33f55eafca560e8636527399cb1090f0e12b42aea5babe01e960b6cc5e1aeccd5304b7128ef0171cd69aa1235ac5645df381f43d1939ca50514cac467d65f8c428d529b556415fb6f6718a54b1bdf818a93f1c5eaa0b7192fc2e88a4343208bfd7d7fb2dd1cf6379e9cd7aa15bde9fb44c18549e0034c379745317fb52185f93e63835a9d8b372e78195db2faab00dead1da0d07737c64fdaea8802340d3a6854dd8346ef7d75f58de62b8baf6afb36b01a8a7f70469cec92cc967b1444c051c8730500bc65fe55ff00a8e4a62c7a358f383d593c7331f764a589f2ab12c4a7f930fccdfe24f43ee85b38d984cd912464ac0ddd9a0c1daade12730f676013e1af2995e2aa3ff12cba4c3ebfc61d2c1229d497a791e8aab464245372c74a6017f7c96fc2b9190629885760fc94dd2c8b9fe77004ccf6428812877c549f44b5350d7e9c66ebb6415e77fda6cf626b25e27ac210197684213ab382aafe161f9f0c6814e82fb2345b7e5ecd973a6c562a1fd5760bfb4bd6d35dc43240e6d8ee2255dce11568979fe22dc34e404753a66c146f34dc188d4b22bf2a5762f858c385d0d4b4a7d482d3344e35aaba;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hb68f36449f28e02408eb35f48aad75379196eb1f6383597b362b2b8c42bf37881e1d1963cd89a51ea3f2038792406212a05e5fced0d8e9c914e0f678682b372d5d2b3da48a9e442084c16921ac35ee9cbe801fc9a37186a7f3a3e6d7d0e1372213dbfbdc31ecc9a5ce294f0081127c627825fc7465946dd020ea18336be680096574ec213e9553d2058185d57daff9cb68f5af098d6596891b98c2d612d2270a6bc57e1f031cd6530d350dce15a52985d5162ee128ecb80e1df43cbfa9dcd8bc27d628cad4d147e01bedb025234e218dd2c9be4a501cedb628282f08e05408f3fe5db5a8e5c65c7865faaee7991f7f05f9c4957f9e0702221d6a64219de7940c910a734a65fb1e1e0b901de58b74f8e3e5d5124d1cc00a9e24002023014bf710e66337fd343140b98fb100b08ccc32cbd06d4dbbc973b03d72c1a18c1a862bf077f63bbdc914a068d6c2e6cb447beefb684fdbbfd4fa586fabe29761965479dbe488bcc53588e71e13cd4067d0c4892c8bd46dde52cf089070431ed90cb380437f16e37d9a8fbe950f802cba7e1112ec6a8cc52c0e9e94084f4597bca992c2c4be53e5a5dde38e5429b4d4e9852e60921253b5eecd6dd03993f3b326a721c44b4469e53972d984b65f782f870bfa283893e3d9abd2006605536ae38d0060d9017604dfc7fb884979bd5e8b0a05cebc50f22f9cc86d32b789caf2f6378dbe736525d620920e8fca62dc223e24749e1c5d945773abe7db0e9a975fb74d8806b15ffd1598d5d45805db78698062bcac8ff2e622aac869353a4368038b48a4e29469784ca7386d7085518798fc577389b61a61ed2d9cb361e420a274840219ba9fdfddc1ac23d08954b9c1c9bd5aad14a88bc646362e01f3b2b227180cc035b74e53e185d6a3784ede440ed79b955b308a31c9be7d8146b2f5d8f9a3b72df8bff8ee63407db1a77657badf2498b98c2c664f42ed02fbf71a63dd0e9b925bf57835d5932db138027dbd5cb9f18af272e1411b23246ca0880f63dfc7f6c5305ab33b14052c528a79f60feef7943f4bd2e3dbf3b305b7b6b0384769b3ff304a08cddea8343dfa89f8cc51dd15eddc24f17715115427dd2edcee048f58333836c08f93b5a8e97558479b17b66c31ed2c2bed37604d4d56e441ec0fecc0b5d00817fb8805758583741415f90ffc1b2b15fd61f02467e20492ed5f92b2e5c38da76ea1b80696b4e0a1e0d387b1aca3eb5dfe779d17ceeee9db323fded669f877b50fdcbb9f4be5b99a78bc42038706b0852805820a7eba98b20c5110f1e0b9cd40136844cd87a1f0a36d8fe0f0a878d8f7bc82fae1c8bd3c1c2a9769a2c2079170535c59707cbc2e401103ac36a2eadd4c34a87980027836337d889dcdc8d7e4cd1dcc4ad33ed1f2398f080801e01675760a22ade9891c34236fdd5b907cd8ce31bfbf934d45b63ad55ca427bc1bf160d09bbc0347c04b5aa96ad4c54835c2f0434a1c6fddd3001154e9ea956c3cb5f947466b2330e6ae5ad1fe4bb20b51d33679c64a35bb9ba7483e3af5109745caa7524945ba1beda5905188183e2bc6b9ed484f68f49d4288cc031faa8f34d3e241582595d4edaf24f1c522066076e63f8222115c6542d7556e492e3df7ed693620752be2251acd0034ba9f6f69eed2f82acbc74c0a27de1573c1a6e4b19787b3d3ad7836e17d1c037744de549d22b82a47f5c087721c1264e963bcdba7cd94d95c6af6cf879166c9bae3fd8df8695f60590533ae4a00f0a522b236e2982e8155dfa0458fb29a3e7611c319927d5352f8702413477c0900a6c593637eb2512b56ac05b0de3d6ee51781488b248686a0655e491bd3802cc6dece6d58d92f8d9df351d0514736f48e9988d77b264dd4832078c657702b54d8ae51dd893a7e7e762d32751414a3c7b8a84cc842d47ede485584914cdbaa4f4be48e77d8807f77fdece372c8257a264db8efc856325bc2e6dfbd4702d480187ef44b6ed99ba44bfffedf429708717e98cf81bdbf9a71473198113b6d22cf87658ceaeba59ade2df127dc7a59d0fdd070218192b9961dae48b2d142bfe46387c0689528f5130fdcd178566e06243335dc424d7003bb5d9e13051325854a7683aae0509ac903481d00b7f243e5a23131af58cfbc3369a90da403d5823b3bbfa66a8bfcbb2d53b7c25e058efad4a6fbd6410686475bf37c9c45952381554abf54e1dba68155ab4aed44e29448e8fdf4b55b4d1fcbf3fe385c2f5bb19a1cdab7895d8996b273205c3303215a90ab69455346ad8131608ffb67a5105ccaeb98009eef551b5b0a1c76a64e8897cef655e4f49f7c5bc9c1f819c01b273b3e48a5a13826e3bbb528e7adeafd068bf5d8b6bf780ba5ae50987f288738990a8a7a534baa9ccaa61500cb47f57b99b17e1504947ee981ad4fe317ab73bd154687cc5c479311f47b5cb0458c6349faa2fada8d92474ad110063687d395641cedcc9e1636190a2293adb8b454beee826ffa833fed36652f2e25e02a8bbf12a8b0e70906762cbbbba256212f96da1ea01fb937252f8558c5df78e78e9af425c2e2abd6d0c01186d0b8fd93c64dac262bef5a6b81f80e63f72780a5ccc217f8f567104f196ba347d156c7c2d76f26c1790ea36115de86ac2a6dbdff5d4d5ff3f62e8a15ba0adbfe18dd92909dd51b9ed9d8232c0f8b61147b33dc38f7bbe8ee8ef12cacef8483e9621d12803cda1a25beb4f5eabef9da4d9f623d736a15e36b9cf1748e14910ffdffd360d99a1c77aeafd6c80b08fee03546ac5e8df102e8ad31faf011b8168a8c80694427e2d8e8f0a6305daafa4b3873b3b8b0a6ec26f48112f0857c3d69f811a3c82d120dea8f1721cb0c5ae24bc51b9b3d7d4abe5ef25a83a86a7302f92d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hcb6745e3d140639f622335a945958e7100658a740d9aef3f050d546391501f89f566ee393bc1a66f576ccfa1ff681262b375de8747666362e47fbe3ac9c606cd4a2136ec60a35dc2620426bd6fb68df886d02380d7b39b445f2e103a4e9880d0750ed4ccb5361eb63a6498842153996d018c182a84098ea3587c9f0c1cf3ab0e06719eb7c2842a161290f59449eceb13d0e52c01af3544ef07b8fd2f00b0283c98fd1da6259f75a3a06e2026e066fa9384d1de66bbc23c742eba63d328bdd64fc747d9baa55d6ec12696440736724f70d9e1f62d6b662c5b60cf593a669a3aecb95c797e87e7f5522040451187c029216c83dde7f6e2b5f2717b877d909a813069a7f2f169e4549f5deb51e070fcb57edbd6f3ec28864945241844cc4db8d5d7bfb48b646b6a48702e1a1eb8fb42b6f52dae3c64722e10c428391765df17b399330973c37f128d651fc57a0b020a6bc3ddf4c88034fbca0d1d81a4c3017bbfaafbdf23fc863de34882a0bd7f25131c0ea874f46845f98ba7adececcb700361a63b50aeef96cf02fc2eeffc74e53edbb4723186cbade4f5e19bbfe4b19805448c8ee467ae01f7680c0229be32286a7790282264751efcfe8b201e8256e4ae51aa2a1c8b5276aa54d492d8ec4ed4580cdb2d4196f9d4bd475eea098395ee9f7cffcdd9214579956af457def6100f7f0f206a9d85081ca732175df3e3e9f06cdd70d9d25c6bd946f25f9e01975d81721c50b60ffe09463cc1b4bfa3669c18d1430907efe178c6e9ad952412436233421119c2b0a21b3e6a42df8c82a062ed06f572d0c6086907ee70fe7954f27487e45539f84a06a4bfbb20a709d2aa780c26781a780cf4787d31249085f0a348d056ebe1f860b051684fd40b13e0819696e391c0f23ce2a7f3b35ca6b3b5e2ec8c1fa98d0d839f3b966547985f2ebc7cc13e710149d005aad0b577f6c689e9cf1adf8f3f9b58ff68112b5d32afd493caaa7d698dff1abfc409ddef49acf24d6833319150a50581af6a86a9b137217ee77ce10aa7332362c96dbcdcefa0f9dce3dd3405e873e3e10671b31c908ddf612005a432f92385174394d33bdcb5005908611c7b650e80c09f1d43873b13341f2a761e5a614b5c04a569c5b5e02007a5e02c5bb12481766937be861cd4b3a779a6bfd0eb1b00ad12bfe37b1945ab2bff4b03403dcf465e409ed6750560e97e30714a0bd041495934e623e15b8d029ef3b47779f821c741d36849d481f7038e5065ff75d825fcad80f644c82b9286c8b2ed6b4ad285151d31c0ce7fcc6feddb68624758669e750b00b1578d1fe3be693c45fe3ee284e5404c4a3117a69cedd869c33d679a6dc1e4a1da2007ba8c944b83c5441782adb6ac40c4520c678cb8fcd9c330d596de0338f25b87e8a0d4b063a891387d2a5d99d009a00165f4c574c15066a596e210ca53d91901cd90c0e42804bfd9d031fb1fdce2e1ab533af897f867994ca0fcc100ef8665eeb0d1173f992ac3028868b46253b181096f6646c5564752541f64c1eb8ecd4993e3d7d36f952f623282a7c8cf5b985fd61ebfc403b017eb8a2826cf6266a86cedfb24001576492de836d8c6b4200a8377e81a0b2e27d0e29da03f5ecbe5c911779acaac7dd9b1ad976758ff15324f2f6939caed15802200ca7f04412484ac54d91da4b0df8df1fd704106f6ba8d86d505bc6df198ca3757fe82f531012a5e291fccaae33240c4bf2e51f78fe8224224d2050671b590dd1b82f293673dcb0de76579772e46b9da80259f5ab86130bb897d8e7585ce5ab1f442543df07f695f0e42a8ed4832923b097ab4b28d77fca08d101219818ad9eb81b07fcdd8fb6b5afc5084804a8a21cdb7c25f6e62b36129b7fd4aa26cf780dee89c41415e2d1703b449dbed17198266c4ec9adcd6a66e24d1ffc78f31058acaf0c16bb451c1cda6c7b4f192a5ba016c238ef492b9346c7c4155f1bbb72df16bc3972e0e196c7e1481bbf371b0a671cdfd8955c4f20093ab39fc993bc576833d5e97bff11e2d971cc28b29ace1b75c207d390839bd86b2261a8569d4ba7d3392edce7dfb519cc14585c305a1b1d7a9622a4ac327ab82e3a76ca631bc71349364eec43c66e670cabce6f7092c53865b683bb394018ed1feb0c7a8da0a815944dbae764a706e44826eed566bfdc9094034a487444fbf45065b5f020eb960802f2d14cb5128d6e3ad9e4ffa45d9f3872947d2e5cff95e516055e05a407da4cdddcb100a0989ece0e3ef8455e21408851e9ea7c911f399ec7683e948e869e9ccc29d54a087449a661a10ae564acc898f4e695f7dd79647d0ba461d52ea53459f2d50f9d80dd7d4c189c66f9147cf2466c172bba7f88a2a1a8a415d33e3a784f1b787f2e2fb122f78ce4bc9d06c8a14fea0db4bbedb0beabce2bb1c33acffce53f78184f3cbd7222ec5b578b15363b48cd6b78174b5197405e17dc6752313dd03bb9c7fd461037930864030d04ec37b7177683062e8446ba1948c7c2ca8261d3373393e501964e89049facbe7f4c083c8fc4c4015f1426f9bddf65ab7ed2596c4d60e339974f8a5afb262b44f789c72dfef9a0f1638f23f7bc96147e65f90c66939962ee00bd615c64e169d80472577b03a5ad47d1f709cddf319ae4cd25e03d1fc92c8ad51ee6c623ab9965a4a5329563d7d3d75eb94013ea0f521543a5d0ae5cfc31dc63017c82c113603b88fc9384fbd91bf91fbf7c4d3689fd6c4e7c7dc84724e96c3e33dbf0ce3f2037c4378474a74da850acba35728364a57a7b339587686fdd972f9551cb52079396d1dd2bc13712778f24515faa9d659ea79e328fa576b90300b27193d8f0d0676a0d275b0e04b91676b02df0edcb57cd0ac54b5de9d87fee01462e962;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc8d9471673d55e49fe53cd33336b2d007b8d83fbeee113b9745893bcada514d51dd58cd8d8ff913bac65fe4ee943eddd1658335d6ed9304b84306eedd3fa2eb80a7fd8e42b16d6dc0fa0a7779c556fe15500c149699f16104f7cc56fcbb6965454e0bd40d1765fee8058ced924f8700ea2a4e2744d284035bce7c5f490789d7dbaf51be4b26d4fac743bd32f54b65abba105422b5afaf0fd82a85fb4aaa4fb827e8d7a3e360702d9bbf9af6fa892d5e459347bfb1fbe99c277c13f96dee63bfd3e86f9322dbc965b2752643a2d2040a2dca09ff8d9d1bf6dad01993c3dc618909d8c5f38845c8ce80442590ed0d5fafea810d027ec5b77001519073a890d0b05d37af5e07be55c6967a8d71814ccd97f06b8337b4f292c4cd99b99fd068277af687cb0be6f6e57b783d00b116f6629a43542d9abe775e0ea534471d99e59429a0a026570fbe2918458c946ffaff2fe71d5f8a41f883180469532fc6bd05e82d680bda57a890d4edb6af9261be8d2a0cc86faa56b0e1c95d25079c5e2c2c4561eab2c417ef8680b7f67952bd3dc334b47873ba0c9cfc28a8a1de12e461d94aa082ebee341fd5d25fdec67620998dbb9a25c6ae3d7e9a1efcd9d24ec4708611020455ada61b4df34747de8a49e8ffda0904784911afe3da82ffd042a26d27d010c6135525b3eaf54d64a668767fe2f75c05a2c24aa903767abf875eed3093d547d31b5b020d2f7f1005373315926ae0384622cc7d19f32cdbd1854ba92decf993e7a13af619c69771dee02aee2d4de3e255f2d626c1b38c86b305bd2d6fc10e0f4fff049e0dd17593421f08653177d1d823eec7cd4f5fab5eb9ba2f3ca7b5e00a0daa072e9353d500e097d20e4f4060543a07651dae79c46d6e3b6a78d8000ee38e3c991dd4d4735f7cd72aef17c746319db5d7ee40138dc7eda612e6cf57cf9591ebfdb1aac893beb4a582c4adddc496aa9e7069a74ddcda339ef0e0e8abec209e177de23c54393ab6174e5df1600371148954b6d268bf95bcff0b071ee486bb6655ad1aa15d88932a2348f613551b031bef9b7da85f6c325b61bf191607827084aae1f953355c363f87739d0c12164cb07faf0727e9264f20e613ed123b2fa2eea4f5075321340cd62af191e4aa17712fcf62e5138912930c2986c8047948191d0f1457aa571a8103d722e3fb7d2cfe7ac11009dabb18d69803693d81dc16fad53500d29fe8555a6757f9535b570fbbe54f48bfa436e18bafce1f6ed79e83dd2bbab0030508d44107a2ffc5b5060105071a7bf9cd650d2990c768eb1167815b364e67c9ec2f238826c60749547a6230f17245561dedd47391cb56ea876f9d60f6289a8e0f8aa2295376cc0824684e1997748c9bed31955df8a98dc9c0f051ae6f3ad2f9aca2cb837c65304b94c399785fc139b6966e0d2bf6f68507455e1365fba2323538ff28daa1e513c5c105c206f90080cec09dec67abec839e6e91adb350e28efa90de598f51feb213566c7292accd265259499ed4a66350ea3317ef8ba7785447f695c9a1caf7fc4973288344f0bfe8cbef7e9e2494521fa0795584ac648047edda336605cfbf4b85cf2438999da1aea5e49df3406d2fb0f58d17f1b0a383933959265f2f3c3993c5565787cf631187e961ac588c27b55798628c3cb86a2aebce31c42457c1a6d6d1cf03293b3ceec659143cbac574027f4fd8cbccdb354c6dc14e2ed0b8505a20c534528e2517a9319593971b9c017beb25f5c60ac5d85e7fa221d880753410f5e770bd306db657cfafde88cc476323605fd5aecc99785df66bbfb18930fc085e73d76a97831c646aa0a4e6958af7af563b2723e3708cca224545e4e7669ce14ce9f4fc2f789d288dfa902ffe6f7e72e72a5dc560bd8dfdf982463880eb04bd3298d3fe31845ff69a9658a2ec6881c34647b3f95b371fce82c38aaeba45eff5b5cf4cbda41238684c431b392be6aed74215fd0ea0f7d1eca4a519d1e5ccd3caf4d7c6dfb5660c576a633a856dac8282cd8221653c92cb336b221b649de62751f3ec45668a2818d49a6e0a583c0085cdcc07bb80b4ce82ed192f9a5134027a0a72897eacfbf84b37b5a55f84a04bbac48229fcf40c66c06e41e6287ae168b41e95a5299157af74fe8b4462f782a83f59fa9f1ed346c1141108bb7d3bfcf0c08325b7a0aabb146fc3e0583ece26089586dfb4a33f6df4d844c25ded746b8a1948194c747a97255dd1bc1a40271ae3317e6a9dbebc22c2bc41680349a9775d525f1632bcb8641eab64b5bbb0b13affbd43d3cbbf637a76801e307925ea389d49c8497948d9aa02a321a2e2d2bdc57a8849a48f8014a7eb9ce32b06e17adc50e2fc12729385a72dab11557b2a72039f4b6e96bb1a62e40999f435302987cfb09631b9a35d97dcc0fac31bf2182787068ff03f142154e6d6100abdb1146014d0439b092eb55abe8d48cd718c25eeba3b3f5c4d9138cf95a31225e244b8bae93071cf4f52bcbc4771e2ffc1592fe8cd913efd54aabe9833ef83afeb4e41a003422b7a20d5f3d5b1008a56b0e874a9dbd06a9b87c9fcd585cb83c0e32bfa483f2a92e0bf3cfc3ed5415f5bfd79449939bb3f5d0941ec85ccb2e1c19bb439e40f771dc4b3b065393cc7087cb5c245a3b6cd131ee02e5665007887275525ee06e76efa921a9dee78e5224486f6e9f2171ff620ddf6829785001654b019ff8e25bc82ae15d99804daf45690910acbc76934f3fdaf2867c2d6b2d1d916b1e1a952c85f5010f768ef48b156481cbc84a631b5b63ab6fd6c83b4cb554ee019d99085e7b65d161086f66707b3dde49296ed51a61e1e2cc15fe0d6bab617310edc0ceea2d33580aa8eaa9c4a5e211d4c165a9ac83d15286dfd0c49a5af2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he0228e2c739a2705d604b9535aad3eb7cbca922682c3952e1efb0b4e6a6c83279efc137aed0fe9fab16ca47e93dfb1f8fe4944c0157c437ce0ea2fc7457a1f10a7ebb3c653c364aef48cc9fe9199c4b1405a67445cfbac246cacaef867f86c402fad2d1ffeea4e35ce1dae1cfda7203d9ec7fb4374b8cf5639a701ee1f4cb38f7eefa1a7aa91c8dd90f490cb2c147c032e3a479d0a1205190974d63f8520098cd123d7d776c5c94ffd63cbc1b75e82b527721821373cc90c7923f0f6227c7c72e7107f3cd370d300d9ca35c6f8b80ab8a4798c6c3f5d1d0c16bfdfe71f64dc7e6498538fded85debf0af34f472fde86b69c945fbe3d992d2046b1d1bfc7075860f33700a557a74c928f5dcdf1fe16d2dbda2f3b41a80b52549a969f9e4373cbbce91a5302ddc054706f74871446fc5f31386d7f1483126fcc746463cc01545aa272605ab41d31149a807cdb4f783d413a6275edbe568e193814bc9c7af195a20109951c9641cc863d3f5db64f752f73560ff78ded3eb2e3251842eaa92e98473589b3dec1322e2ac3890e52cca662cb8118c48d9a6fcee4ee6c3072313fcb617259f9385d185c81671024fa1f0bd2d7ebfaae2408ef225cc949c8172237fd2c5330be399e0913676040a2539cd0e49c656000e91b31932c2a4ed524b26d7716505d2643841ee9d43d3b99a96d4956a9f3864419fb206f63ff2c2ef4d5cf978ca4923f312d89356b6e24295978ac91d8f236a435ef974543df0261c3a0577a3ce53944a04eb7083a115a30973967c072eef4a80fd5b8f26e5c1e1e91e2d891b35e7e66605ac6e14ad29a270be7b102bccd6b264850e6450f1e2078e83a3fbddb0de9f4843ddaaa24c506166cce0001dd0e4ae7fea6696ca0a62aa31b7b01f7fbd901e2e1c683ff9c58edc42669d64dab94c938c9bb4377f2e31763279d7839cc50bd340af5cec070cefd0b33724375888813778f5f1bb6d5290f5ccadf7bbda4fc902cb61c1924fe70493b23e5cd84c867b28b30698b87df147725a9047b8e26c8e2cf29f284e602679fa05e4606d51c7adedc627acf262852b4877ac46169c6e4b991eea32e5d74ae32f8d57bf92bae66c2af853f774b1d81c28294f37aab21b6568b24c6b9846e581026af0c74a2f84a82e568e4153931f2942de1dc27d284eaf291231fb1f52ec3c78a3959192a31a0a008dc76a44495163451ab5ec5cea49c6fe1aa1f2318a796ca846dbf147d38dc18610e1be19eff73b9e0460cd1dd79e51e7dd25cca97efabb6b7c261ac878629383fa3b44e844f0f732563d0605286fe0bb8c738057cc31bcd427a43f902b5fcddf98302755dadd03f986145aba2717594c9a4a72826dab7a96d642cc8d004f7a634abe1f5808ad140f50fac0e1306b55105612870cd6ec67c262397da2087642f721bc2afbc47b50164491aa079b9a17b76cb7d8f7f1e5cb067e674bade8d24c34540b98b9438fda79939c0579debd6de3a782ccc5c9ff531a5a2bd5419db21e16e6ef477cd96bcf2e9e146343847fa2d4fc0116af4840c5f938b95cbe6d3f2b5da38f5ba04b96c38b9faee208f319863507a8d3993293dc693e289819f169373537ba6caaac35502c4cd6bd9beac1c55d9fd01071f59b548ac5c72b8340f1bc9268d77ef13e5cf49f6a59b294de445907341629ad2d9a0fedb3dfb01daf3cc1a536cd11c24d97c850d3c4fc46ab4fbb4d13a343cbec6fffcf1e1a353649e75bd9ceb8581749432c7340cd9c2bea2131683c9b390c067d547ca2572f205b9325de980f0f77790fa94c24b41fd9259949a1cc916a4fffc9f80b8bdfa40c550f33d5dbe3a453fd87218cec471f011c9e330794e6098d6c96f4b3f2f39baef261f38d498275a594b2c1f9fd77bf7af674e753eba0318eb3190f2f508ebd020dbc3a6e78bc61bbea5a0d8763f0b00dc144c5fd7830efd9f35b74e376688c54a6a948fb1c2a6a211d0c3355d64dd6bb57a353431846c8124abf90505730f0d74506e16b05f1f811491d87ae4b33c50be97d5ee9264d671c5a4580565140828169101136de4fc262852c4056d2ef14130325a89f77b727e48a09d97ebf04b0f9c9f786afe28323a6694d71ac695861fc91b0444a4e02e06330c9b63eb4dba6cd4c4a37b8efcfefbcc099778d7392d6ece8e567690afc582acc0887bb8998dce910c00c4c422e8bbded87908cad744b4061a14b73c7a279676a9c594e871978acd05fb2d73058d04cd19955f88904c3c9987610f95933c68dbbdf8ff4dea2988a31eb6f415717f9b9c5eca7b0dd65045617e4dffc2b2e84a5b160badac3363610e1bd5c08abcade3cc2a7d70ab5f5aafd243a51a9b340138622330c0e41530b1ad8c8bc729c5155332cd0fc77603411de8a1dae07381957000e5448852d078ed14aee49aa73e429780a990b92bdb5ae2070b765ef57226d6e1aee495ccad42f027966fd642075c20f2489bbb143315134ac1415277862467415f675f3e71ca5b91a006410d9eb354b560c0364cf65e2bd942b405061162177746d30c9e904ac8cdaf2727c05e82db8c3869c5948a0314d5e3d1d8cca7a14d4e0a4df34ce25ee38395603e8cd55d220800ad077fe9d48b5516f2701642b41fc240730aa0b86a82945d54ce9bf3e4516a6dd11ab5bb240be3ea4b7dc6d21329f04ea444660a374d24c00cbd761fd43a8e4b41ed39d27db6c05cd847621d0c30dbf7000a90f0cbb1054cdb15e7626d12c5a497a9c4ff5cc56dd384c403f094b652461cdc8b47b3f1d950a08842cd1a0343599c2a383c68d9a3dd59271b4bc39eeb36678900ff769a9a9bb93a552dd657095a5d24e8cd82e883f76e8a91a323ada892095696e1777ffdd0726c7e729cf69aa73b822b0e0900201e0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h1a28ca182b6786654613329ba7e9dfd04cdbe561deeca7966652719f2b0dae016a8352bd2ed8a9066a2086dbdf69b17d5eb22d956fc6b08f6688719aa8f311d26f46de0ca3a1858da45aff44d89328e2856bfee52d7c5a1d1b013c8d5debbdc8b8b1fcf5353022cc411c335ea67a2ed7bfb2799d51001d383cc49c83e326129c9822fdc440601fcdd11e4b9b511293dce1b80dada27f107a9080df56e0504118d3da976c3b6bdf1d5d837914309025a2a8febf3b34f72e28f30291a7efd43f4f3902721cddb75ea24e76e618d961eb8bbc02b36a900c0fbe40e7ce26da114c5056193c35357d257695d533ab4fc9173b5b566bd2113433a04df09b3714625addbcd692dd91bc4d2982aaf662c58b184c133cd63a487974aeab405a488725edd528a31580cd992b1a32777505f9c2073b2279f65090ed6cd37505d83a67299d11c9a818efd1617fdf11419a6fa101976b5951f492961aa081d184a42512f952c2670885129bfdfcd375a95910abca1e214ffc3c340ce1868d6f78c6cc7285a7f23e9fcb8f9690056ff9bac6447edf246b43741823193fda0e3681fccdde29a9c29a6295d5a0a4cbc10d59e783f55cc42286f799bfa25ba312541133d92b290bc150c3653938a3581e297a4cff101438764416b352dfa6ee05251db6894935156d4c88e636fa82cb22a1b8b8f67404bec2c0e1fe2f2877d26bac60c1c63dca941f1c499c174e2383186dcc9ea60fd0cf6e805b6c59e0c36aa6463a71709e604f57bc5e583d60ad8f76f2a38dff9db2d0ddb2212fbe7db47f5e0104983018cc432c9b06785b99a3bda3ae09724468d01c064b272eb6a91f68abb70e0e3e863a5cfa15aeefb77db6b153e44ba700c75128c8e8a65cf82b4d58541a21e64cbd25eab913e4fbe9d38591cc934b5cc8ab622d5ca2ac5bc3b91628496bdb7128ebeac52a4eb36078a57978e07098755b5837946038554cca8d7b372f14ed60fc3aaf85f9823347d36eee8676df9b66fba578f70416f4347aefe0285bf2feab52450725c738518c63b839c722e5ecc7c163e00e041dd5667ba4378c7c0f9d4794c60395de10310d8ff1ebe6021d2d182bc63bb61b56644f9f5a60334cb5ef52ef99faa20af3b5231f13f20787483ca809a9c239506666ee00211d710ecf1ddeb744895759a98f370da0ed035f4bb9974df1447b249aabc2014b9fbdb7dd838a74b1653e62c379dc910b82dfec582ea96b70f7f7ea7211f7b388a2c7e8ed279ee5681669e857589201f54976d93cbc3bc3efcc4542792e7b7aeb709aaee2708856ff9522264e476af7ac442ad24d15eccc18e3af9dd782ca7133cf264fc838be358bdf06bba6e2419bb44ed621363776bc532d30e14465a3cf33377eb280a17f6e772e207e2a907c710388ab2463439f52f3e907b302d02ff4de7bf6fe1b6af524f3bdc8536f8ddaca4f05616d0728b21c11a96a9522666fee27d5f19e154d25d9b08e110bb0f74e5c34c663dab1edf18a6d396355f5f892d7106fac9dfcac15be10e31d56085c92a38ae5bcfe7c463bbca0c825a09bc35f2b87aff5a3b121a5b7f0cf11b8d423cd0c6efe92f6eb5d149b96211a29f50fa8b89ff0a4cff0e21d2aa1f401db6496c74acec53ba65d22ad13543dade606f9d3681f89c5fa74279e6fb89961dea9acd84a60c74f4fdb91579ea38943ecb89afa52425c44855dfde32746ed5371a76b659502cc6666c5e6dd3e3c5b46acf33fbc340c11cf74022d0e99accca3722f3b84c8eca27bc943eff48c2e0fb1318b312e11be727bed8b4c18c18ed305277483823e094b350befd431c3a597b62b3980b683e0dfd5699e9a82af930a7ab9b81bec78defaf0b05423d2a00a56fca3c2683b1497e991201a4939dde3022733d3e8e8d917f5c62914960d1f6570b99fda3986946a3eed80df66d942c00e062a7f7b18131e95968fd22169cdac3862eb8efb3b4baccf818cfe9c63769cade9342edbcd5d42eb8b4e72c7fb1110e564c91ed2c3b86ecb2962f7c67c67cd54d7e064848b01c5452775510dd2b8daedb72d5e8134146676dce19ac2161fb772434ee2a016945be776485622a6b5083784945acbe47d2c9367863e2f9e552c4f38bf55ef86cba04569ef665e9e73f865938dc05829196efbb218ccef33897707906ff820553727dac107760b4461fb2b17bca6e74b0315243a09b350002c6b33bc87f340d69d8f5bc8a486fa7818f34a1ce9cabc9755060407e74571f8026127928f0081536f0d20c674199066309f85acd9d4f203e2b376ab43a98e987332204c7dedafa9808043c8c4dc47eb67fac34af86063900434258211c01ae942fb9d5bb264dac453c6e90ad2b111f52946151ceee9ba6af0708dc1fbbd4153cbf3bc7b14fc84c569d478b72df5bd92715e3af9d42905876faa3f4de0889cedd142e739cd5556a5b89fc10b75ed4b2189b14a2f8fbe50ac075be0b52eda08029355237e4dbe156a9a9f83e1b609072bbace86a4fc92d2f4de855e7be48891b6801c088b53bb2254845976a448931d124e2b11de9e26a9933d7b3f0b506c72b3d939af66f15edb4ef3b08e8e3ad3f5dd24c338fda0c221b6287a3fe1283f144b760a651ca011f0011e79ca1043f0692fddd0d94010be0591bca2f6250e4345d12f5ec300bd1f0d70ac9af6afee48b5251d6ce16c8171e27661d6cda243d9989927277e6b757e15163d3f9444d3f819fd60976ab90ebd0b23f775c9646ceb4769d64db0913f3226830f26a280b6b0639dabcff2d28daf7b5012f4568b6cd6aedd98bedf4cfd8ba2b19b85cf87ffa9ddc66b619c03ab0ae4a7d1c724003ea7b09cb6e1665d700ea7389c150ac16376b45adb7412d46bed52f7e55f865bdb87bc60259fdf7f60;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hdfdfbc65c2ffd2a9104368a598b9f6384e4f44083fabb2b28a70c5c3cd53eef9a0bfae68bfb949d5ea9d20d9ef84c08020ca8ceb74a2fde1d890d4c6a6d311846c03c948324dc4beca732157eb808f12f00108978ec26f0d3e2ca81dd5aa5c40bbdd7aed740d30e9d3dd5bb166a86bf49c351cc963f40597a70eb112faa50280d3514f7fe32d7241bc6825f99e5ff0bfcad892a747c629795cf898d57fb702fdccd9c2a96d16c159778bd6815338bc8fefba69bb630c37a1bd1c701e1597d20637b27fa9674ba4ca8bda509dfc8bbc3eac8b830596b6a86b3e323ec3a731b8b8a1433a397cbb144b02c4db525064e6e06967c5a81ee1a8b7b3694ff5176c48da2ed9826f33a105a9b735c6fcdff34ea8736180a06989a0941cc820c5dba2493c2b96724781b1d56568c0a248576879d6f125417db9be26a8b2e304932f026d755a17c9c39f464fc5d256711a8155db36f873898990523b0ad8b162dbe758b020378f66c1f92560cee5fe56b76571e5b3cdc3aa51e5e1c806b1d688921089697a8b93f2f26b5c32b82a54f0003054b37d255a76eb95a3fee7e70f3e12c0d0e1d7183a9d73b616384b47fdec4c0ee120d7fbcca45cea1c59325a34216d57d1a758d3970d8d41f335d1ab936dffe04be966ccf72224c9bf528b277c164a3864e245cd38cc432c2b2885b4e27db0b09c2abe0be06229fbae5b2815f0b48673dc2c6d7bffec836c733081bdab4c340e47df7e5d9194d94a4e6ce1065d3ef110e8bc7c986ba0b843f484cdc587b945f3d7f61606625ea6adc6aa039e34c6d36a7f7d7cff6003f21abd2ccf9535808fc189b7fe8418fb0757ffe6300d0fd94b4a230abc4716f0f3ee48240daa2b14512a87f8935ee7e2b6e4d901082b091ae66abdd2ebc9afd92f1bead1aed6efb24f32314b96ba46461d306851e292706f10b45c9feb1ca15fc3859baf85a0fe1c08c5aecbd7da841965b6feecebcb4f3116a40c75641f340d7395bba2c293c107ce1de4c2a8b195d5600a873c0b176915c3f0a7e3a50d459d7fac19ff38feb998c1417e036b0ec59635373aa284e867024ee4c8981a35c4a49ced8fb29e05d2443b1a036762844c9e84346438573bfb2bdb1d117c5cfc0f72c3cfd4a6e33cf2462d4f2c7a82d48366a086b0fc8f5f5744cafd8e8f03122f85e0bee756b1ad2c6e820bcc7dc098c0825cd150a7a603192fdaae95cb3932630d9d2e4d2f55636f0ad14eba14c1220873c588515a34a6ec45ee93944f1f7ac5e9a6c596da2535b30dfea2f22500caace5b1d3aa809b16357300b4dd84f5f5f7a2dc511942bb4f03db9b876209f83c23a2a3f2ec194f869a15cf999d1bbb7be0ff100118f526bc1fe68c12e34356a88403b3cffb59be62929457557de32b61f3c3454e5df6afb126c9a8e1bab4c22f4e039e5dbdde75c654286cbb0e6d2543b13a1e9e53735e67a4ec509de52caacb063f0474051c2fd6dbaaf2f4bf405d1d75e5053eb423b99d06776e21f3b55da10b44ad7cd394391e9b20318e79ba4274abfbc68efb5bcfafd7815cc03456636e42ed39aa166366c5e7dcfaabf83a54a7bec6ebdd7467a67b3b8dbc9ede20f80457d4d13ba7cca9f3b50b4be32caec4c6d4b3858fa921234d45e828ed4984e1f88773003f7ef7c8850f47b111be8090b143ed0b8a4c990eb2adc727c2ff8fe2c254ab16e89d7ea409d806a5e00ac3a2477b2f67eac736d4a23a358afc0aabf4bba2815315bb51a93516071aa6709cf0c7c2a864b5d855026c5df50b29406ef195eaf18ee65aa527555494c79f213723bb174b62c4ee7f193505acfd20bca7c82cc369eb2bcff218d42946d074c6e89dc40cb476238af5a6bf2ea8c925cbdcccf8f08e2f1eb5e8b0c30ce9630fe64bafe4b0fab21a5ba92dc9975760a50a7eb51141414bd2e5b0c0ec950f547a07f9a7e66f6a67daf0a2b8232f7d673f58983ed7141d22371ab87d31498fa378e714259c5cdf462d3054771b135b499995bec4c18a4d901b8fac25f89ed3d13c0c5d666b98fe01a532fac12521e0b859f7bbb5be533d7714faa330c540dfd0d713c9bbdeb78e72ee569d6bd36d3ec14718299311f92c09a844d24e10bdc6ac4f4e30f0a3cba4cb3df99b0d6234110507c850012712958675d8aadd6316c542be0f6834cc0393f3fdff30cf96c6cd7fd1411a572f5809b553dcf65913a76859b0538ac77be5f401ef6f987a6f3b531642e90427d21e6c616bcb068e77f406ec7c21b6ea3a5bcd1bc904a7b91b8877dc2716823b95ad0add7c696ad3d64684c25ffa8716c9041d960e50cf662a5f30171cbf01321e73085e0fd820802557391796515c2de232b6886c975448382554e127919b6c50910c3ca63b2e6f74cf8fb2d8c31b0d223820d418a8ffb23cb05b4507c01af07d172b7ab21336dff7cd6c8af691a1dfc9611ea27e7f0ae7283bac1689cfba918df518b5891d38c87cf58fe2bb6d822c92e7fc25f00c82e77f055c726801fc88ff0608fa249fe792f8a9ce0bd10e1199c3853a5a1b3cdb949b3ca3d87d25d370b5664069e5b2aa669605bcd7fbb634231bc52768b44d871343b476210592ed48c11180a4a588e6d62c48a327ea3848c7b754a0da0848a7418035c54eb40723881a2131278c3dc478649e3b7a2e6fb9d996adc393d6d50f0924ac5237adfdb50dcb7d7db4c6449560288ed1d4899cd597519e78366fb62b871e1fae9639a6e045a49bbb6c646c23f5533d764df13dd01d2692cf86d4f09796e914d9e602288af4462acd48166df06c8db44333ffb569f0d061d996347b9287ea48cb5491206e7d86a3f68e2b80f816cc4f2d45802af7db8ad377258a7852c0fdf7b53e44bf011ed78253b7f82f3c56be8d81d50e5e4649;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h8c11ec6228c3f1f2e5e6e75f44863c899b7f6d0971cdc3b5a669159df6e057f57938875cb6e045af85716de6377b615e6f87821fcbb4b00711dcd56bee55953430a6fd798aad84ade12b2053d44fa89cd0e3973793a190ba5866239c2eaeef0c850ddf3778e649311502914e436deda41b68f07513008f7dfab85e68cccaeaaa4a6ca3deb595c765ecf8bbdafa382a2e80f2fb454a6a27d758c39528447b5db8d09ba0192252062eeebfb8deecb9aff313a39155f9d74840e45163f1eac326d6a177ab7c0dda7bc310c5da3ac867b3db8aecb5bcd9e81be9b4444f163354cecc39f7f08f7907dd92dde17dda9da3b3f1663f5f7c4e6893f0088218a51631c73b6b3b41c8f2a4b91a39e2c375d1c537f240104084bf3bfa3869000c971401a16e48fbd10ba0422c3dc54fbcf3732e0b3499c908131a22d978beedc1177dc46ac19979c8b7dec7c88e52044c10dedb721e7098b91b03d36ec320a84ee82114780b60c2e64412c077995ee2b0f1f588fe1df5925b82ff16a53edd170e19a6b3f058b18cdb51b82636de946d748f63672d6ffec2cec6a81c6f922917f7c08f2558e25e0d59548032924bfba00e448c2550bb9ee4e93ea32af0863e2073d3ab826a03c9a873e284e2ab08d88af341bb88b6fadf30442c10672d0fa36ec1c827c864f7dbc6f6f86ea6de816ff87b3081672a877f0dccb5dc826c125f34f9e8bd6c2ed7a793424628d49104e0641d74295382514d1fcc30d61da6afc11c30ea84200600756cff7b7c21b997895ac3cf5ff1a9533cfcd6eab417e2aeaca3e2d52505c9f86f4d54c4b1f145792e0180d078eb3658ef31a269dd0bcd2b94b96ccad0310fab960733885e1abd005774c5164a865a158f75ad5e2d07b7e24ffd8d6e7bfb52c2dab8b0a675d67f605c0cd185d3fe58a0036d59b3c9567ffa304eb68931e0046e0ccb2e6090261394d97e16299a552dab9e97f616fd9b15e82223157179ec844cfbd13bc3c6bfafa346fe44b4f7df750273b8a53f564fb7547b21170ddc66ece2a79497d81a9a95bbbcfff12140b4e5057be190ff97f831389aea1a0120b2182e8ff87c8b2f398e8a59b597d7bab67cd77f97b30158b991d0e3c490209ffaeff3edde77c665105925e09b03c38c364df91e6e1dc45f23d0a62ecffe0cc1bf881c3893c544d0e02c2fb3718515c0310c2e72fc2196a73d495c142d72afc6e95d86570f0094f218531e98d87bb2f27d5873f8dc34a91421f169484f06b33daddbf4c16d9714eaeb70f33deb824b6eac62744e3218185730da1731492f2587ed782997c29ac53086dcea29013c3688a1f1b0ade520409bc6748d5a87aa26e656a82f07d6841338872e5c307ac09e5d02c26d793f8484e2f611d388d96f37fbe379d8cd5970b383ab99f1cb5ff5c93068345de5f123d719ef79a4cb245ce7c19fde9334397b029f5e250e9d5237bc330398aa8fcdf78bcf02a5b189f36ea5c5a79d38e1247e830fe5cda165c228b8bd31833e7e53457d30c9b2587df2c1ae6ec7d0e8f368bf76e1cbf9d044e09cc1f6fa3f8d9c207fd6b83e81ef55b87f4fca061b7cf7acf775ca53909c2dd94edabe7b40e3a7348e602154230b7c3b816fab9d5bcf2130d878d5fb49195e6435cd5baa4807bae9bcfa2707ec13941659198a2a7b5cf0420a07cfe9b8efc8b02197d4535a6d7f9a950dd2867f96345ffd77bd7b7e01f18f72401e9642cb3e2ca857470a83892b143827abe57fde290c031cdfb8c1b4d2a547a648c14ef9f3f0d2dc45ae14cddac1695c4a476338dd902e59f6faced96f82c5ffaf690e0fd089eb873ee234c5054159b74b152e6d1386cdd34264934b7f23dc4d88c141ca8dd16d260d114a5463e2aab81608d4ec587ac64f450c8308533963bc1e6f37a3e2b0cc5fe04eafb86846d95c088d590b93664c28a98a2802df36a04cf044fa0f3436d3391eed7db4ac0d9f033589ea3ca0d694d5426a1301c4b1760ec1789527232766bfddd1abeb132d74142a9c273edfe79d4c4a5dbcace485707eaf205b2ca047aa39237c650fed35aea1e59a8c6aa874ff6707fff29a5451b5e9da081f50c03285f1a341377bbf00cbff9aa70400ec22898ff6f79284b99f0527770ed6cc487ae0ae84c9a999ae0cb675a565c9f7254c87a42fa851f7fed3e08e611cfc28cbb60f5ee9106a47e262362a194fdfea2f9a32881b0c82bffb1d59df646005dff48e9c4d56e28eeb46a206e00a85c11c540cffc9cfee77718c2d7be2df81b1fb79877576c5ed135689cf03f10e27ced36f23c219c8abdf4ec9ad03b571e0db6df7a16a915c68f3978888ee800bb2489f6a95f7034db409ac3fa76488198237da93849662bde7b3ecb4bebdbbb6a63f0f6bd922b7f19e0a4800f62571bc4c49965dd664dbfc82437e3d9699fbd872f17a53c55b3f217fe00e2f2423feb8bf8cea331cf6ac716df372421098268103729aa6943a166efc4e0139b7b5846f271c89c4d4b9bce4e8344974f261722f74bcea289c942044ab18b5b7095efc2c4b637bcdd0752502e1a32727cf7211126158afcd4fd1912de70666ed4882b2daadd391f2ab9b049803ea0436746745e29bda2ec96f7f882c4c06b5ef725a549df94303041f86a08be9efed137ba4adc6e56018fddca907ac9a8b2204a9391dcdf23c0464ffbafc53d15c6afc3b432e3ec2a31d0568119bd667a7caae1127f62272224aee9c529d3104f844e630f8aabd5163da00f5faa8773d483aab9995fdaccf1b58ae7d1b68ee229cc31192b36d5c0619dc7fb94565ba7310b175c6026b1b0e53f941fc1d7a5ea76e4fd93919f7f62d7ccb102438abb81fe677335ac0bc9a4c7543bfa15ec236d95d702a29ba627bb247755ad33510dc0700c0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hf551df30e7adadadfbe56a3d5357fa3b80db9bda08da2cb198874aa36e336e017866dd9df8d9265ade83086f99e7464fabb7a77df298d8523756d48f88da3f544fc334c93e5850834be03ac345022624a74b010cd628dd8cc122ff9106d7017077d6a8ab4027fc47b308566a96c3ae66fc6957a752b4cdda62cf3830aa4b36fa6baa0afd8e31c38c04c1a0cdd90d6511a94001c847c62af52eefbb80c680cee3316bf9386e712610ad414077ba0bcbe2f7b7431a8b0cfc3ac86472cca2959c56018f473646ca20faf86e845d436849443092d4d4e9b5b82afe2d2e8fb4c7d32ca171d44305570737fc63e0baf076f651cc71bcb2b0cf7fef990ead3748fa8c52f2ced604f27b654081b21d2c4a4c608f332549ff84b1b94d684fd18951c2a0422f4d8f187a7afc0abd1255f4e1cf7e754f3a46bea6489c4c403c76633e3f5a935f90103f1c7d639aa0be80318fedf62eeac2e1364ceccba122bcfd3cb89325525f6c3b059b738642f8923342a8faedc474b309ad405a99a6fac1d297cf576b409091b31d32062a95721c724521710c30ec12f9be1d5c82e7d75145cb9e875668b8648c176e5abe6923bb919a4cffec7526c5ddd4ede700c727cc69f1cc9a47079647f36f442b8beaf5311c746705b726da3bdc5e863816ab16b6c7f8764f4cbdf3bbeee2f19644defbd5299a8f2bd44c60331f09be604839847ca41377e8fcc97bdd4eb5cf398b572637c092f5fb6a8579b7bc90b9adf72534004311d47ae79319a491acb43ba91398de2afa694a2faf74e0ce57d1ff592d9e8e1a776b491a306bdc6abcf06f1df79b25628ad83f210d258d18b052e6994f96663229998a59f821e6805b15b68eab88a8cb5e64a6f3ba6644aec5b0351aa5fbc1dd6d7be9633488e78f11273f02645c308182b60de5d08a4a7ac902612b3c767c5ab32736960f22fe904bb2933c1d9616bc4a37257d3144d7ed169877041b0fb84ac0010bba08d0669e7f1aa53eec70f3af3952466ba9c74a1fddb5edf12f1cf107e4a3ef0f3bd0b0a6f34bc9ef289b0e5c72c82729d89c9e7a6eab9d711b605c8456dc7c302b58ac495e56f6d0605c63b3adfdf5555a49d8d8c54e6e75b03d40a645e4d78aeface3ee381b774ef8033c2b5bf116e1d97f1ae5310f0060bfa4a18f947c7d1533840e4fa1fbd9f2a4e44155c9cc094135128aa9b7d2cbb8c35363f6ea960f02958d030af55c3001b3e6d4487a451a3e53efaf23743c5e6628efb09036fea411ce5808daee6d2497f32e05e55bbe07c708f89492d2468ed0eac08897d46ee96f6e2da7b8abada0d3535ccfb3b5bba0286cfaa9a44db3c0537b1c0c4da18f22afbf474b908031ad610aafda82c4be7256f7c2df0e6477c3e89a9dc1e485a1606b7029add2665b4a4b708bf9a3afc7718d94eb3f85053e19d977b39e71bebbc7a789f50f32a3c2ae298229056c75effb471ed8a73a352db7bd92d6696643abf14585ae799c2bd6ebd55a7eaf259cd21c1c1745952db3de4d22b94edd8214bcc2fc2b2ae8dd19cb94b5b1564ba2b9607f94423da0953ed612ccc6720e5157e34277aa3f125b251089e192279f98edcc1f639c8ee024518bc83f7940c884f0099455398caab8e9f599120b2ccc2198a7e6c4bba065c4550c07d11a96274cdaf09a335521e929211802107b03b3a134d569b17aef97e84c65ef1195f1a083e996ba9a513a2a89c01620506eb9ba40919a0333c68aec4ebfb0da039b76585be108d3a0a64b6bfffd0fe4191811056401ec8057d6acb21bbd98cb014c3ae5047ac9ca370886e6a273d0b635acdf37d56f01b4f502922fe2666b781ce522c9f05c11a842740e99c5ce6baac9680465c45963ccbd6687393f2f9d7e94095dddbbf1a11566ab40f0a0f424429c94e83d5917b1d858d858a86345a3f6aba2a26dc6510def963a2c8680628610831b8916950f594a2825b691583f711cecbb19b0894f76f69c0321ab374e5d07aed84a0912c6f6ca673a9ecebb774a0de0ef13b22b20cc9f02d3d81239d56bc25c0d56c28a0a44559559d1cd8eb7b8dc0f0102618d288b2582e0a20fbd7bac1c93469049cedf2f8290755227ff1fdc28c94f65abce0de6941802c6876ee2272b3d0fce28ee217fa925e431d365da8ecd0c6b2c6a12a5b315f375d5541c0d9c5271bdf1ef8600114f27db81656f574095ae7d72285c88403452ea2bc00c8db40373c30bbbb2dc512091ecd8a0ba66ac87f221f13b48fb671a2e331b5a3b67e6236a30e2eec2dee1c96564f57bf58fb256fa8a45ef3cf905e2fe142c14342e6732157ded374fadfdb343f4e1339cfd7ffa5b84647b774c8fa23bbc5fa552a0b9cc3ace41f85f113fa465e5638e0051346e267fcc6f220b5c4c2e079e84ed2643254d6414647590553aa12123df2f7feab81c344f44706909d8879162b9c5cb8b7587de9f79082f08d90d4a664dd5b2c36716cfc5075195e742e71ec5b208aa88b875afeebfaaed0aa9d64f9656064379d4cf38301eee6f2211a3b2f35f6029727e2b2c8ad13de4fa99ae22fd4d1f4577cd14105723bc148f90e9aaeefe2caad8028110a7226dc134a296d235e5ec7284dc8e313f60ba9ac8921f900f6235ddc322a06ae49b137ead2d19208be3dfdd7fda5dd56dfa4ce97d0c5e625d6429bcd2225ad27397d808cad132a39b8555d702fc50812e5763e69723865fe516781507823a0664ab8bd4f1d6d0e122f091677cbf616c338110694b3b196c1c7d76f5ae1bf2c9f80ac86f82a1cf9eaab1a4d97a7534435a783a49fd2456c7986bffa5e58c9bbb343107c07609909aca4fbd898fd437c3fe072d625c0a0a044a45365b785ead535a73f97a748bd9bd932a9e4426056f07b54c626b94462bcf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'ha5a69f33dc49e4e419ca3ef914bc73f50ae87fa008e3cab925d96dcdb4ff8a014cf3325dd39f55f5d1aff300e2ec2853f7c8e8957bb0213d44944e0887306fce1ed33d4fddc6bc5f5a7bea8c91a0e0ae008d5649b6a3de8f83cfd25d7a23ca543df71f4564e942d8b732037ed02a9ea3a209bb837fd1895be94eb2580c62caef24465c93bcceb7756ed3c670cdee0a284b8eba7bab0bc96180ba0485cfbf2b691a24b2a2639040f60e1b91e1a5a59e52e10da78bf607e3809c783dd90919cf90db0f3440f43495f86a1b24b9fe00fba71e64ebcd566df197ec1b7382bb011323f7030c6a7e8400a64d7d5f5fa627ca812d589621dd36d82b636ffeecdb31b056a98ccdbd097b8393a196a834a204dad9076110223e82315fe1931b0dc4abffe7c5a00e3ee8cad62c2bba8ad7bff0f39df6810e37cf98e2dabeeb29754aa31ec3e88d1c5d4af5c0f8f3645bdf5dec403589eb3617ab3b1b9aa65bc1f97a7bcd99e38f52d2116c08b05e874b1b1caca5d10a485d7ad5891793ae8a113bf055eafbb3de2f8df5834a407e8a05a9d068b2876f4f9491cbdb5fc425c0acd8ec0cab258116db205b4f22961f3f3b349f8cfc103ea0f76533cdceab1468552b9babee231917b0c5a4407e46b6c514a0a38ae39200de2cc497f35c80360f279ae933c386bbccda8709a85f18f2793076ea4a8ce74ae7c055a398841d8a3985dbbd6d5663489d233a64a40cb5b46d4f1ce578d5f8ffaa520d0e5d7afd3c052915fd5cf7e826fda650a0607060f8b7cb53a5b2f9c478369a099ac9c8f05c331e66e23c7d9e597e9db0cb7f0cfa1ce1eb5b2403f5e55e520bad927d02f9d5b47536b21de0e89fd9a8fc562857a803eccaba3d09655978aa7e4fad61c92c2c246e3ca069a11f27b827be3451174b50756df7cdff4e73a071fafcd6dce5827ecdd8012190c00fc35e43ac37c226c14727c6d07820afeb2c736dfc1901431dbe41179c45d5a60f24fbfb819941bfa4b89b15e2e08755d36fe390ee3255d2a65db3991e3afb27e50fa6e6defc2201933d565ea078df00c4d3dc9e19cd3fa9491b1d9cf289cc0d091b42685b568b4d6ea9cf4290e2ef19ca16493bca92b045d6cc338e8244cb30ee5deea8dd8fc4c79305ead08552e93efa836a916f6baf64c100fed7feda59512cd90dbbb3f39b4501ea937301ca5fa051ca74e049209c1553c7c89d1d3639fb71cb248624dc2d1caa740a3c63499a0bb595a4a22c100e54de8ba3f111a4fe8d1704e4252e0e8fcb7b05a4a2524170d7ca4058dec8d4a614d60cfc320a3c54b1f6bfacd923b76da83f2b57b762d7b0ef6cfd5909291623159982e4bd182b1c5a7c9d89f12daf172f676fb262f6215eeefba80ac81db37a48d8b334ce4025f2e66126ac0395edc73038463a5cb57d1e7fad0c3ac773e42d129d39f8a09dacd862bfcb9620261f2a135c452070b304622f0744fb20f323aed22451a30f37ff0efa10541aa23f20b39d7501e0def745f37768be3dce78fbdfeb4018514ab911a7f1e2dbe583e8dcf2240f66b3c7e3bd13e0a7ee80356952fe0ba649c07fcd35111c3a76777f4cf8f48885c84f7548398e73389e7c52259e80a9f60acde0f9ba0fd3f2ec55cca781da9536c4acece5f152801da908cb0bb81b90881665c421f5598606d09da24fc7b776cb3d4be5adfa1f34446fd6393c3c6b472ee1b064b601e7ae0b974a51d141454f369b55ab430a5edef459b86f0b2e309addedd230c8058258ff75725f74e15fdceecef59dd9152af1284f4c7c8d2b2095d6332f2159b9650cce2f3941d9e1899572f0b24f7c55f3c49fabc7ab0881c43aa976a7917bdbdb367b387de57961a5c4f4fcaa7913912c32577eddee3b5a45d5632277af2d81a9ca0b252348debd0baad4114c5d187195e4a09e3d0e558e3c7761ea7315ccd640a7766beb42a4b120e923f0150d87b40b83342729d238d6a22ecd31e380be1760702df31d44478dba835ef57a054ae9566fbe6155ac58ddc10190cba52a007752ae79ef2726c31c2f70ee2f42c7e1ef1f37c0e4206a14bdafa7bcea7095af3d7ae77c3bf5e9a833cadd60fbfbbeb72c15dd6a58addb1b4798274243561d76342d4e25124eab66ded1a4ec46b8d0631005e63dc1b17057e8936e9a9719f1692d209839eb14e36a3a6963bcef6c3aef4d496aacdb496c61454ba8435304aa00c69c7f36801768a9ca2cf50c1beb28580bf7a16372dd1791d55ae0610a8b61a98591bc07226a9bcdbbe921a6ab781d7a8f6541a3797730ae89389de5d8139adcdcb895823867cba38c439ffe77685a422c391eefad55b65feaa221b7feb27756cd3875825b9b0d3b6309284f52fbb1d39c9c8835f5e3f2cd061cc82d697a7225d39c61c606079cdafd4fb96e2a5c6e4789cfc39fb58bf137a76b649802b6838a37edf87cb5684ea4648f0ccc33d60ba41eb8fa3e36f6815191016efc96f1e4a7e49af80e15292ddc3c885ecc1176e855ebad10b2a3a1f8a7747d60fc121dcefa6d44a597148e7302a3daff3c92b9266f51923925fcfc4a30c927f102a212013d8d19333be307bcf501c1285a3aab54c20a3aea21297583193cf21cad98687482c9a1ada5a38d0bd8682a95d71f8331da555e17a8939f52eb5463405ff77cae10d580e08c756bb3e0c7619423476dea48c0584d0013545e37142b010160ae50cea033155064fd5fb4ffa18b26ac8c0f01a60667eb70b2f6537d8f6dcf8ecc0d8a887a8dc4df47ab2ae44834560e9e28c77b447a1855043f2e27db54acfc4811daa3461e5c7168d64625323c6d6c26f1e807cb27cb16f453d73289c950af84711e805a83042a5bca056cd928f7650d1a3bb7ee6a225140f03e63c04a893cc500eaec840092;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'haef2b77e57ce087b1513bd66f2500049cb8335ba1bed643f2ca749529cc2abe40fd99a8425dbfedda29e9a715aa8f0944a02d29d5221c424a593c4327cb4e018c026a0d1fd280ba50c082870feabfc6263844b21f4943e39c3995d7102581be9d0d174f095a2dbcc8b74ee6a1db413073fcd82e0a6bc02330d2e6b3360b45153f8f57765ae158687787574638e0cafc006ea03ace6f9015ef3fe00e623bdcf93c25178fc66fa3ac82b5ea22331cca715bcbd9fd29122cdaf23fdb0e46d0505ee2997753782dcd820870e227da6643f6f377c84f4de9a0766f1b0168179aef8e32fe6d55beab2651b69a900647d55884924c1f76a7c129ab0994d037526c3846309296c9c3a1e55ed0bf66eb1eef68a5552bcc7a246bc0659c5ce820167a204e3196aa168c1be926a1034badd019ee3649fc691decb39ce0e89d671cfde30592ae023560feabcfaa6ecfec9e71c68357350bda131b7056ded4e8c155f2edcd610a644268c659775c6a8cf5d686b57bdabe544a4f852e5763004106fd4c78d186a25b395cfde769f17e8b52d71e264fbfce55688d0ef6ddf82b172d7823bd461db7e493e56785508237d927b1d4eab03376f024a9d57b99f4dbb575635d3b33ba6c353781a8b4ba87a0c7d82082d4d8cf307b60d33587ca4d9fdc319580933413adc10fde0db201ef3cd030a930dd71f9aa90a815fb8bc38b68a445feadb75395c2f0f90712294cea5105cf1571e2e424a8dd4bcf5255d6d2990d851056e75c4df7e87b4012e55db24c03cb09763e1e1d01a99812b31feab7f0e0ff35b7817608da157cb485764fcc92bfade39ccdb976efa6a4cbb35191b896639381b52072a6179ecdf2799dbda8b79a14d325a5758de0fc4281b61f48f095ebb442548f2496d1570d1eb3bd5637572c338f8023f1ad45f49b7b12bb4a2897eaa5b6abdce18168d384df2d75eb3ca7209f794fffef73a40cfa1ff96f02d7239a12c9d711e0995ba358194d51f4b06577326ed7e815cba2fd9322950dea83a9e77d53284da9575e77acc1315d6ee879bc943e8c9ffc1d98e123541bf6e8002166b965757e9e1cc582d1d6d6556c0a83c9a71d56e299bdbcd402389c74d2933180d5f374717bf67661dc43fda69a50efa0f6ff6b5140e9795ed1b7211fa7a1286722d9df194988ca5590198590e256e124debbb933e9a2d3cbd1e2161f83dcf3274795783ff4a72cb0849a4d7a6a16511617432c23fd8fb0e20063ebd62c2898635d728b146fab2d20c26c09fbd463f7e6bace6c724258fe8bf1569c45209aa48eb94782bc375411e4b75d4706fbac5aec7cbed24ca248a9ed4e870be11757378dd82360b7304c0414a021e2e306fc9eced1f222b3b067e4d2a85c4707977dec27db50c2a8d2a84e9d33f128c4c72cc1d93d419f3ef9d02660bee8dfeb91360c1265bc8d7723b7ce89d992f8fafdb9c0181f03277c5b839748e9dd8e5a88731c186dd0c24941c4d7f6959ae3f8c358e684117124956d3afaf2fb5b414127274fe2c2dccf8b85b97368d81bf0fe58d40830a149e3050fa6f6f9f9f62bae1df4136580662ed8b4182af08d980df0f3b622c81ba3515c4552678f4db470178a2f58fb8baa2df674d8983130e7a0a43aa420ed1c4c59c403e9aaf8283b9ae1b2265291e3069f3edc53ad5ddef89f49a259844cf3166f772c7b92dfc1491a170fead06d5bbeb0681ca23cc12177fe029b21e54f2beeb0b08bced84730472e30aba24d0b63d0b360269059f4ed2d9ddb349b941625f178a2b555b73d0db53deebefc487be2b096f93f989d257708916e821aa7396e44377d7878dfe6d70d83d1345d221f76a5c5e3151cb37f40f9d72399c567b370f610cda43bb8aeeff9a85b4c717a9aef52cf27fc1761a67f4c01d242b9c1b1d63e9bf77b07f0a967ca19806534514bf3a7f95aacbbd2fc028a1c61168b8ac41b6513ac2beaa677f556ece5545f45ce1281ce27aee5dcab96e62c04858459f7a06a32e0a5f8ca955b1523bf47d8e1cbd268657f83e49eb7a1ecc0f7cbe0361c16768941cc8d218e2981a04365b65e3db32264b0783504800e4bc6ac13840cd3bea4845093e9c3f1115100f768d526b3f72301695b888daf513269bb013000ef59372325033c2983812c698f7ed7dfd91be94e2eb64dd5b978ffe261939a1be2884385992bb6364fe6e0d3473bf3e98ab7e372d2ce1b2d7a5086efe1cb3af9a6c6315292299bd883029f6c6c2f0273732ab270e78d942f1d76f71a97c546778a53ba7b5bbf89096b448c81d799bb75fc16cd8e091f6448b5b8597e8330bb3447c834c89595c6a57481c089b352149898dd2632412dcdbcf1c245987cefb30aa7b525161f669405b7166dd1e9f9be5f670057f82305bd4fec8f3a0f0a12a7b73bc51b04a781d819aed83bd94b70280f4203977af2874ff154b08ef6df7095030741ca5b8cb11f53ebccfd3f1419ba273890997eb559ff604d4be821c53e865d0bec0cdec5ae871cffded0ad3cb47c61b95eef2d53537ce802edbc196783123c3b3772ccfbfbd57ae617f6bc3791a0bc0ad5eeadc55897f7fb258d3a718cb60ece68e02e7b8206f2d2b9143cd1923534ab31a6877dad2d280ba34cbd7514ca383a7671c368164c4f0b911431b8e4415e9304432812de99b307c47826403373773f48900a3e7dd5eadc0c353f495ad542cba104c6040223df8e1485ac6c172df20eeedaf617150477231f780998249f2f8bd77ff601b5962e7de15dda352f4e3e46548ede74cfb7816874e07b11560fa1e5ef17cfbd3103492331d649847c1a127927446a361beae13c38e7ff9b4fb54655c163c560fd009c97d826243da7c37c61d9af5a1ec17c0aa6319ded66ce2167945d4f199c3c418;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hc68e8b54a4678d4ea7eb44887b9f985d82ad186ff9ee6a2d19d87bba53902d3884e2feba5b1e50df6c4363662f3f9367cd7ecdd1f314bdceaca82acbb75763463a13bb47dffdaccd73500614da75e07f698a2e8243a5e920a1ce9e5ec7e69831b2705ac1e2098668412ed4942becb54a7ea8d2246b8db8a895163412a76c7decdc79bae4f0f71ca63c1f9213264fa9042d29649be620fc85300a82c94b8849037ebd1232e47d6053d0c11cc14fa4cc961c7db3411c8bc013f74c87097992fb92f2db8356025863e72127e8c19e011f9fc9ffa7a3b8cfd31c1be0032ccc49266fcebdd43791e50f5dcfbc792f0c27d8446f18b91b38ebb23c879596ec270d3a29c13a24f716fe8e86e0bfe4659fd35aa772daf481b83111d306f402ba20f511ce5dab84566d558ddb3b00e7998dbeeb2811198a3b175644e00085677dce50ac3c2b15b8911c15d6484703f3f9625c49a7c4d9e3de761c7df69ffd26cd5b9c5b42cb843c4f7506503e057ac6040f77f98f31d34666d6258ed0365e95fa2514330bfba85a6a534079b77e1dcac56a4669da3d5f69623aee63ad42c3bbd76c91b7bd07bc074aea3bbdf3fbe009035d0106b21674afec36906a0384b6b83bcba3b78eadc3dd8bcbb5c2e62e69128a613bcfff35c30ff86929a490b6a3a11d98b1f79d1f131e7c1be906b89dfa8400c2a52589c484b1ecf3f0d9d080fdcbfa266f4dc094f421e56be9a1ebdeda34224488a910a9b22b4655c9bf6ba63add428887ab3aa5a8482223ceba48392187e97c698c841256b47ca7fcca1b652fdc22a674f9f6263953c7b352a7ce5d87dddbdda2c80e8ef3447a9a4527cf15bfa9be3151ee8e9c87a6a1557c42c58e1f77e4684605573191f678a7010920f90e7d27c4c424cca5d403263547a1d36709ae8cbaf179e60bf5047dbce8047e9c32d66ce21f53a0fa3c1cab8fcf42fe7543a09432c2b44753854a77eda07bd4b43f04d38b8ed51be07c52ddadb2f0aa69e53539acd5359c070ef684eb2a00f64c54f54e0edc72e094f66d434cd5e12a67c5146bb39085101fed2cddc22c0d8afa08d09f56d9f6aa5b5101b9489f47a379cb80b43fca0c9fae4ce303d031084c581096a7621e09b84395b77f6ec98624e69627172c32d353953cb4aefead91dd04f60e0aa041f141e6827ae3090a6e0f383f6e2282d6bed7121046e71fb5756865a33398e6ba8cfdbd93b723c995f6819f81c49c9bb2fad88c5a57f995bdb69f30ba0ec4c286b035d001c954b9c19f20d350ceda51c2b13759293d47be626bce176d48407b587d381037a3b384ab4e9a9425749d47a9e09859c62406fe34fdbe683b840989378ecdfc901f424936993ca4978afd08e1e225f3944b0c130d18cf0ce9b8f941d35e00f290490c55cbac293fd16ebf4b63391cf4494460072ec6cf37248d8979dd900d2adbe5bb8d790b080c8c501d8e41b370e1f65ce9b40ebe80608cc4534db42a059afee2a7761f78aec06d81bfea4698bb1a4fa17eef2593fbe6629ac8ca8fce3259ebc6a14de8a940b0fa9d1b38207ebefe38ddf5e533e93d0d0c63658a994324194d606f22c5f78d44fd2837e7a22991d281e785b9d7adebc455d2d52a16a1f897a13dd134358b2c0114aeaf51811a91be61b297d19d321dfa8ecec185db78a8097c3d434289b54682b07e60033c548eeff137f8bde5afec2a6b55bc1a1d21701fc258b985dd7ab0767f85dfa121d2f1d4e5ec87a42954a11029c68aa56bf3ff07aadeb04a81967830dc73b4038b1eb9172d9a0de577f750e0af06f623f31c0f0666b7f48b8eaa1266437c659f65e6dbd1527777b6495f294b3ef2bd05a6253d157890e5dd01e1c6eefa1145e5346e3c3d2693bb40fbe56d36f05604dd02c47d8579537c248f803eb4cc8bf92ac3a2ae638d8ed29d8ee68c07ed407360cb78935673dd7a4d012e9802699a0163b841061f97dccb66affb1b4e4412e634337996db5449c20ea0e73d37f8ca048c9b374a2da6d4e29619ec5f65870ff9345021b72cdf88e36b454e4e29759ac1806fd6fc0592b33c4ffea393f86bfe243246754df52447c4434c81fd6a24ee6922c0c69f4e7d22ee2586e4efa986cf84181e593b02c8c6b21b4f257d22fa5bd678508f25c31ec09d438c4cb55925b3a7085065f7b5a4bf4fa7f1c4bdbb9efa7b647842539ce9dd6b636a59697f8019416bdbb0bf5fdb03d6198fdbb884fdbaa57430364dc82c4dfd374abfb132dc44ef869d137ad4c970ecf9cdd6b3b6eec683c85a8f7f539b2223c592f00238161418ad8c7c3eb7c8902801dbaf93e23ccaef5cfe5c2db76e3390f8c63542a729453cf40648bce0b28ed3f2d1df15dce76af2491989ae533fc6c9f74077b9edcc2e83d1624d6ad4048cbcb3d82485d05e292cf51f50162158becc86eb2c052175b16ea3ffd12d29d5fe9b6ed46447efab9eaf8b452a6fe8fc402ed0c98787a5949fe328808b6097b0f0a1cfd100ce622becde0883d08f9acb352b3b83a5e902935b06b2bf3c02366e29511830d884f216fa3d94a88aa5491bef89ab3cd72151effbab99cc8e13ed5e19d9a227927c851ea2cca7bc27958645e7c2fc5945fcd5e1cfb31c61483e1c8a20785a7aeb4cf9888532c606128e75342d14a3ac60692661a5e3a07abc3f9e1dfd671c00cc052cf1a43a94983ec952ed844f730de01ce52fc441a7ba269e8263d340d749b4fcb6f9615f9a044ef7343294176aed473fba2b34ab16e85da13b182cc53c26b8dcee73ae26401577c50eecfa4fa914f457c3e323e6ecddf6970ba547de8281eca3f60bde0c6baa59781eceb42a19d4b941bb81b806c9f6d2764dcea778537f0b84ccc3b4b59f086c18cd5cbe4668955a024b318e9a6f9e2101;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h6a0ce04eb020f6ae6daf02c4154ec315845b56535d4956d4d736666d1785c06f981352e3ec5fbaf3e65803ea5adc6a2c65b671e37fb888d5e40fae5fa669bdca52db9210d4db0c58a4e6b30ea9b721b25c292a647cf5eed25022d43e9ee383d3c811cff8c18081dbe28e516fd08b3794123ce871410188cb95632f9506bae3b3654bf169bcfc45430d613c7fef8faa1b4867981cd9c7b104e5dd086eac017e448955bc46aa02e862c45e89126e099ff4f911e8c055764db6edd1de5388cd4bb5338709be4115e3ea3bc4e07cbfcc2eb1c89e225968af93edc264e1c71a16c9c53784696f5cfc9fef66a3e3a76f9132ae8a9f9daaa93d36aac359b089d8c6018d4235b41c76c58b546353021d849468e687d6997ea297ff89759ad14349d6d688f63c75db6ead36117e5209b1e8e6b9994fdc13f1cb7c8a1e7d766232c31a3c59df69f0840c812aef49c9fcb871679c0ca29d75da7888d4f3d5346fe400b7521d29e80d10593d001a4c64e7c22925867c34d0c569a2b28947ca7fdf986e2ca85f1580e94f5c60a2d940dcb3686854dcef20825ca0fa4cee595a1b15e112f8c64d99df486abbd280246930e2ceb3d985e84dde697ce175abd77ebc5058996df1d349e74cae14b92aece16190882627cd9e40e340ecf5420252d2645722fc354ff53b2045b07f1fe1bc8f53b5dce08f20ab958fe6650bb5973bc98685da4db224e66dbb1552bf800646edb98e2011975784a4a9cbc00d8400c292c9ed11e60738c3cf4bfb0482e86bdf2a1793ce29fa3074a6fb0670cc6c8bc57fea2002c04a4d9404fc6d303e336b33790fec9ba2908fecfcd70cde94cdb749978c157fb3578b4e2f5419571bf4a9302df594df0b5ebd79a20c4af681ea60a2c184474c723c6d7891ce5f457dd6de5d8e8136dde65aa66bfe3a9bbbec04ebd2a3fdf17c3ac1df35c5b9417eed72f089906d9b477b91ad0089555240fed3c97327f1af2561a328aae753f406dea791d23601e60f54ff5361cc23fc8cccd3b6e9fcabe964486cbf299118eb30ca1076ec4be116d9e913fdc298df2542aa9f2361fe82f11da91ed2cd33234fd4e1754aaa9259ab50687a19f4e946ed2e3305b1ce3f85ef970b46b96af989ac72c10cfa503b1808d0f95434ee1f9ed2d2538a47164c7f219a5ea786260705e65ccf5c450433dc6484e22c508d1ca91e835c2ece1b76001f2bc402b542148a6c4843b9d7d8ecc956681dc86436570dd9a67ad955dcc1c6d657c3f5e26e88eabfeeca58f9aca028a906f6271b06bb106f5192050fda546bded06461a6d50940e44e486fe0fff5471332285260a0c21b15fa9b6ffc7b37f7348ea63998763bea5b511a44c0ebca374802a0be0a2b4b20bd4b64a8b5719de24026d3f16d58e9404e6fa33ba0ed52ae94c564127ad7223d1979874a28ba373f8eadc33185ebdc6003dc625f87276445f3fe95eb82fc27ae3362c67f93dcc4c0a1c5e76a7a02fc7a4b11d24dc7e965f14c5e6d939216a1e62f76c112fdc8b2dbe78d9f49b6eedf9e312f97b9ed8ef3e228473699704bf7cd4cab85e73b54172a27005e7b8dc7a2148b27c6ae43b5b361a73ac92d7675d13860cd16b4e7b086f7d931ad32eeea379350ba6ef4112991accbc029954f1a29194e16fb98f487f98e6bc3032e7fe075d74d4dfd6b2c554e5b123c127a0b270a8e627239fe21e502e95fd5a5d71e77e3a3a9d34ac3b3cc8a1650da3a429b80b44f651bdd782b620a1e9c59ad345d9a9ef4959aa88be58a15320c1513a04b137678bbdded6dad844789e3d59565ceddac4cd317ffe1c24f2d8aa74459b345519ff9df9ef5ca1a05be5aee0ade832f3f27c58e8a37ccc22c561b6f777eb0d8c990ec71cb38020b61628dbf86332bda7f418435b815f7bc741030b33576d5afde18f899ff06c9d781b074b1eb2738259d6952063550e38345134e96c905e8a80f73d2aaf88502dc5ec97cf10f8427fa8cdc1d06e8f2b8afee195ba94c9855c6eae381e70611b0b8919db24d75bae9bcf586d1f759cf3b99d9d41d6e0aec7d7ee82f96faba80e03eee0b7e45f11c53e8bff2f9b5cb2090d7e5b464721dd64e09bcd9b3896ef85e8f4075633bbb4ec444455ffd75f578d239e21c98a9bc39bbbb9de2bb069e5ea93b4d7646ada22d23d8ef50bed82b12b52c7f375771f22ec4a0662c98e54f833f1c5698c8e85298feb3d884e63178f51a7c71286bdaae5e665e1afcc1f1ed6849ce19c5cc300992218819380919f08407d2435b958268f471712e2e138501ffcf7420774265971ffba78f87a2ea44eb77969daee61936ffaf902c0c8d4b6d705842b986d1988953a409fa489ed4c818794fa18a7eca5605cda47c5b16aa0989ad270096efda728adb29e9d714ac9f182fb26b09bf9a884d0a955bc0221e093cace759399727fbbb8284d49899ce3fbfbaa308172087485a6aae60aed61e966456131047faf489e5a21a324873be44bc6164e2f8c5daa762e11d6b82e7e0a5fda68167cf9e4f29269ecc7f0dd8caadc183a4bfc56c6da19b232f8921eb02d75653f04081dfa73667263bb91d8bfdb6da06cf5a46779767f89618ff1e2d9836fb221811feecbfe34561fda944919f70735854fb6475a0f4259521b5b726a037f54dc8de29fb5f706f98ab18e96c0536527c898dce7c0fde75a0135236799b2c695c2ed33f5216c1b692d11cee33051ef45af35888f8036659371a5f34440e062b7b097e7cbb6cf6e92397f8ebe3032556e261b5586a42850b285d77d54271fdd832d56788c55314619cbb958f06ca9585a086fe9e47584f3bc27606df7641c528595e3abed401f11610eedba547bad3a0ef16d0a7ad0ae28bf48a4f1b6644eaf49be19d10ab2f700e872b26;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'he7cc6448f8bbff285dcc009386ec06c2fde16004e713b4043ab38b09ca1d052dbf178358c0e0c980cb14202e5a59061c5e54077e6414d76f1f290b981e15f37c93ff3d2dc031b5930ade8fece81100b9e6cc7a86792cd26c69e5b1d79f8992d1b4bf2e1bebdedf9e0ae4ccba8a8d2c1c9a31dfbf4adcfd31601ebda361295e62d2cbd46693c0cf75f5e64390ae41b3aa0ae8602abb65a669d7a0ed5720cd1a815784e41836b301b095c724f6de1244ae2209b3c6088a3ab9ab7e14bda8ae36387ef03f19621e9b8363e620610e8edeaccffa947308c789423bc83437dabe48322a44dc75942719425ce6c05479d7a98e040cdbe2700bcfd6a66ed3b0f7071baa451c1b980c2d98bb63a354909ace435dd636aaa8c7e9de513ad809b5581519103ef73a543e2b3bea25b5b6deed6a8fdd4518c63ce6d84ec4671921d389e8d415542c1321139a7c8f54ed7af91ce28b4ac9e177de545a14b26ea08154d7c1dcdf066c50b60e8f55e801b87d60be50a214343081702d86f12b5b423f6cdb38029983cde3ceb8331070a537ffcdc3e5d3b383bc0e31c579928bf54b1a474b1b8075b57db6a84d8a75206ca58750c2083197100fcb1fbe92b36bf4aa6813cd17ad02aae608aeb2a6b39f0fc24bdbb5e4ff4485f8302bced03e53867b813cd527d471f90b4cce632147ba4532d592f3b4fc98491625956f57ac946647b5320a2f1071e11c4cede22394654941b8e0560e3645f42e9b4b54ecdca2c99e09d59aad1f56197ae0f2d3843722a8ef7903e5a75389cfa67014c5452a2ec73a19e516b71b1f7eabece1c25d2e4bb7e1ee7c1cd4d703c70d55d5d31e49c449b91c82ec6ed009111bef014a09e3fd1210435b209964cc168cb05736b4a7e5414272513244ee815ef1540f56b7f74ab4125b7f0ab836d3cd228487747e626a407aaf115f9f8626019e964c7ec9b4ad69113a305199d8efc7226ee0d21e3e913aa0c400d73a372d1fb148a21adbc23aafea094eb1e165609b28afab269a2bfe1369aa1b82e7bf7a689722b06ee792fe5252e55864e82cc27b113fd1370776ae2a06690fc0e9f854aec8146ea0c83b24052bf466b44995664f53a7fed9f547718f64a4fcbe9494c0d89266e9296150e09a561468a5715068dda4e0fe0ced5c3a336b36a88bb52cf222ef8fbca843b5806daf198232c23f7b9cbbb4feeb6df087e28a159eb7fd1370f8a67cf4d4e1766af4ce38a607cee66446618c25ffbfb857e7ede1dbd42065aa82b8d72f7597a9b180ae866d14c5c9b0f2a1bfc0a746163dfc1a33e07589914f3a75752962934e674e1d2b6531f37600f32f6308f3168cdb561168be216a1c1f26b4595877c396e659eff5e6e73d36441ecf22687aec676f1f48b0e78984529a1005354eaeaf92ed7f56e7079bb9b3070a64a3bd56e55ab78683ca5d1419965f70e69818d9baf09ead6e8e9d5debed2bb402ecc601fbbdfdd39e03cb7c931e04479bf5d7b20e282543dc335716605951deb24954f91c480c8792a94ca12319629a038303e953252ad45008af6f7950303475753f5d85efde288f4b515ab22c6eabf5a0c69d2ae41249129dc77518200c6941a1f38725cd7998f59cf4e24e088d07b805f492380f28fe9822c19a51ead62ef66373e8d871dc56e2cb72252ab21ad3b10c8c5c066ca108e1ae07311a4abd218bdc7c09e28442a6967dce6b382bc2b2eb4b5e8039c3113ddd247d4723c9f7ecb91a49d1fc3c161d85f75da6f71050a3899ba3b1ab3b98145b9d392465b2962d47c212487ead9ce12867758fbd039e45448131607d549860647842fe8096d64d535e74029a8ce168e09617b63045059b0a5668b631b8711c4dac7accd53b4ff18a135fd2246e1e2a2dc31e1662c5a1a3f7fc535dfde54f66b3e7d0afd856aa896d8cd973450b24d672bc519ef34bbe70549a1f7a82bfa22601dade416ab3f2f589345bbb2bea44f6cf90bf3214095b60b86c332935a85186074af8bd9ca9ecf0131b467e88aca9d3be6c2585dc388283f957ee5c647622e0cade5a71bbabdc739261eea62b9dc6ba002feb8fd1be0decc7e99021d9906b3db06c2e6f1c028edafec6e22f8a996e08252427f605bf8d4b91a432a72d8f6f85d819bd188f4e7116c038fc5fb13c0100bba235148e49fc8496b8fc0973857bc35457f0cf49b0592452e51490e8fb622cf97b75e4d4667c0082315c949ae81ef46d5bc351bfb1bed66469516ecd749d12076b8222ab49b1a629cd56a3be13a3e4eacd4fc312fc8dd7cafacdcfe707c959b49b7a9f9e924f70b895d1df1bd6d4a0302ddacfa7ea274bd5ce5d53d0800280961d02716ff089bbac0b9feee5b4201eedd907f32652ad61e29fb6390948aa91ff451ed8276ad9fc6b8bd40b625dd5dc2d3fee13b313b992f94382ea625ca3f4bb298c11b9eccbc75e315a1ec177c2899dab80dc3e68ece01ec20a95a4e7b3bdeff6fd3a587ec2f2a859d311b86ee046e741e10087dccf648f808eebef60449d2c12705768a9b31384f2cbacc33e2be2daec3c5a53a78fd7c75050247a34f74e5efc0712f6fd6a892e72073eb9855c1f96f32131d3484567ac2d8ee4c8f1c59678a205d2bfdd5389e207789d7c6a744240cc03cec9245da058d96fdef93418f2d0f9e230206dd1e3438a25c18796471eda46af78959e2296b69ed9d7b93f0ded132cad64dd6c7691f37ef6019493195a684501010ece8bd81328eb6ff53cbcb152dcb3b063666293c3cfa529f020d6f16ca1d8643741078a8c4efb9668912b7225eacd5aba96fcc9f4b0fbaac5491aed861117837457862206b30a0ba58860c9fb233a86347360f20973c9b0e994bad35e9ca36fd39ea7ab4c68f8e8d1e4904b9a0f524927bfd5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'hfcc5e2e5c475cc1348f4891efde2bef3db8d1da0a50cba42b3a8f6789bf5743a55be3648935a4edab8e52ff6a5baf8739cf359b291b2cff8f5be79ac0cf64c93970ae10195757db4eb9505bc9e3122298c411168bfc4af69a9aed36a7fb13281cbef0063381c4fd3ba0384cc8174aaee835e89ae7cb3c35023c1554f145ab29e1da8d61806b04157ab676b975efb2e62538e80dfeddf260470b86faeb19e7054beb849c0b1b6a33b34470731cbb4b23e9899ac0fca6a397442d5797f8a92860aedcb07d2873cba0317e802cbd5951810b4c06d6f86284c674f802f6c4171954631375293992adac2accfe57e90c7d7a1960b97a9bc44dcfd357689fd8238b817768a44d9fb16e5ab7e225d285666a5541f408163ff5feefbf53ff6a87419c4b77dd3a23720623949047e24c2289f60c2b924d5cb350e91b7d7fd3861b25fe46f6e25d12ca104694f41d2e19b3129a45b79c106b22c90ccedeaeea9b05da9297123fa562557cddcde9d0273ed363c92991e2c22a4da7bce759e9eb9cd099aae3080b558d4573727c7b8393c87b108ff7c62c50d3d817ae5bf31e2ef90ae47fb4e2f68a951ac9be2a657c0ea3a3f185fdce3438988bf1e570948a0ff84e99494e8debeb6814f8ab67aa72fd09b5141d74e630e209fa7a0de04560312e49085745917f710232a4c81c572e0b118b4fd6a7a106a42e0a92a14483becc883e5be7c0c79434db3c28a664a76e020e987f990e0dbd38b00f65472088352e39bfd6d65f1fa6ba5a14f464bb59e88d9690e64882aca419fa16d1835840b08888b274cf2fea7f4411095d06f69b70ff9d894dfbdd5f90ba88aa49bfcf3e6e0c9af09de45a9cadd72f75f77f8f0c398766cdf6bfd188d4ae7af5a1614030ba3b677704e8ca281a7c3b4c0811ad29f246816ab4dab57a7830df27f0e866f9b43a3624c432fbffaf8774131013da27e110b3ecc212d66c28e6ec63fe1bf65370af9203fd12caeed46ba973e665ea9c29f16951af35c6088ffbc5c4b2bd0a4e64e1e7abe03cf5c96bd47cdc2c9bf84829e33eccecf89e0ff49e31c7b6f89e9206047a1e484ec8f53112a10c44afa9747b233d6aa7ac8873478058a481f9d6e0a67230f5dc9ac8c9c56bffd9ab317b673d74dd8e9f9e790a4ba9a8880708acb860158e55f938731e6cb67dcc015145951756f33b103f020b95bc4b7b583d23e40ac15c10c792c8d0cccc5387d5399de2ecbf1f5681e457d74fc94973f51ca544ee28109d95a42e63e67896c08d9ea9bff5e18cb0d834d21280d09eec65a9e7e3cc159e92439fbd17dd3c82b0f49a4aa57f618091e53dc624575c7cd7756511555ebe2178b38dee60bda61511a16f8e7c8e5d6772eeb11e8360935dfabe4d23c43340f175b6808b399ad13d994199f2764d114d517d64634bafa7b9d6f3febd515dedee5c922abe4c8ca633ee8a71b2877388f7072eff11c9b1dc5e51f451ab30e7d5564787f0ae19e5f8a36ce6bf79124d30b46825ff88f6f7fa5804b299c89654ac9b77eece3bd5e4c928842198bffae751f5e05e22c98efbd0062327333fd7d1fda810792930fb8feb1e59ad8101d61560afc1766b0098f6547f114677dc8694b8cc4628627b0a80deaa25ce22145916f6900e9d02e5bcc6bf1c533366d03488a61a9c6088b6b81b111cc5599e27122d0d429336576ba8fdb8d86d60d5c1d1d800daf2384fa85e64ec39b3eff22a21c170b8a6d5854fd0d03bff94a1e5ccf69972b36c0e59b6da39b2e15ea30ae5b65dd0ba3d77141d52cbce6f0fafa53358e35e88e6b3dee9727dc0086911994271179b28188c6db7195b2b5a9dabf86653a28a33588b2ae94456448d47fb494a492c604408e350fd17a064986252ec2afc1ab4010821e031c7bb38560c99f5c559e48f38a6b7a7fe09b6556d98e6be14a4480e81da4b853d13dd01e98c073aecc180ae5c5f409172f14bb612eaf6283eb0f44ff35a11eca4cb74cb3ef1016e81510d01cd8928250170aae6f212a8f02c80fff32ea7526c17a483f4fded646e5ba4ca3d5214dfabe9f4df86fa78a44e074074fd20a5fbb277f5fc4ab878f846573ad6d3671bab53bb74e7731259cc4997a481100d74c65a6b2f35ff5236ab72e9020e9d1e5c99320b2c3b61750806e6d8029023e18019cbd4a0f1c3f65e2548f76621f569a90f4abb479d0e4936ee5c667252b5af127cd7ffc8e4eb3018d23126b57410da9116bb19c0fa21feb400a382c3f082400695296791bb02d1d2ee06a4b304df511e236746f2b1b9330800700be2a9c2c2818e0ef280f7137139e49d0d5489a7ac69d91cfaacd65608e94d367064c66fc9a1dd9f52e681eb288a75889e00f0e4cb9220df1eb9cd7b5362e66e351e994997a55d4c8e4f96170ee22fd1513d2ba666d48a17fde6c63efb438b423a9334ff30d46f392843909389282df18fa53669b0da61035b5be4072fd9468db0dd34e4f308b25ccc515332660059fea1d42cf48c39058588350e673fe92311b57880beac6f177cd4800755d2098b8ce410aa08bdaf1f9ce48464cb562fa64da5294de4b27f774094777a1d9ae0cba777f4821e324be69ed6389ea3383412b8b724bfad9096f00717fba7b5b8a49390dff2ff3e15a0f1ef7e607fe5dbb192b2803f05cf24b048cf0822362b3985ffdcb0473c3ee95f99017333ed8e42df1a61b4951a00bf475b8f630d5a9a760685a6ac8df96656fc40dcd33854192ed2e54ad724aabc30af195be66c1d951f0a5a732fc44b4b8dcd00c0335b548295f6bd92326b64fda906df9a9842527e2ead829a9499d80c2996d72bec33f3e7250af27d2eff3a2bb5b611e79184c08782f6284ab67e1d89131ebc22dcffd27834f469a46b191026e45257fea1b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 16384'h9f5b7c94246ea26273e32d574b9e5caa3055b15438b19caa8df1a4603313eb3726928e12ea5a17163c9b7879441c32b3f7a51c99a09e29b2aac3ce5ae4dd1b809760a88dab1b61b78470a6e953dfeb7a5e5125cf426374b0dc0b3554e1e58038a089875079a876d930fa7b262d16eac6389c32760121e406ce8ca0c08449d037d1951757ad1fda24fed967e570bcd3f2bb88b3ba75605611ee19e311f8691a4c84bdb884811c16a1143fafdc4a92745c635728fbf2f0009bebf1db957c45f76a7be33ad5e2ea03cf2fdcde46373a66c1d99560a21f9bb6eb5daec57b2c1ae0b74d7c1225ecbcfb347889e624bd693987c30e8802ce50677d0052c4c44a8b7cd9fcae47d430bf8336fa94c9c16a3e5c7c2cc7bed8c9a0b228330812f3266420cb152ea31f8d5edcffe5376d9cd8f87a5bfaccb90a27b1db9f641ded9de7fbca828d9e57d9c64a453e47eaa19a8c5c02d180f5694c4f75ab7accfd839e42f9a6ce8151cd7fe9a2a709d2296f1f07e27d1929d6bef6d291624ef7ec0ac26d3748ef0cf83966f4feacbb9280c9de61e7dcafa19a448531d7a22607081e31a8042d16b413db247cd21ba08139526a3444430c44ed36323fa39d0e8a73ade403b0185921138036c81a4e4116d40b236525f8bc6d7ae68820b95da4ae1cf068438773647c21bf1b26425fcfe5c80a47aa7673e59c61b78bb96f3517bac7a525d87ad11a05b1495e40fef8476fb4ea564699122104cc020f06e8c4b2f7a58f7d4941ca971be44c779a0305283c24e9efda6a8a179d6641bedbae8c53c9d5b03c4ab3b184c999414b47f5a19392e50a327a73fba88797204476e6510891c8f2807632c68aaaedf7e9c97c9f27d215e3344217cc5808dbb8c889114e5cbb1f0224fcff62fdaa5ef232a38c1661b2c8bea30d77344a1f9380e3a94dd8ea92ee8a6ba6fe675042215bd7a2f3ff615f983a6fd5bf1eb99b1ad349e2030eb9f3c9bf77cb4952596c424996a3ed00c81c38d616e4124038b977741ef9733d861b3bfb4a7d925c526faf7fca4dbb21c657bb61f7ee3bd547965155303347a9e35cec0aefeb1f0a53dcf51dfe40b86a64aa79ae4de02d950e0f934909d51cef7d3872aef6f3aba7ac41708908bd92dc4f4ea763f98d1263f29602e450ab5d92202233c27ea3652a79fa220fccc7339d305dd25589326a067351def2a76b3bba9082a0b59fb221c415fbfc70bfaf43a2aed29b6ba8e56c3cd647a2ee05ba4fbc7671ae439d326112b57cd2fb8b30248b2bb1a47dc9070a43862ceadec414489709a949508a413fa9c07326c06eb89400016b11399b671ea25e53303d5cc15011390de8dac449bba01d22178ad4e77ce621e59559a4a6f5a4892552a8311d48b6f84bdba9c5870c972816b9c42f117612d80658c5d78f69f5006f7b3a47ec87ac0aab8180ed4ac5f4e5c1f1e042fd256d10e8e3d8e6f1a9778fffc2b016da785b0f409006eab8d38b4f1ec0b7a41c1d4febecec3bf9d133cfcb08da7ddf7a3cb29d90a47db5d0547843a60fe93fb35437554a0027b04f73926a99da6d3223f2dd9f1dcab7dd34d7c8273c42499f7492486e7c96f40de3ef7f6dc299241cbd72d3350306a1731c90cffb9dc3a34431aadd98beb60e21d9bdc2cfbaacfb446a32f9fbb10a8e457895f2d10f180a542c7515d5c8a62d03abc903200c3f182bde986fdb50eaf32d00bdc530b09038b0fbe71cb9e12f866ea7350332876cb1ab83373a688afc7498653d69495c090a385b736bf2299c3832afbb08d72bf0890c5519ad57a98077c5bba89bfa0e2d1b85e7b5dd4a8d57d93250d09d559bef5d55178888c349d685d2f00d5e0339065c94f978264f4c3f45fbf2f18f2ef444a09c61da995b0e908fcbe18b94542738cd0a2dba82168d9b813fb1db9cd01b6013ae57946bc641931071a1e94b38330709717f87d81af90b6140e6b33c968e618ad2584cef042862d4b2c09da60af768728890bcf14cb2f69fcdbe88047c117e8dc84ed5811ce0e07981c4d9bf80dde27247b278e19982f3aec84636f6cb3830fb7ee6bbb51617c1ca25576b7416d56ca4b584cc87ba1af09b9f54cb2c340b58be8ea88d8711f9f706ac78c9c96a47651f4b554bd97cc15a79d1212bd7e323f60dd6c2314d12910c0295e0751e4349c1e29acac3728f946e538553b27c8c30750b4e84c4a328f7a02572e39a2d5b54b0e249bd697fe8aaa4087742ecfbc0864fd8b043702a8cc5032397ec968340fda5806383cf90d93ace940d2e2b0e8f3cde7f5221536e5e0e8289b7423a27af832a9ad1a09fe040271f72926cc0759abbf02dc4bf46c25b554fd7a9f9d6f925f505a5bedc21fd6b977af5eb7673bc26945ba2fbf80b976aca6b0941ba1161d41bca1942d0ca3808eb0e6ba859dccb635cc6dd9de12152ffbe822f82fc6740987e71b63705ba2879677d2614c13c38af35ee263f1c8a3d85d3986a84ffcbb9184c7fb3fd24361c575513141d610f61516504f548f9c23b4ae2de63b7a7a43b6fb2d1d3df2d58132c81ed5e6fdd98f56832980c703087b56938903de842d14b44be8ca45cb57b4ac52bb8c935b154e903d0a98877095814424a3fc93a74f128794b65ec1479dceb1a9253478074599bb09c10a1764f71ef2c0b234d5675f99f42601591e7ccc8a1b64b81c9ebb935326e0c6a288d8e62b1ace3812be108f6447e1be96b750a95a2a1a0b6f07d8dd7b2024feb5954c80da86d568dcb9428319be73020833d75f2103b6368968f85bb4dbd90266c4bf1c667154222a35df6e7fad15c2a6365ab2ad831c5fe690740b861ea38da90586139964dda099c22e44bca1496a0282a639f739f4d04f9a460ffdaf6b69b3d332220058486a444541e14db8b;
        #1
        $finish();
    end
endmodule
