module testbench();
    reg [22:0] src0;
    reg [22:0] src1;
    reg [22:0] src2;
    reg [22:0] src3;
    reg [22:0] src4;
    reg [22:0] src5;
    reg [22:0] src6;
    reg [22:0] src7;
    reg [22:0] src8;
    reg [22:0] src9;
    reg [22:0] src10;
    reg [22:0] src11;
    reg [22:0] src12;
    reg [22:0] src13;
    reg [22:0] src14;
    reg [22:0] src15;
    reg [22:0] src16;
    reg [22:0] src17;
    reg [22:0] src18;
    reg [22:0] src19;
    reg [22:0] src20;
    reg [22:0] src21;
    reg [22:0] src22;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [27:0] srcsum;
    wire [27:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h584b6fd3d99027a33e126e15417f55714cfc2a83676ff97fec32b6df2635ee0f757d0dce65d5018cf5cb45760a2b304c1cd1c939b762795fe12953a1a8b25630b16b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h161d93cf570ea613ccfb0e28bec684f4a8a9465385742e1347ec290950fdd6106711fe2876c6677c605e94c15d485c9740245480620e3fdf7f49976a1f71986c76a0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h35f075a47a672fe7e78e53b141388b0092568d89546e05e105d949b4741a577eb38f72cb638276500be51ef548ea43093ec06c9a31bf17c35904e8cfc48abf73f9f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0b93ac43652afed38b7eaa1a8bfd4727de01f6b72e5b1d61b0d2bd5aed2fa234de810c3a4cc01f8c69f2a210d810e8ef60eac8012a5d720bde3023fde5fa9f1740a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1917e5dd7e6c994e8ed9af160ed81a2833e17fb6e90cf7ffe896b4421cf9f6665ed184fc256bf032ef2e5eb27d1426ae186d8af869f42ac743043317c230efe3e419;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a8a58384cdc14065ef5d8aa459295dcf388c0073256be862245d5aaa020ebdf09574089a0221df0180ac56798c002fbf4d894ed6a157ed4b4e2b3149656197d0de64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c96c7edf65453ce8adf460eef50e949b55948677c5a7d14746c266e06f2608395d9b20dfcebdcad1ba07df77bd30acea605b1b7c4bc9b4e306e98296ccf9b6aeae1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha8bc59f6e4cd87def0eb9a734938f220dfdd1e6092c39c7885c0f4d5384697918144c0da3fc072cef1cbf896ec70d9f5ea1828bf10ee45becd619e756d198c52c345;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115212b97b0f85628dce148d23ca95571b499ded6d2a34d889ba7be0a4e238791402fc4ae57dbedae682fa53f0af8287c1ba54b0a6e70ef26e456727981f90d0b05a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17e187189052e0a60753a0e3672f32651b0cf3d045db213632afbfa7afde36e9f67b49baa05ded05cf6bc33966d71a229db698c6dba0f4a8aff1aa3acce7544d87c7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbbfa8d5362f579a9f7f5bb927f925b6d1a4502b89563b22054b1e31ce65ad49f58d5738e88ccc18ca0cd8c13a9af3d2040c055ab7f96ff68629542ebc7e90dfb7df1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h80c32b53500482ea8c1a451d2389eaf605fbe2f94625891b83f2081bdb36c12a3beac114b2f3e360928f0375a230745db512b93e0d5e35bc0d324b3feac19d194322;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2f1d79f35f3c285516687b5ad697ccbcd6d7c9b3fab499e3192d436893f6a1850587fdd19f59fa323bcd464380acfbe46a7881786577164b5d35d6c8493a57777ae4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e97d939d467a8bf6bb2ca0bc81bcff4214380abb5c2de7347ff8172183a4e58ec75a52b53c7622cea7dd9e49aad17ece4d8b20b98b1ffa1899740bb66cf67736a28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc3be48bd6a4a6855fd371baa958f775cb2f3ddf7a32a9ef94a55580d3d2732bb4f5d3dd333b6c6f6f67254e0f095a9264e891ff9c83704b824a90ea91d1d8ff28f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ee30f9a633b91fa6f81de8225950ef5ab2f59db10f8448d144aa3c5b01f1ec32d927a0951d4d1f2832e6db2835116970cc15e09cb751165d2fd9e56ef239c4d62baa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h580eeb64f8aa17ccd8246e05734cf5faa7319568b55b01ebdb7e9f6e15d999955b42784e96ed12e46857083450c75351ebb055bb9ad9ff5ae61639c8a23fbf7af16e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h189e3ba37a33e7b1250aa9149538b1745433de234a0ee95be7ecf096734fc653058971fe789049f7e72b7237a95ea43b995f9a517720d889491e49459c70900d32d85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3d682c3821acbb5ef3cb21c009d3c66917e2e545a244134911717c90b2128653d04f5560dddad4736d43748c240c81952a1dd5da5d7d1f25f19167a0378911708e9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a918415dc1591ca4117424b6c4dea9c68b8a77469f14ddb6ad3d54a7549251cfe434ac8dd43c21cc7b1793bce013679afee75c607cede8334b4d4c7c34c96d49b825;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10374d3a2469d9a3f73eaee6d7d7ab1caf25554dcd57ea6e9a7b977ae4f8bf3348356eab50e1f4351333d042267e957557a20171e25e45ef8769784f3a161e89cd97;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4c0e9779f4f0685e5c2ce3d2b533fa17c993808834d963d7f3895ddf9e271281202f37c2714366a9fe1621a2e4b046f9135cab2060e507c04ae4846fad745e384550;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea766fa9ece721e2373e427d0b3f855bc1c7003c43f7ab8fa8d7ce9956fb4a960ed4a37cec111a900118d9603569caab82d5771cb35cced82083f5c5f9bdd9b8f536;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd92b1946b2de496d52f928cd5657af0e64ad3e86559b1454e6df8fde8f277cb92f20c419a4f62722dc5a7c6fff06f9560b84bbbe6a57cc16cff0ef6921ccabd1bebc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21091352945a9c05a3eb9891340ff46f42ceae95a0c0f5aa94d7c8197ae31b057a9de33d8fd4beadaacb747b6ee87f9c4f61d95710516384919cbc0e5832f71303bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e5a859ef3476dcda8103d6151a30a31c4a495c874c8edc42086384513643fd6b0f39b94bd45ec11ae1807945cf75fcfa4017a50115384d2517f2a04464e8742a00d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2936a8478c5bf211a198e3abd931c3f305f40ebb724760c39083599b119dcb13c32359a34bad6774047303de760855649f5527e4b2a3b56d5e58d594aa2516e01319;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a9958f97c577e9b3d5c67174e7e13fc2b549886d68e7ecd20820d09ac12585d609694cc26339bbc1803913c4aee2db87c18eb6c4d7a93906ab2015fd61beeeee362;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3269d781ca7c45a94ac46341d4622d8239cf3d36fc5903ced08d3e772e19fc97a3c5fd170a1f89ae264ef862b80e504f4072383596d664d56d5521450c0de99fcbf9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a22ac18f39a4655b4c645edaaa868d13bc6985d4262b4a14f47cc570739e3a9016e171a1f53847f13e06bba822322645292956d9533fa3e6d6720965a0a9d9681a41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16b4eb1358bc75a6dcf9296527c9b6fa020d2aaa43270f2c9798861c14fe8db9ccfc3d3465e8e1ce43a6307da8e1e2a3fc82419854b6a302c2f26621c80634cf32494;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6e8d3624615b82e67fa128713cfe915b3f1781b206bb6a75fc8c165694dcdc1f4f00b46fe437c8aeaff1d72363bcdbb5128d6c3ac9dc5cfd5b4bfe96eb283d4d2283;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1323ad69b5d485091c8f98f6174e4bc5e82b92eeed37f6833234f93d13f294d90fe5f5b1a14cca54561af7321eae735a61ca1c26f7a309d05091318dc072f5f93430b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13b6389cedac12aa7b19ac575c90baea5fd0a3b7c76b58e7fe2877f3484f2580594814ace40c74b41ee612b73b534aa4c1763eea2b12ab7fcf8c177ff3a508fccdece;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e9301c2f64f683deac76afa3541a4814fdb83e6f94fa4123eb9618968e5287a9b75c240eebbb4c2d45dd145c09dde63ffb86991ab0a2c42f61f62c90d5c3b6f7da8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1045861f22bff3fdbd3f3616b2d1bfbb9be2a1ce5bce95742b0053a58e4a5098174fae6c8584255571dd3b1dc3e772347063c71e5ec168a0a8fe936a681019b41e1d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h905507eb1dcc729883e193936febe7b612f202c3de33babe3610a55b39a4819d3861aebac3259462bb1e3606c89da4c18c758db3ba962e5b61f5047c3284a55af4b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85fb916612d924b6e893d0a61cb761bef75ddde9bb65a202bc7fd12d21b040c8d59e1dd33c89ce18fd1f27a2f2f241f7efd94d2e1b1c362e556695d51610399aa205;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4adcc716ff249b6c4ddc67a7d6169b1afc87bc34dbdc8fe4f504e1cc8f20cdeccdcbffe8850d4563b610e212ca6a173e8ef5a5944fa4667ca8c2a6fa6e2d1d180f81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b147898dc35fa043a11e7f33a6fc6399279f60c3c44cb635e09ff16252544ae0c49922232173520d10a45a9336bc14e07ed981b9eebddc7b7ec14dd8ce2f0178ba2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2621d8c5d3174f2f347e0558bc3ff549bf19393732c5683125a97d1194567ea3818d65f4bb92d10bea73f160982488ba07cbcb563e65a8a159efa418b7582f7f01a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e2439620d7e1a03b2271832edf734cbe299eddb6b971362f460585284759a4a7a0e61bf231305dcdcf42005bef75868cd25027998ed670cfb398f7020b6b3fd80d1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f405da1ec98cc0faa021e67950afbbc2a4ad7332c2276a9d2c17c7b25f578c2cfa811a2553729cc0584ba84e65c95967be4ba7c4effbad392cc64964d47a520bb69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1876199c857a02c6da694f8cbe9b171a49c6441830d0d0baf6b9d418faf832930e9040f3dbffefbefd8bc0766ee7699074b4c8855f63aa9c580f6a5027818d655b14f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1526c4f08356aa0f373f69a05b13a26d77d9424bf599d1d4179744480c3f560dfc7a3fe9bc1987cb7ec8d5d6ce5b9b92efeaa2530fe70b591180c42c351ab70b5581e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h670a4e945f14269a3a594718960765f557247a5ec247674294e08eebc77162b1d218e0c712a5545e50adf9aec0dcd29219a85470aab4e307c02bf1277110da78233d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1672c7b1efce5a50d31b2d0948cd84843b655baa1fdea39a55df8fcbcb8689e28b6c04fb5bf512a9b59b57b246af0a35ad31734f0c76d5c845e1b8f296e9c7c1b4f10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199b3a687ddc25f6c93f052175430a9fdb029e0ce9f56a82b4e8aa6cf335b41713d99c04a9ecbddbd178b7776251b8b12a6708fa810ef1a304398e37520ba5914548a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10aad9e5e52fcb979e0aed09829a5823e8c78fe7e0730bedb485d2258602600a5dde2d5090ceaeaa45cca1bbee68aa5a57bf616b9fe13e5ff30b712f9f022a267589e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d0429bcd9118542368d1f32fb0c46d16b31f54d067abbe3a69e5ecf77b9523d9ba7f25d7a6d471a2531347ddba8ef939dae15398992f4ecbef864e0bf0ab6b22ef2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea8f2f553e056b7e71372b5c0ddcc23dbdce0769d9d49f15513cd20886a1db46c5dbf677f4cbf5543ddb153bf7e4b90eeee74dcb45bfb3055e89ab4febd02c0758c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1858bbcdef1e52ab0942c25214102805ad41ce4614559742e7242ca96486e6f5100db1cf175f039dea05a850d75acf6a81db3abe7ad1a2ce1c010233b15dc00ccdfec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3fb016453230432ae79e1dbe0b4bddf6593edf0035c57a506132920635103cc7dd9f38e39e683c82fd5be2fb94a3ef6726b78f61d84603963d580fd34ee029a9f22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbdb43bccfa9d16382d3d1e78c65ac052e49174cf4ee933ec20940db08033d8f55c753bc8bd055bd88ccc326a131978818963a7f1d3f809593ed3798a2cc00e02ef0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c2d4a2fb470e96b20fa1d7510d9fbd0fe2e3238195932d56771795cb07c421c9a3f7954f64cf763bf086615f80a906912d3bf826b51ed97ce3642a6ef50d92ff512b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d4ab8cfaaedb9e2c24a25bd89c3117c4aef24304680f7b89b1ef56bbb14d16e674260a984bbb69c36bed00bdb6943edfe12c0a6c9b29597c33ae0f70255534da1f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc282042b94a4ef01104033488bf3024af2d373442d22d995509876376a78012e138856dc0bcb3b3d5ae3b29f884a113c22cf73b91455212c027a28bddc813009dbed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1def72a861e4d0358ead5eace83f1a38445be147deef9878597041bf9d3a8233a44e5164d00d7f4031e8cf5f2f72b5b9b114e5b1bb5e22128ac40a5c1f2396c9f6e8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c38371e981e6519c82122c579de6eb1f7014593cccad71bf6a9463257bce4078e45cbbff440c5cfa27777adf3b8119d340f9363da9837bd8119f81b7c213e340d24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfb57d291b783eb8b724f1f5936eb190dcb8c47a236640589f94a2567cf0a987ff8a9ea1d32c9da6612010766a9518443b939a6c133691fde3591604b1b8c0fe2a9ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d6d1aba058c8fcf39dc07497361e6ddda86caabc5c9fe7f65127a8ec9698a8e82904509738f8f4720c934417b3dc0e71d0f71859942b4f67f2e82e0e3d5ba0ba1eb8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h167eabbce9bbed03e6a05b28d0448dade8bd0d557637e8c501f9e684a0feb4ec35084ca28ad740954195f4f000f747e999851ce085fd4a77235e0660238f6d2e3a5a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6b33d7e0391800a0ab04e92cf75a5723611b9b905d48a04d2f2bb577ca920396758dbf5759007f09a7bef82816ef904f8c15214988dff4bfc663376d15e7058c8ec4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16fea0f6456a97a72bce87c56305d1d70e1604ce5cd5ae2be1be2a845e3d2609e0968e7efaa0d465aa0862756be7f1e07ac76f6f5d530425668b0934f8395f3deb495;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h112cbd111b60be0b80236e1af94bd1d9c8af8c733c400c033ff484d31579e5c518a229a9f8e41767d7e7fd3007bffb55095f8efbf702d001da10f5adcaa5f5a2e9be4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e533d148fe3de857cb5c5ad4dd343b5590cb90f8a150cba69a041ce9e0a0f387144775eab1a281c5e7def390bd1e801d209eee6b3529d20cbae697af2e86c16feb69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3908d606069e6e5eb4d4399dc6e8b594c9c15489099d2c25d84add219262fa9707107d22c0e5550a2ecdc817476509d5f4c188ce166505cca52d8c45f58f4bae2aaa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7376cc9c12987a693fb88c449596962269ec91c85cca2c4f51f520d06d8726c2397ec80065dc3f024e446e990058c0e94b7df23e87641160fb6ad8aa7bff3fe514f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d1c69c3a26d989b92b20105e366a20349e1e584481b555cb0f06a433a530a488f5a56523a57512d4dae343eca7d1ca1525f993400f5e6180ee6c2b46cc48e414c37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151da864bafed01f11c732ba0f3b69112ffdc2e4faa1bccbd577013331c4590fbadbfcaf419d8ca73322ff5de914a856bc3d892b1a6f512e1fa462bf7655ad9b80cb6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef0eef8fbec4bd931bc1e6b39b2536066eb3515d78ee85e36c6c60493bf6d1feae3ec2e2c40728eaf9047c6c799d5240f71f7f666c62ec60e16365d7dc977b0fb093;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58eb356c0fdd2ee5cc0f101d676b4e804e4650bd1b493835c9fd05ec2d087a3698f5eb5d6cfc3d3de67c815fd2f433e9d308ea69715d7a0c8f80c2078022d622d2ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha710e3f821c228bd450b6d79385ad5c772260085be9eded83b1462d1ab7b947646afc8a1b38696bc268e884f6f6e3d7eea304bd7b3311159223b7998e5ec9f5ad97d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h77dd4124d46e9e349061d8d5218d763d0b5a06a77175bbcbdc3241b40916e77b883a6052212c91e56dc2e4061707561ddef5e5ecab597d4af428664a65f2762390f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h188abe40e580deed856d18922dba6663c339587f4fba33fa3ce2165c4196eb55dd8355e3d0f8009c1dd8fc7a44f377f04d5b563730054db34a25041bf56ddbbe448f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e54d7ef10e5709ccab2f8ab1a7c835146c1012d7c3f7d4532087fabcd83719d38b1cdc0e9cfa9235166eb4ec7bbfc2a19400bff4d6d5e5292cdc14500c35cb0ebc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49c93a092dc4ad228d688a31ca0b9220d4df60783c234dae08423a20cf9a77644610d8a17b82f42a7ae5c8489850fefd419e9ddba72dec3f7922d49a3b15bd506e20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he009d632b33ed837496ecfca1b895dbf5ae79795d11f884a0b105b79a597290518c1bc62b9e29122a3dd030d09eff741506942a7f2ac1ca37d59e7700eda4ac3ef84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f419f27743c8fd4c7195632e90a90a5279afcb07b59af71ccd71fc21f223c9258f57c3f7bcdd7ee41eeaa05bdce5d294b1d64a634d01aaed3c84145efa1c45dc193;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c5d4af5016d894b9481a68f3889425fa08bcca3412231d9bcaa98464f1159051c82ae5125deffa73fd87668ffcc3b8a6d83f3842aef21e49ed362ec294007c0598a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14b5e27998a8070516b82555dade69e8dd0c10f5dd83534cb8f1efe8a882efd87185e824abf19f33567f4d7437698c0cd4ae43ad602313436ad120c53a9b0ce9344eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbbd8766bba4504bb98756649e67926e1e45256a96cf21449c7020ba60282d012eceac8c82961e2616659d75e664bb24b1fac0b876bc6ce27a6ee9a88f2d9de58157c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6c95cfbac9657833347af8b6248c476a08c56f2a440247207e906bb80084b930b8ceb2c707f09afbf0c7b381141d2419ff1e5ac58c69406c2ea629db82661dd139a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb99bdb7232b10c5a241d3ba20e1494f0da0b5c6c19f7f9f45439801efd9b998a797ed8691511abcffefcb637772cd6d604a4921e563d851021ad5db8097a64b0c46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h173acc949230725c12feb274e806bdf6e5124fcb8b1ed3999daaf809a6f6596f5815ca25bd7eb5c58a5abdb80331baef12ed655b0d3bf9688be2ece9a9944ff031122;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc46be69ac6ad3f234e5fd46eaa66d8d875fa1e0ccf63fd439a1c36cdf4e99bd8a28d666e37e0ec45553ff43253325f5da4f988d5a522d764685fcf3aa75066e89fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cec9bbea42aec5f17d1690593e8f3dbd4a0e35c65bda8fe1fd94e2d1a3a27da3d4479fb4e0b9a000af621a884e78a95d4e2db70546dd9b8461dcc671e284c57aea0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1910987a99eb03430dd2d424d8c3fa9c0e48e5325daff6b383f063d5f222c0cac7b7938719b21122afb8c35f18b15e96a9d5c3921eaa644cc0e62ba35adc7a2900486;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc68bc12c3212ba2b1c7199c47e92da317e396b0db74cebd2bae5811255e7c418f9e8fdf886b1d785eda1ca198dbf7d2f4e336d940457d560d36f8ed2b728c13630ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h23dbf88b7e0b37cecddcc1b45df8e9771b075dabbebb37232d94c31ecc62ecfd2ca46f19d75f3d9c8a992a687f848f1b4a438fe5ef4ab7e831bce82a90c16a934307;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf02f25c9cfdc8459c3258471ded41301f4a118e78736c6dc2f6bd2d710654c65aa3f897d651e0044014b18e1cd471d322dd451ea57c09a8042f70bc429caca7c85c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16b0132e7202e424839376f4f3557539f77d6c8dd61fc5cd32fe9b8c81d0f3aa7e906c78cba519b91dc31d5adbad1fbd390803009bb41afde616f8ad2027ac825cdc3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cffb27fd09151c1e586ed07a3738b7fc075c46a3360bd8380f67b911968d50e01ca6a44b52f4d9dc658cb17ecf711cd1e8f8c0d07eb6d9688a7cc9748f7876d1100c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb03fcd1a6ef7b938fc8864d6e64ef9b84050b92897fd10be1e47054e7f70247c4f0d17bb24c0a1e27d39fb0d1f1fd4d2a17b9513bcd64e3918b1d65b72aa5571576f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f80a3ff6c9e604aa1444a4c6e67976847080b69353ff46e7d1d484b46327bbd95fa30eed6fc8987b3eda5268c8bfa901d0c7aefb35600dd669b030f48997ffc5026a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51588e1f946264b67d51b904f8929768cc3e85c6f050a3ce474da7523d36f8add44d05bcda2426ea4e7c0edb224cb68788958a7d1e88057dba34f31a293b4c4aada4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c68acc74d486986d80c1b150eb214c54c198cf818b38d23d1eebe51e17c7a0a753da9e5ae3feeff756f3ca54168ab482a5dfeedaefaad161da561977a83c81f0cf14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h34859ed38dc0e6b622e5814bf53a5e25ce778298dd18b96c00a9b94adf4435aa77048a8c6dcf439ed8e4bfefdfd1036c14f3ab4a431938911fb8b8927883a7bf86b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185d723cfb2bb4ced104bd7d71c4eab45ca74ccea8690ef41d085d52eeca4ac548c118e3c572976c729426212fa15c6aff8f69ecd3b7e40ff4a3712bf604cae6f2a71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1165639f33453c37e0f57f903a1d7341836d29d6dcf646261e5276eb6cf0f469cf6551a8671dacb1f9a7831beaff7add4aea8ec39c5c8fdc405862db44f522697e590;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h55c389255b1b268ef19ac1b9764dc0d9d99f3e07e903437b8742313d6167dbd276bdb281345f2c4f84397c2b9c8aeb7a720126a92855961d431975ae5412a2311204;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b5e800e78210e219b66b1a2270ddb37908fedab607a488428e2b460eec7f71574cdba64c02ad7862f547c7830269e00f1376e41b58e86eb1940c3de6f5fd32430bda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eb10b9253bfd03a537dcf5c18001cc55f767e087302e39dea114b1d888524130756cd1b2f1897474009ac8cd6fad3c65e5201ee9b7c22f6ecea4f1509203c3f20285;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ab332c1c6a6e5cd7496d118a5d2a87e65b0ad50485fa20741cde13f813c924c8d454d3ccfc411f9d70441c8656afb038bafd4d9c9ce7b99f14a8f4690e5de3b5b184;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f4b5a99f95bc88a5ea6f1e08f0a67e0ad4071310035867a22c12f9a0463901941559b8c91bd9d957a19856a8fd2a0f075391d9317a6577a6d7f8d138ba07df2e4b22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f9d8b106bfb4e3e09dcf309bf388b566e041b7d543f31decad062fedaace7e9a61e229568cc463190f7bfbc894e2102fbc49ded05aca23a0167358c38930eec52dce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a015b07cd2b69542554a7051c9bffeea6374e156953884648f09f7ec3207eb906b406f643850db3e1ef07add8da659ee784396f5ea9b8ba1af54288b5ec94d31245;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d373a4a4872980f9d7537901b68beb6875ed96113aaf2520c7427b3621479e1e3d3e2544c1cac473b9e0804b6e4fef5552cb93b4600b70d0ee7298fb085055af12b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc3b077d34d6c2f2bf8bab367b7e776806f69bbbf7ae2b625360da970c0a21dbd9de9c4f51a1e4e791ac88bb5122cc9a2cb6b8499c8c35ad96438dfbfc67aa8eeb298;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1057ef16e3ddd5ebca4478b106ee578c5e14433b58230a90d231f8c9b209dce08290181c2d0ad6dca75afe2cd74e14f09cba644d4f6d4ac09cdb723b382075eeab23c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1283d996a9f6fa532218bcc98199cdd3e6c12d3a05537d003a82410e7a8517914e52fd4036b21fe8cb3482532cc9c8c447099511a73e9596e1b35177a11d189ac168d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54b76d626cca20c4ff0adc3bce8bfd4c5f409650f7a2346b30eaa260233992bbb1cdeb32d5a3a64a0c7e870a10093726fab2a8ccea1e713b80f5d36ad490cc39db22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a7425badd88ed5f45f19228ecd0b17a601050ecfb04d864a7b53d1312b0d7e62b4dc26ec4c062b34039c9786371af0bcc68c1f6436ceacc1205d438fa79d0f08f40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7d8ce2b295251e98174fc0ffbc3489f5914fc9e3f065db441b43592b8a91a36d78993e0db78ae5b579eba8548d9e9139db7896737e363d81b2bf3a0f5a090098ca3a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ac61d0c9e08b339a74d61b21c2260c2d35ea9fc18a6548f5f39960caa33bae802663dc0fd91303d998fd6ef3847dc56478c75601dea15fdadcf8a7a35de3cd51dde3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5796c0cf0608317c5f59cfd6205db0ba97c03b957e61cdc89045994b021813218404bacf73a79fff25eb9a23c25b5def90aeec0c4d505370af7c15ce0fb7017beffd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10ccc9f81727cb4e22d738608bc1fde5d623c11da1bf4a23ae9423a8653d2ef3ade508d2ec75267b1b968de506b06729229572c435af882c79f59e35d8874e66dc3d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h320a9990bfc133c7a936a56721653dfecffa369b20538e2587e98347eb3820913d0dcced1282287d6062622f93f92a3bc2108a5bb9e16b04d89c7b794432c77607b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h104c0975705bb2660ca79df114951d9d605a7ccb679a3a7a33b651572765ec1753bac75035e26d6bc2df44108ce85448a2da1cfe485de23255089f25c3681bb65edd1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc49473c313c19f7d86b5778ec9f071b3624beee7b4daa332954c0f38c23156a3aeffb02b31f10d7b519dabeb44bdfda7548a83c7c30f3afa8070a44b28be5c1f0fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95d716575cd813ea2ec8cc74b3ca8fd7633c7a1ecb928b65ca36fafe69353303e8e71f630151a4cb86a5f8a9dbe2f797546b1b51c33e8b601d5de19d9cc71f606cd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7bb1a2ad1ef2c30000cd2e6858b47c0c77f0ab41f53e7ab98721683074a7c55fec7b04cf857ebba46ee4eb4f371b2c98395c6a9603672d451a361518b17108f97420;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h635c5c7cc0b779515386f8e88744e837edfab492e2c7a20ec50eeeb422930c5143bfe9247149ef1a92bfddabb4ba29b5513b0147237105d6c467a4629f96cb8516cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fbfda9d7599e3eed303063b62614ca666f5e7b5cf40df519628aff0adac541290e6916e6bccefb7098e9ee9147a4f1655073d4cc22cd2ab08a9ce693c0765703045c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2422ce3866f2452c7dc3edd248ccadfca1de927b1baca7b8fa0790aaf34e40fcbcc2a4de2d711bb79256dc4fc122ce1bbb21cbb5a8cc0af558502edd3fe375fd9034;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h468a08b6b92e154dbcc8eb0c3f13394e6d0b1c6c2d89fd1e08f801ade29c0734e02987e7c35b338ac0d2e5933f3bf7e2d452e6b2fd9df17187e60a6ad8314d2f2b01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h137bccefc2df1f27fa2afce176a3bfea7bbf911991714f23af9a472bed5e5aba7df2af6f81ff9aea69b5e5689e6aac9e7d93cf21ec4a2e4f4b253bc15a60a221152d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164f3f5167a2de0dcd215cee77241ba0e02f823ad5e14b97c84bad5ebe2662fca980088c9f8a91566fad52bd0a14105624a4e4c33f70a3b137e6fb45cea8ea2857648;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14728d0eea10b3511631c0f64543d37536a97fb32ed0c617195ed17c36b1ee7ea59fe7ddcb6698dda2f4b9bfac7a893f6a2bf71b4facc5d3fd726e2aeb4cfd3615bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a60173d2a8fe31a8d038ad22941b03f81fba5dfee7c876534c6a120be9377ea781d65a42e61470fd833f7dceec2159249a61008be58013d9147ec28bcf447c493694;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb90ffd894edc85e71fc9760703dae0b97cc30c6708fa445c9da5ce4328644bfd01de1510d4513894663cb48fcff56b10943b8981ba36d2c15751e5f31f72677a31c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1d47cdd9bf8d79be0a59eded5aa8fb3ecf68bc4bcc3dc985c52ff6f81ee2af3cd0dc830c10c9853ccca4d4a9a97bd92d05d1b330918268719e20c9f0dd93ce68f11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3582da2abe91f4a033dfbbcbb865f7f84667bec8db8532cab40e7697bb6422cb09b890114344d9e8c875b0f352d3cdf2e24389241e414124eeebf3d06f7f07bc6c4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f71f8a00864eecb50a3dd981a67f37f3c41469190536efd8bf4ede01446cb2012a700931b93327a115d540bf2ada94db98f44d6a0c9f2e87f58e191736873653bd6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11605ec129809aedd01d5b737cd16d54294e9b17deb70c01da8e2e26cda396755a25ef3816b28c1d05d7d862a1b6c0cbd7c83b2c0c7524fc3d42699e2c625c93a3cd7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9dc544a6d208a833d13e32e57f0f05d5c4894ad4b355f6ed13943d2eb825becbf4c6c287b9044686a5dbd1f8da18ef58e5b2ad1e2207e5b5df474769ae8aa34d1c0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1850507496d843420573682a6b0098b0c1b0d8b85c326e4a3908a51a3e101f79ff6cdc96b4c7cfe71a3bc26e8d61f1b9963ac33ff1d65f9d6bd1f57f7f208c5cf8799;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14b0ecb2f08077f8693a5899ea8ab79f795181fbba779b299eb1dd71b01615317f3fea038fb67a6702150cc48fad86a3c73f75e0c89852721f54ffb3da79874661120;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h52d20c03e7c9e1dcc997c070038c514605a2c623080e8ab345725ce1c5339ec8b49ab2dd9dcd2befd489d1baba69bf8d7201c6cc593fe5d7e2ebbc35d0295492327e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb84044968dc0111eed76db69129061a8f925d4a7aae05a735052799d681051104b005d1a5f5232a2a5fcb8cb746b0b1dc4329661478029505696c2bbadc6c37afe2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a5f86be87665ec5787ba7b0e2b4875219c1fe1564372e601df4989b6584d79a310868f72f256037a200443e4bc77450e6f4521892d2402a786ed6f3e95a2e0625e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129c9ca76d7713b03bf1a33beba5242cd172b543092ae3921c843a82dd8b6ff6ed41638df75cf6600146d8f601fb1539a62180c59f495f2af831e2bcd681b141c6e1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he6424b12a79ccdb326bf7d1b680dc9cb9a69578c7f3fca028039aac3ac735c9846c3a709968a9c2f0df852fee4a0a4f858e42e07c3306e942f4ae606b9bacbc00b71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h93e90a92a68c4a4f63b65ac627656be45f0aadb4ffa40ad21b042d49a096caf6478be0de77cd9d812fe05427227814263ba14c2038c283ae1f6650218f800ca31f66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b4dabb840f59f71e6e9992fe5c03ec9d33fb21dc2aade464fbe151bbae2f86a1d8a6db8821472e9386f8d6dc29e16cee62846bf7d5d78c90f25d88b7be57a4974168;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf1a35a7ef5e387ba0f39c01dcf1c3ca52620592094da7091571dac55c34b8e966b4222c0d28496895fea46a09369e5ae526baf9dda59d1e28f132a9e3d75baa97655;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19848a0ab0aad7db3566e54019c3f97df7098b0c7e40e73b40f4004959ea2e8162574dddb3b5e29b24c5a6982c522b646e504ae7351e9181ba76f21bd90052fdaf31a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12649a2c30dac250b22564f7ec5204eda1a43ecf572b18f08f74005065866578c9ff1fb703f55a90bafe5812cc8be1c3e103b41b4579a45df669874097dc5b1c238e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h529a54ba91a1b9fc445b9075a47032928ae1e6745f93f63af69ccf6508fd61b9f5b19634a9c586b10947ba414caea198274d48f86933e41ecf0edd20a648bb5ff405;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h72baf87081aba63e047d6337f5645220a5d10e7461d5005b7c14874c669c3df0682caaa37cfb99f27c910a9ace0cf2510c33fe462481e864a1a90db7fde66709ec12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3460d7e61f1e67f751b39c8e52cae8363681c683af513c596d26b3e5eeb006bed6e3166307d1933404f00469f24e871939bfa9a10cf0ee647211808ad342c7ae2332;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h114b0927855003bac63b616c32210b8982686e6e425a5de33b52bcc83dbbcf909f819d5344dd1fd9be344da01fa1980edd2376eea8411cf948ea9a8d1626459222e5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc7d12bd62f832f45ee209a44eebba1b36fbeee19d4f146db8e0091781e9c16696543265232465c56dc649476795bd2c3af86a017b131051e10f1cb6e9d74915c6805;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a501721c8fa6e2398da97c769b27065597e81e65bd077d200a44ff1958b8aa491c4c2ec4632f270416001e1358a4699cd93517313c69e3a725fd706e464cc2422a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha0f7c1700164d15b378002ad9c7a41e8a037725ceb3cff363778295320f614d174ecd9391876c9bf996e65b882276f8fafd5b91c8491c9371e72ce03e40bc60a5a5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h172036fb8e6d7a738208f7ad557dcf5dad7a14293fc0279e1bb8d5d48588bd74c112e6067920e75718bf47927e43a2289cff245d1b7b07f18d78062bc7527ecc10f68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h52a2fa77d1ecd6ee9d84a91035bedf4ec180bc67cb46721df7907b31f379f411b3cc5a6b8d0d3c60f0cc8cda9dc7dc86e18eaba910511155020d4f88c24d2b7eb389;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc61a393e366a582086791e2d876c75b6c3f50e90e049701420d92eb5167d3dbdaafb2cb214902408e53a26bc5093b00f6e5ed4f3d3b373a6bb5e53422d87b8a2c69a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7fee460d6fae74c6a6b2f9cab8c8dc97995f241fb6c94f2d59736286f98dac4c612aba6a54e8df4b3ab6433c62b2fc0a9640a36ad88d376f66cb3c7ae7cd7dcb2cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a0422f364ced2fdb456632fed74e74e4a695535b69f9ba8b28f262b9a700c7a6324d89b7af1fadddd8b9f37368341f921a0eef3d6a70b425e86b018715d74f40cae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heecd8a509edc9189a641c3aa87f79e3789dc037a850e6aabf8095cd4cca8cea50ebe311a96ab27670dde4c12eb13418eb0260a57e6b4f9611f7f2a37a2c8c5e29b39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he5c2ae9f1476990459effcf48224007ffeffb800a8da5b91ade3ff2778076f86b6860c3de8528ca93be1724b1bace0fee675531e3a0d8ff818a5ddd348b2c2dc71f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10e1c4a0f9b8bdecbc951ed69ed3dd6e712f9f6f29b1fb38b8f004bbc26248f067736b13884ea593540309f1b2e65293aabcfd5f63ccad7b772d18b195523a7c3e13b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155f6fdfe19b7d1698d7147156af33e62b582cb2cb64dac12c91d7e197d1e5f368a09f41b2fb290d3cbba200441d73c8feaa59932419d9daa389fa3522347e86361b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17cf550bf243b201e1fec4babd9b876608e9ad29f13bc1c315ebcf98cc163eaab0c85948613a74647f9a77c424553ad977a064eab12756def09f1fac32ef7a20bdb48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bea7b86f6ea572e283503e52247886e6c0a1675fb177ca929a0027b52e64c5ab77e638fb3e2b36bf7870881b82863264444ea68e04465389820ccb6a85650c03af2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17805a44e99f1d3fd320c311258bb8d5b989674b2d8be20520c2346a4a46728ef1db5cac0890c209a4e4923088e1b6544639e2ff053b101c2554e0a5ade4e51eb834;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19544e57cc138bacb0cb7e92e4cec24be8eb4d3d4b22f8f613bda6760b27b302ef850f804e62d215be812ddce76d97780693bfd476c3c9cd5928c398ab97d94d2933c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cb32f577c0a4da938bb65b3b85d97313fe9867ebf81178ea944de0a3f54c4d5be59a0e08616949ab8d0f1b5c7e6224423bd8995b1938f2b1dae53660175ac32191e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h152ae5eb90cef9a2c4bf32fb862cf29739daeaeb2397df51521379f0267e1ecb666b022dec2b08fa106c25822e15766b6cca91e51d524f4c68d21fd1b4da114eca610;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac5e8cf47628406bbf11aa620a300fc5a50e6d32d961c558abf1078dc27729180d396ca836e7c1050eaf5fad77c9eee723aedeb74a1774283c9944daa6943aff7dbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had5b2edc108b3e4fe38e7d8a125bd502f3dcdda391779354f98f7811f80099facde0029d04551da635a6be6ece171fa452b2bf07b9ba92253e028eea4aaf3c9f1c44;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1be6d8925cc9a7c69e092e70730019ce81451743f4a32f66a6730a9741564af0fc9cda79597e76731d54971bfbaaff2dd5650f28458e61cbf160aae3b8d0e293fce00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1300cf1a6b795ada2935cf4306a64117e42c5f3f8237eae9c0bfb6a4874438b7e78eda39d3604f6a131e19d67980b21367178e79a7d4719a634961b6279591451ce85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15f734769766d9779fa0b2d4dc83d7e67883bd7d346d170f7d9bbf9b58a1ae2a8d9455f834c584c2b358e66fc1b9cc8bfd00d8d627bdf1911380fe98559d176e7e9c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fa8e5e0cde736954c3462472a9a1b0c29eefeaa19b5a83068aeb63d5c3e1c1e3c36ef316ef580fcdbbb50fd2f28637e71b2da31963cb5609532169fcbd88d81254b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb2f0f4c9f281793ec581a032616f32d8eff30a01f0c59702771c94ba13889c1660704bbe6fd1ef94f675fa71ba7b3d1290c2f98db4f177477b4d74d6d2584a2776fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73267bd40687c35aacbcb24ee34a8c41b5553c1b8fd1d2091d7556d7853209aab6b8cf75e532c8e91c16e91577461db07d7bd7ea396bb6195914153df88e8a8c0d80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1db9ec2ff04d4c51e5a18e0664a4fec5c0b7205b8d96c9777b2fd7a4119232aeecb0bc9a41d1f59dd20fee9830d10b8a72375458c4969d16737c0884446560a002272;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18009840c0ff84a1852fd20de1e5167477d52fe2cc6e937fbcb7ee1529fd6b3aa48a569fb1060e760fe6f908e01ac7387a27c59644ea82115c4bcb4f461952515667f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13322ef4df9a51d5f307e936d9697c374674594bbd53da95ad4d71140b0f8c78fe94763f99dfb5ba18ec5cc46dcaeb186df4f903deb30d91cff3b14e8c52784fe8ac5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9d2632b5578ebb4ad44b1aec47f53d72c342192787889b32739204c979fefbdef1450bc2d801fbd0e98cc6e15e679843c17eb61c625413871caf02bf14bbba67bbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a92374c3833882fd95049f37963b95e928da10a09c60e8219ae4b1e7b2bd08c8d61f07c002b67b0a0a96006bfc1a5610eaf69af7d10db44eee2cf75d898806190e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163b623ccf1d05e705a9198f07b0c3e72ef2b61d99167bb4cdbb4f49037a1ef8d3584eb95aee3d9f41e8482ba52b8f4a02a6aa71cfec12c02f98b6471ab08365df969;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15bc4f8c2be3707b6fc24d4330d7d2f54c74ba226912f1fc147933c07321c7c9a037c39c56f9b57fa2f85b47345ab8a4404866be7a8c50c2bd7d43ad937aecd3f5786;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b44b75505ced40c3b628804988976b926d642900d8a49c4708ecfdbe36a86dd0ff5cf4998b926a642c8217ef260fa85e4e5df2e4aa76fe30c7ee0dcee864b013efe4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f23cb0c68e8b6912ab249ffc842400d07e601ed47e160c567f37212b73df8d448eb417b66c1766c22f077eb73306b5c5991f89a10932b56e60ef3c734e6a4b8d89ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a61fed229a748eeec4bc371b85315ee97aaef82f42dc2bc6287a1b3594e6e4498a8b326583728f6beaa8d6a9fd0159fba4372a5f804c886d762c594dbb7ad19347a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12fdbe0d0647e0925161e5b82c17ecd74cfab2a0cb10cf678dd22ccd31bcb8eb8bafc727d78555d5a8ea9725e2a900b7d54b834c5e9b3f170afcac990aefb4a65b04e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1852eca2416a1bdaff1faf564ea8ad453f6eb69e4e6225d6bc6222fc1465696d21ff7380c49dfdfb3e58c3e5f5695299d696e5dc90252dfe1a79500fe1649090195c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h748e2c6effc0fefa6606956eae4a143e3ff05a58134f408f96171648447f5446bb84d70a1eda951ea5c47b41de3ba656c17cbc05ca1eee3254c5b6343803e425323a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19ec09c74b7ea74330979b5c719d6fa26b626e71be32edf18cc28674ac88170e3eee75621373549592af031962df3087f0968c144035c40cc611ee76a14c3aabcd558;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dda2e2ab4128efc59b1ee25f909a1e1b0958b5eae9f2ffd8ce2bff02734cbfa960b8b4dc820f717152f52537de886342f04d854cde73b113e03ce9635b8125bbb00e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f6c61eb34d41e988754890ee2fd0ce5431081f5c155cfdcd0753f10a77349d98e41bd9b3d174878c451fd43055ca68a4ccb9ccc54f2b2cdd10f83198b9a4e3a034c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e7e474bf9fcc0230c610907eca677a09ac1a58e711f5ae8f816a5d9ba4013dcdbd5619a8980039dbef2aa4e20c701373fc557256f458c9f856d190a024d3df1bc7b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198aa189b90677ab6bd04a31fedb3ed9e45ad5138366fb5b0f1bfefc0503419794ded602833a018160e0e76a9f86711847ff564f24d260aec6f38cf372ffd7132c60f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d4331651a579a4e7da3731e166f6196f18e877dad67883668ae1e7cf354366298a38b570f07d92a480cba0c9f898ad99385b68fcc767c2189990a4d5f91cd8c84f9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h125a6bb12416a7cde506bf60480d7fa4975ae75098619a824e1d5790de3a40061b2515717881c031e9212b17c9bf9fad211e631f99ba2c0432e5954f39bd9fc867397;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f40b0dde5afdeb8c779f9d657485d4a541d5c8249e76c0d5dd8087e9a0b5590782e48b16344d5f1ca69f49daa6b54d528c994c99b109c7f27bdf6a1a1010b9c05f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf5cae1cb9f827f55b3dada980ba27bb713bfac003f5877dc48872b6bdbeea58594b24c6041a6ab051b71da511460e62f16d00c1eb9b8c4a495fca419b8aaefbbb12b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ad063826856a5f578fa7173a266e11061e4b58c2dd058cb59e9f281a2e30f3e6dd875c0a5035a7340ff30ad0f1e606cb85b899a1f75abf4323853ab262c3d66f1ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'had843b334d2d474119390755f839e19eeb8da11b0d51acbaa6d0a0af695d501360fcf7fba1b05bbed4f2f6890997238e476cba92c0fb51ac0877c9af5fbb41db1fb5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2283daeebfd752d091795774726a84bf56253636026d1208fda4ef7c8b55ad93a5bef1c73a2a2697c6f53c845412928a0f4913fb8be2fde5f75380ed0561fae737c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19d7f86ff40939d898fe03ea798a149e4702f2f9da89fb28cbac484a597402998a99f0744edf77e795f44b063481a8624e4038ac101e2d07270c025561a47ac4d89d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138e89cb61ee8ab629f2ce282add9a6fb1282e594b97310a9aa87fa21b59112b36716e7d3379b8680cf6f1eef4a6bd04b3adc3e91f51bbdfd554b24b41db0565925de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he4bda1ce6829b70fc0e19444d9a958862be4f52f77f68a0c5743f22aeb13a7ef81979b7b200f3e706bc1a72ba1b5b5113e13b4f57c73c091febd4d24e99f9d3e30e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bf0fd6019b5f00596c0b3bf67533369b2a3fd4b20044820155271dc691bbf1b285000cedddf8dc1a1b945745919a95c9a92b1d38bc4d9f673a1842a8c944a8a20186;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a7e89b77e1173d8ca6d45aefda962376111f242b723177d1b403bd152c2f01fea6ef2f364f63ce4d37df8f8b90bc5dcd97a68c0915f6c71b2166a8d4446c27b21854;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b96bddca3d5bf3779c1b6335dd22155a4ffdc767052a6dc4aec2965eebf9eda42dc939fa1ebcbdf81f2eca6af60eab3abbafbae8af76fe390d38118a414d6b13cd4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha7f47b25aace8be0bbfbc70ec6ee41b21cce0e0dd232728e5ef7e9c18bc94abdb0273676f3c1308d93eff9bbde021f02197f61cf992515f831f2cac863bde3710cf4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12522d8a1c6ee4696f70cf2bc04a179ba61c6f1ad5c70f87a4ec38b05034a3980b8ce6c9a6a66738e322f9dc059ad2515a673150b013f9a03e382f070da8fb2dacf4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h73f66d55d6b73fb6b2078ae9a608e336ba22cb4ba1ee2244ea7e1fa1d675f0e8884bfa757fe5a8d089cee97a37a739605f430f5762255b48dcf8704041e4d8722646;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he58119b59315ef372a0195cfc484b02ae2cff2ef24f18440edb134aed1cf4ab6b19914d2bf805a5c129f2bcf283d68cc7c04275666b32b1f9ee02125ab3f1776e2ea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ac1ef223eefe5560aff3194272dc2ff1c4bef748dd5b7650c2e048aaec7b9e2055a7bb8e47b5c36cf62b3e9de4ff66e55b181d8186a61253d7d6f187f51adfa7480;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f87496859f0738bc6e4a919b52b7219be6017ca703b35c7f46981738c3ddacfa2958225281e1ce7009172e7983e39f129f9b557e208e55787cc559cdbf51a940bb8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16b8341b6971809596706975a07ac1b3993c846b2cd78c2fe6108d3e4ecfb8290c267f13fb248cb844135add21dbe47b33143cddfd1d11c422230eb5f5a6944290cee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17b83d2a9dcacaf95ef34ce6512d4769643925dc53ebb359672690a80126a917bc34bc1b22cbde780f108166544f026d34edf1406aaa2d6b9becc68fa852248e53da1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc44fac21f4e2a54fdd7265b7d71dcd7259758064691493c7f9a1192ec8434706f9654e98c499b1f83b443122fba24615fa5069b17e3ad996294314193063367049da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5b60cbb6133d8703ab33348965787b8015f2475c9cf51e3344d5e60abd1dc6a66fc15c4c8e78a2d43bb30fb6d019f85de2d9265db7c8c696b3f5955543f38f0be46d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1893f61f47ab908addccfc8427663c8e4b34bde134f4bde5a777f64a776596057a13e2e0fc3d4bbaafb3ab8375ef97e4246c5e48de48d1d062fe7cc1ba3f35745347;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1435a12eaeff03b87f6ba566255e47ee607420720a444791132fd8de9b7d57306050904fcc9f200a15fbc142cda9da0c9df133a04d1f0fac781774b95717f12b7a35c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd934d548699fb4a60ef13a68fab2057a29758b771bbd450b1b810007190f40e68d63e43e1ba9b0784c21099c9cbda684846c8b22e8790e369aba9234c13388a29ab3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17e729faed6cbcc2cfda6adf6933f2d593069ef23ba1c699ba8200bb078a12f6e0901cf35b0c6ebdbf78c601c965d067005c91adc336698257fe22c5ae090ae25f4cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10afd4e246e862e1581683493eb75a6fe37af94b35b8d3e0f7c22318e7e02ce3d1a712aac3c8f5c525c8e9d5fba5bdb0f2e1fd3d87e2a1106eb0d60b7cf4a9a87fd1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h42a57c3adf30c2f7b664a340a6646802dbf59c040f91f288d46913debcb2600dd5667c75192fae0cd397e1cc90bcd1b6d042acb531f741b819003c6fcd2b3476f388;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ee0e2cdc2de6a267125a93c7d48d8ad6c603ebf55068b6f4778db1a601a24fa1653f770460a4eb0ad8456f0f89c594caeb885da5950f3d54a04f47d59b5f3fe6009;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h129fb7085e35a955b3295c94b793b4ebdcbeec55bf7a496452af626b54fef7ef47c0e0a9edf36155cef6d6fd3b5a8cf102f7ee79bb3703cca375b597f4497360b9dee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h23e9adeecba16c4701cfe7245edb4e103cdcb1a6863e154571a663212960019d599b9788c8b3a8954adbd92ba4c0df36d366c147bda88da60a6a13ba318c1202bc1d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h785cf9c3e5e1b5725d37e1f9e5c7b01419653cce15a3878ba1da4e0765e807a6ea1c8afb7bd6c23777b738a0ce0f97ac454f65fe883522b2251c678a561546d2d19a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf77610ae6f53b6a72e54c607cb80e7d0b97b250266c7db717eb537e27851895544d87487e8a332bc421d56564dfd8979fd41d7c0abd2b472f1024adbf214c21371a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ed3bc2476b8438ba0fdef9ec7399ce92e99c28e340286327fc4333bc3d64759b3cd53f466b257efe229714c0727a4bbb62526cab1cefd54867834afdb63ee0b9f46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2da324e1ff66230d137c8beb8f5a9b62b2d4135114d93fd1d599c9bca1fb74817924205097d7916602ef19216d576a8a2fd1e6a36f021cf48537efc45260023e2ff0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f50807576413f69f8b71dc787d6a883e8dfddf251539f37130d720b8e5df8445f508c16b693b8635ce9ac3b1bfcd6dd37f9c73e3eba0975427e4109cc1bf9da7360;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h618275e0edebd13ff0e99aa913a79574c35f0fd11abbb03946294045aa6d7d29e478b9411d5c1d700944e8404cae445fb5bd094cf18e856672ef87a76162a10b3744;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h421d643b9e1b6f1a6cc52455e29b282daa6851ce18616fe7612208bcef3511e6ff0701b4eaaf9dc10a6ef228e947376cbee4d91e9c33ae795c8434ab6d165f3d6b02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h190504c7a2d32b832cb0ac7726a6da1cae55b923d706748df0f88c1f357b211b0e0229924408d84598ef104569b3fd94f9ed7b261103b2bd6b70d72c30beadf7594e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h867928f5aca3557db609d09c048f5bf362d3c79a8772e41bcff99aca7750ebb915f53b4722389f2481eb6c2837a0f3c0fc0100d027579cd3a71d894715b4e18f6bbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h378a55f943ae93d7afd4ccfec18fe69c6db8346d807388040df8232ce65180687a4473d8002edae7c924301cd6d0ed00956e122bd5216bb688c3976b413c19b5f9b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0543663b64d2616c3574e1c2662039289fb66c789948da49489084c369fa299619a9e28e5afeb54d48a317a18091cdc34f43c320db57055f7a93a3f2ae86e0ce792;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f38f970a02e5898b8c36d2694a5ab97fa27f81c1d84ba9421a3475b607a4784e8b9f41bdef9c0e28bd7eb6bad9e549ab355e76de2da1722aa27d3130f4db79a18e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab03358c07604bafae3cae6e3b817e2ca4e2000e9cee735a4d448c2ae7ecc9b4df29043e9da197f213d6e64749f1801e1ae30e638c7b6e5a8d4e5084e2c71deee3df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193455246ba9e6354711614101841c9c7211135967c2678c15893b4c7c9f713527716e7f73d50102fc21e65beb1b24af454b1888d551d0afbcebf610e6a8ce929b3e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h542eb8e44f30f37f0db5c1e84b0e9fa2237e9d93775f80334d5b7931fe46137bdf7e241fe1043b80cb6e3fb60967a34e080a8e077179b4a71f58897f35d1cece7ca6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13c91d705df28f1ed164fbdf8ec259bcc45c5d6f406e415b33b1430d35d515a4c9889acbc29a166c0692206784fcd090426089d0ae5b67209e8148a8fb60ac1aa9da5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133001ed43ba820ea0c1b732c891f339836cd0fec2d60c41c4fd9627f8b2bd6371e23c3f94efca9043c0101780e666ef9c2fdaa6ed9f02163439a57b6da4828aecb69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f45588584da366209a75f8dddb8db99d1c78d0509e3619aec6c2ac92fabdea3b2871b0ef6fdd7ff2e11dbb1acec79ff03da1764ecc548c1f167ff6de84d7052e85f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d297110ff7cf196170fddfc18a220483f60071b8066601b4c705d2c25cf890bc6ad3b2622cffd47af7b838ec8785701a710a92a3cca8bba245437ec8881bdcd52c57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hde58759c73f3585f745a121f64fa5c94eafafd1243c4b79ecec0525e192842392b807f0d1a6c4b3f56d299ad194062f94721528ca9594079e4245398159413c6e1b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e1d3a42c09bbf919b45b3c1df5b90efc0f872e0492afc27dbec987062892bd9ab543cb4995daa875220413792d6bd6dffbe90b4ad6c8dcdc7f58a4b7cd42a35f6f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h961cf8c0aacee887534a8f750a6aa55395e67485975b3650e5563cf440cf315967c828e321dee196f625328cbebbb829b2852c90e12e45f92b9dc88eb3b77b47ea9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a12cf74a11667ceab416bddf25e073c036aeb1e52638bfa6ff7b17ff7c5fd31858e74d984564d80584e9d2314f128fef1be11b050d0b04eed37e13cea2ebf1fa979;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0241f901d7b824b24f08def463892b90d025d43dd2adc08c1c8bc9948824818cebb8688bc0ca052dfaa8ebbcb1b4ad662c39b7d85c36f39ca5f93a9e7da4fa4ecc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h112d410d038c515f56fedfeffa122efebd69e9a731e8feaa2b866adab7fd38e8eaef7703b5932f89a7b6024adbd6cfd2570631001b650a9aa5805f27e2405792c04ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10abac86616b06ac36d82069e79c91b2b8b09ae2a2b6603f287a4e289057b169ca046402d77d39ec797d887c8e14544bf6514dfc005c3365270e4ab9b66492f2029b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdbaf866d0ad7e217d39d81b127d13cd15150b4cbd6794aa4d48bc0f68a9d7482aaae0563a4e21cba7f2f7b565364285392cbc9e07d4832c744ccdcf6122448b7cb4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h77c34d35b783b4097d7da2dcc54c54a246ce795028d8bbec00aaaa3a8162e091ff1d039f600ddd1e099d3a6c8083837fbe680d1e77c5b9f9ba9bd02e620f2c54aca6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1264964e65ecb3284bb7f0f6bd72defd90e62f40354f1161e73c3c668e975340135991fde15e6c7a34364f9f65eb2f710ee627abb08c2ee7c3ee05d1371ddafcee36e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc741231845014bda1e20326942b9252a31e4c326ea9b30058c64465d09dd3b4b95edf02fbd8e634442a9648367f63d25e156344a8b11238bbd9504be0c2026d8996d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c924229b3ef4a95a68fc5889ce59cc112968ddeb06576317acea9c137b6faf39b983fd68ca7d084ac53fd85509ecabf61ef64b3dff5408f0b446cf9948f550b20cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6e62518770bd2e5c1a123665d8de2416d736f516dc5331370aaa50d6a0fec6ca95cb6a7fd44a98b7c4bd7eb3515c7ede12fdbebf3fd24e0e0aed216bd51d1ae94a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ec602b62611dc3b2c757263bdc05f8f4ac7bc629ebb8b56d47bd47affd55f3171099bded75806b4bc74c53be6002b8011a92890ed6d35b28b02d1e77c51ef9cfa97e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h118521c8b6b056072ec614f0b2ac72898dbfdcc67630d95461b9ee15f2b50b440b9862140573aeb556179117183be75bbf54987f73a6001195762f434b7a8b2d501f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf00825188915b7437e18eec9298a6efa8f110e39e012363f1a4b4fc68822fb18fda1f0e4f63b1e31a2a5625c5e320e19e51b41a11d9cce36cb0aea4b80bee1d84613;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h276d014a62cc052b8047544a95b81b4d23676bf15e868172a1de7dd6aefc14e8495ed506bf923b68588ad2f42bb3922e350c066c67b7732b8bb09169e4401b0773f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd01aca6c4e7f80073549e206119339c1646af360d52ae919b3301ca86f2e236697fe78aaf986b14e895d9660aa9fab11f97f8e799a66428ebdeac50cee1840f74d75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cab69d04c6c24618a2883f1377750f78832a81cbf5ac4336380ee4f086a12af5ff95543c0286fda2f626a5f9bcc3a2cb3d686191966aeb9dfb8091fd129e544565d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9dc9af2b8131474fa5b79a2a94bf3cca475a2d6035facbbc671c2bcaa651ddfcfdbe8596a168adce53b1bbf06c549bf26305bf16fef9641f562d61a9747a15a53bab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4ba680ac269aab0724e0ee3a42a1acc3aa977fbc686101536c5da344cfdce2a6dc7c14bc39c4f1285759a5d379a6bea81d8106ea5bac4e3cf59d464d1dcc279027ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19c679a6711e59020847e38e78290e7a3dce7a9ca9ae53ec6cfeeb11e25902bb7ddaf9521f7da0357d3f60e3b2d6077dbbb2989729ef8d1fbe8bb371b54974da49b5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h203cefdad2a23c38b14eb1acccb268bba00ae9759d5ff4bc8f9c0e7c0242f12c56315abb465101c214f53a754fbb519e14759143eaf0d090a1a40d261724d0922320;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a857ef7eda74149fa5256c6fd1e1d130c5872385b487f438ed52cc95abf405b05f46b75795f36f4aac26cf02f9ac4f2579b8603b096d1b58b5732641356bfbb6af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb32a4a81997518cc877f2c85544cbb3e851b82deeee23b760807fe1bfae0bfe86291d0bb520ea71cb9fd7ea7f7a0b72f7fde25b7507982d47ad7cc4b35d0d9488e8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf84c84488a944873357a7b2edd3221bb8f79309d6d4cb49ab90611f51d33284c9f37b7e63b78fde4fd6fbdb572bedbadd8c1a89a3fb1a48b1d6429a0f96ec3ae0c75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h23f3d4d06c4759b002fbb22fafc6945ceb8a17366ce1a3badf533ab334b8c7669da3b4ba48a0d2ab06c759fff5313515e1e39bc1e7a7b5bf245f23c6e10f22399996;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6ac91823bce2d1b0f4f9323de7d9c4905b49e61af320bdc34df11ac4ec31bb7a34fa400d17f0336c63ffb3632da9effe60acabc7d7e40a443eb7e28fc76f8680e4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h252ce63c1c1913562f88b8d614a50ca64238a022b28a749e5b76f46448d4ce7c74aa0fedbf8946b6d98a59c24897a22140b62509c576bd9e156dba6b990748147913;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aa99dfc28bd327ec022e68631113e250ef1c5fa202fcb0a1bb379084357a2354c49a10f4f06d09834b4dc9106ab8c4ca3e939d8659508021da1aa004e463fd20a481;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h98a5ef22ef0f83f0d8b0d3d01b7464f7bab4bc050f2998f7668d3744e222bcbee5fa8b3360bad58f2b4020e8994b624aa9629a92806266365fa74bea068a55f99a7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f1be49fb790c10d2514cc3e3ee914ff0d1d6fce269852276adee53b2711588ea4044cc9c3899ec7f1f78db5b633ce621ee3cd3959b575ca1f8d72d51b66d0f8df168;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12bb218296497f33e753951cd6ef91bd106f2a8731106a2ad4bde8ef7789b8421197ccedd1c20753c24b15f6dc3704b21dc668670a1b3c5dadaf91d5b50bc5e626e78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf46d24c9e51c6e508d2505609ef8d4d6ca7c4ee1a73ff98a1539de0d132cabf6a20a6b53de5cbf59645bfd9abf8935f01b3fc360cc9ad963bc235d28c8ed31478ef0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha55379cc78d9a3d942fdee5ceac08125e359e77382c6342cf264a26740ef454726d9cd532792100135d976f2002598b389e011c1933414b366595e27482cf994b8f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11918efaf7608a7c7d00abe52de1178904ae414433ca380edcf6aae1530745f5a4855eb196323346116feea70cac3a52691c225f7668eff17b4c681bb097941896501;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h199cacf374fc9b5ca4afb427ccb391a05df98e8004ece3539a79b5206742cb3854e91ae75240f13ca6d379f6de399a4e1b35887db0088872bcdf8eb2520107470bdd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11506ea59864b5a958dac56d76229af04977efb8389909978976a1d146547484c5c86763b106bf850438cd41f7454fac6f6e63fd8bd8ee2927c5eff8d12ff60d5357d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3220b0901a94b2b454046a8f999057563029e30d78260ac3a2f6180e1bfaa156205363d4723b9b8b82f5d895566137785aae747ade00468d858c1924043deddbc31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18aa9a16ee8bfd157239e0e612ec27197236fd4ba9e6066aee74dcadd89ca871abab6c2a4e545e91e371647206dc1c5ed3e9b1c912b0487adaf5efd29ef82d228eaa0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h50560e72b0f1c19b3ef569707af5c2b282e77278062d4db5a5898ff271e8ab511bffbc09fda80cd4cb580e06711e288f2d237f02aaf35c3c3a7c24b30499e433a9ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128d7e4c78935b26c5686565b762f6734656a72d84308565c7120022d5f79b17abf5a2b1346820c280b13d67c6ecef2228bcaf9ae4eee2989bce81f138f501fc65c85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h155ceee090317fd1cf9837983a8bb85e7442fa6e4a3c088a8a0faa2dae8e6a1a552135a023cf720f4634da1f473f8f6ec2f228b7917637ba156ff5174c104907b3cdf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hed3f1b676a396aee3ee0ba970f729d43491298682da208e7c44cee04dd17a0270b9d1a00b9faddf9dd5d8d844005c21cae32107c8b740cf66abd2e5cc1a730fac21a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166515debe8621ba90a523204fe2a45fe2b44c5b9c20d42346f9c558115b4e2824efbf3ef420ef1119dd3df9c5cb4e757550b119fa56df10a5b4a28a59f0a220e21ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h139dacd6f7e75c4ba8831f6a44a69fae196533f92b9242832cde7cf8734441f3021e536bf49fd67a6a74a2446589b7ccb2bbe961793c9ad8eb6a3e9c24c75d072c629;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19575705b51d36ce79f0bb0551dc916501f94de5eddb77186c6fa86f9c1bd3f54bc2aa13c5bafcf93fd2aaafd6899238c86f95ca4bec29eb4342aeae4c286e010cbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d2817ed8de1a34a7e19180a5b3e8a006c8c5838eb306a92a323efc4156d38f7d6985d66833a47b20e0089f9f3411984e129508d7ee8c8b8941ed71b0c52309dab6e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1061a45c169b809f17c5c2a8d53aaa675d9f3342e445bf6b99dac6747a1d1d924f4997897126096bea445b5dd62788b8cc32e0156ba7e3f35863370705cfcc63d8a75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a3983bb3cf6d284ca707996c94f553861ba50430c2df34d0dc1ff8da85c7b0ae3727b3627959b3baf8e44d88f78bf88d6c17da8b85e5a05f596eaabbd74d1a98859;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182bfffb5fd83432084f6bfcbbb1d9a1f0fd56ed40b5a682639d81cf02bcf772724e31020fe3476dad856b27cd113abf58b0ce311a321b4b38744883cc8304e4757e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1505028c787d0b5373cd3e4c3faba0fa1f05e8b1bc2bda798024954ebcfaafa9b2ee561b53762c93771b835422ae33c4db80de183ea09aca62854e39d197acb5ee9e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cbd5048bce07032b057b562b0a07ce17fe9ef55868aefa05d84a12c0179e403ae1506c8d30f5fa84509f15fbfdf48f16e274c1a9dfbe66313f2a354ceab724721338;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha0f48af4d69491b748cd76cca7b1f21ccd439535dfd4868b14865790ed2890dd3278fb59be1f3d9f6b3fe041718d1b0e28aa5e4a6d43b0da1a3e4655c10039f26616;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf98e3a6929e38e46dd5808174570c3a69d52b772eb0d52535bc918a9712bbabae2aa1f9be57ec4c800aacfda5012c3878dadce86a5e8c8c115a8bed248303e36cff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2470f0df7eb875b5f8ab59ca00facd10f661fbf1c1d4cb25ecee754a824c69ad30ca8b01c0a9b305f0f5fa01312437121e372ddc4e41b6c833dc3d06e3169416fc49;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15e851ebbc2b0370a983521a250e1a8cc584771426ed81b756a262407cc4651be413f1417cd3e9bb2b47a97e0cd44bbd7e0ffe8c5fb6c2413ee5d7227799ebd014c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hac329c9940f456def9c1bda624e2c0f59945d8ef0c6132d58c21b639e9c29cb00e5c17c909c5c62f1b34fbc24bc5b5bb2fd354f2b083cfd2851162363b2454458a7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h88a66cf348c2065c18d29d2e462cc2fe703d11fd00862c47651b1303f65f631a4d7b768ad16257687247586064ef4b04ad5f0454fbbe4f59e4dd6d8ad7bee9a11027;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1798f3e29a5556b62eaa85b3865c92d8df45bde838a2abb01068e99c80cbc015d3eb813db1be6702618908292b1a972a879a39e25875a8bde9196687ccaec8144b1a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he0f4956c34fa20dac005ab83e13b736b4c6cff41a2801da22e0a8d1f55dd1c74fc12e85bc25678849491b17056a75a4dcd8dd251ce04b56d5994497900159bc45e8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c2a60bd420a7bf726e1b988bded1a3460cd1ca6ec52f0c1450e860d1380ebf92691f5c7b3da12f523f29b45bb9e1cca0491bd9977cfea82cd9a5f1d764d83678756;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83d99a1402a6b07046e0a1bf3fcf3d54dd54353bed62bac105e7b41880d9c4600a411a7f704da8d76e54bf2e4c323fb6bd0b7cf60a81d6c2726a5758147b463d272c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5296ab99e35e8f829944cc14a2e8b8b8850202d572467d93617c48520c1b176b3d5997a80c96df654934d7738ba16e786f933a3ceee155b8609addcb8bddb6760168;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7b196b1a2a933832429595c7c4d7ebae01ecde4e0ae3c5b459531757016eeaaebe44bb9218fefa3a2e3e7377b0fa9cb33353bd78b1003d8ccdaa0584f097d3c756c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16f557d948effbe7633a87c245410031f6af1b7c96bbcdeef80d7de89078ceeb048031cfd08b54e2f7b0fd6422e73430d52b8e50ac1ec6afb282da244d4d9e8a0961;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11fbe04a87e1fb02dc2fda5aacdc13a80571e95006363d226e4eb82228e686b0b2b9a5d7c5ef117d1539cdc510c0bb2a60a216d610dbed1bdc871bd44d4d30a855153;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6667072be34061185aa04055f314d89427eed71b51a5d5c850bce019006c6bb71b5c9ce326b00751eacd225eb79135b3dc298f9c03e7aaab3db0a59112538e87ad7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66a7d97cdcecdba3566ad5b6bdf5b80822146500a639e89dd99787a39bea2b049b2aae528f364542caa33895ec69aa2c111070b6623e47f64b1e1b137eb63a40ab75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb35f734e7465818fc241397dff2cf718a0796ce9fd6a3f474823805527f97941570b532e56541749706e1c986465a6d6a1b23f1df5e2f3497f9750272c83f1741cbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16bf158fef3997cf52a58992dc6525e32946a23cfe77db7666b66694e41a78945f2f263dd355ac69b9e7483b952bd275ed2015c28728365ee800bb448106595eee89e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15eef37e12341e026f979a58d76099cac46352899835757ffc67f9f375b42557521c6d4357266fca8fd14eb19803e9190d20ff749cf252aa883a96301b73998269c90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef76488b8b30d9b7eaff1f5b6df8b8abe2eed8de59c9922f8d827a26bed2461ecddb3b0bd808c8f358f269fe8cb8babaf15f0efb414b3bb8defc0a9c5b41f730b5a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a98a6c6c68aa02003b16b75a8c8892eba53b7ba274de56f3bb4c192268ca9a5387cbf8915224234418cd0fdc1fa32d5df905275f3b03c6557079f510df320aa844c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4586f0d4c3a4ac07507922d073a2849dc8e118764b1884b34b9feb14b52e164d10fc3d721c921b42f8ab0c6354842c85274117e96f7747d5d1349437352654229c22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1074b12e7907e8a6edaa6ea87178b6a937aa5722a2706272db0317cba4a4a8421c3d2fbcee428706e3bddc87c531a7c53419d3bd68634f939db0ba5e1400e7853d608;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16203cd27eb645938689820e83d0500da6cf707b9b4bd320cc0f37ecc5223aca35de98b1e6af25fcd76843d9a097b46e663e9249a48fbed18e09177dee8b4c083f8b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h159755fe6a7ca50a635523d6e0aa7e9a6af7ca25f0717b964623787009015332762764d5842c66ff227fdbdba8983806bf4e9f900751040432d77859f5509f71a71fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h721e23b5097c51a91a82f875ff1219675fed55baf5d342317a3b8db72a7392e770c803a101b4a7abf2f9dc5ce0b519001ee08d421822d7a0c05394ac48020529209;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8bd83fa70247a4ca52900be7aa8ae21abe10cb61cc2798fa25b1eeb033190ee5869002a11c163d20ca6e3cf9507dd8239a380d6309acb7eafb7126784ab3873dd441;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1017c7cbdb8ee9ab07d38fca543f1262ba1be6abf50e2f3235bc6a423cb59d98782f24a3413101eca47474e276e1b7a0e9ffda84dfa24692a34de1a620277493bbedb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e2b5e394214f1309d00f3a9985f99baccd6461b6e3af43b1593aa0ac483d4c87d9b7a9ff121ea9bc1573459744939035450cd68138ecc7431acbdc6f20e095de317;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12f1607ceb29afee06f9132f0f8a1ae19c44898c54704d84800438cabb46e7a3005e8c023b22fb4131689693ff3d117618230dea097fe67e90a1a43ae4bfd2c38ff88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb4747a61c601ac7a48804670177a371334120d50669c1b6664ab9dd96463608bbe6898df987df0e581c55e70fef62037c5ac49251de8dfaa14fc891992c0f89ef4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dfd131b0c92d0db6eccb3c904e7ef05ea3d39f82203720c3dab7a5af6cdc097c4e4fc07e93c8de089645986f47f5fb87d63d33f3ccc0a117cf2976253070f12e69e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h47d6efaafb34321fc1e39428c46efb7d10c08b352cb9f18161e3c146cc8add3b795f02406847d7f7435cebbe5359debe8bd658349aab3bcb6c6477b4bd8b9ca80627;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d5096e842cbbcc14b8c3921c2085e3beea27546e0798a6998fda57f5336d63e4d9327c4e8d3c48ef714868081bd3926ceb2e44af9d27ddc1a326557764eabb1658f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6db7702a422a1ed29f3e3aa076a79b48313167960b002f77396b7377c126f4858eec846aec8fed28f1336b514cc38de809843dcf05c0c06e357ffd5eb0418ce8698;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hade72a7e7e7c9872cf9b1e33b78a98164dfb60370d598f0a64a4ec3452d84c0abc8442a538eb5e7ee9e6545df5b54c2990d40964383b5433bf698d64ff3dda6375b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9af46f4fd345679ddec5c8dc510c86be4585e31aaae924e8a2ca77a47bdb50e4dcc9d4e0ce3875822b170cf0216968f58716da55b226d06b48bd60446d30b0fe8637;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h364aaaa028a7cc1b1bc123262b27c0b2cf7d5f2d7cb208d7bf84b35afcc202adf66005e21d4c2806007eb2d5b8851ba1f7175c4d526cef5350c7eca136bdb772ee97;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcec5124b4331dc39d033777d3f3b2cd5e97c54c60c97c1ef0394be264a54f53d36a252ec19323651f4ea38bcd02b24e38f6dd26038ba095152026934cbfb00858e06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12adb4587c9e7a1f3b67db637569401213bc00e07975eb5639a48ff4216575be248266ddf1d12f4a2f96336c0f05237d7d35ca82ddc633654c13276caa0c6243c5ecc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h39820735ec4d6d9cc9e42039a1a78971fd9a8d428b4bd372b7bc743e458871194813e3c9976b2c9e06f8d8d5fbf8896fb62439fcdcc326e680a6ccddb9c2db10944e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h388ec4d29d61a02cfbaad86bf27f6795d5ac6fdcfa2e98cfb148d513f39bc724121057d5920c9157eb4dc8619a892f07315059b7c16ef9db83c4958904c68c5d594b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hea0b12a45fe7a9bdaea29d3b7bf6f7e918f71774c837494d9f39f03cce37a05c3f5f804f17ea1e7dc3ce42306936728d5aeb02b47f2a197809a497364cdff16923d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h145d1b25c1aeeac0ff95a86ad417ac4a4889a4db4e7b72cb589fede679b42e76fd5ea572a00155957ff5bfe71668618334f6413776c5d1e34154feae2380c8be22084;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1818e576690d0c7019e13eb26d8928b968e52ff4a1435a90de346220458e1d017ba299e5c2e38cdc3647ca00dc6cb99edc77036c6f61d860cd66c5fb0915c2023ee1d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10abe0b59c4ae7084a5050bfcdcf2ced33239e93f4eb6b20badde1e959dbf4b360cfb340b665993bac1369839707e1b34b9fec0eec15ce7946c53f67be16b0b9bc695;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ed6397d79e934093146b483c427ebb8bd8a928c098942b1243f4b4d4100672085fd1a4ce8a3943c6d1606ccd397e816d790b011eeb0291e063515796d3114cec873;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h182ddbe3e24e3fe1b0ce21dcc8f6fff0b236edd106c9be213b29443512ce2f3c34a3d8d2bd939908867d85f46a4ca8ddf8d3707d42fe4b255ac9102477a2f24a45c4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f86368323c9d030cf6df5babbb3806ce5deb50345f1db96127fcad5acedaade8c34d1cb3aa6d5252d1b81a5933ea1b664133a99ea30e7dc6f37ff0b8d771242cad86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe1d0cbf8b67800dae060623e3da4f3effa6fe510ad9d0d67e1d1e55cf9b04f86d0d6a44f5486cad6973d93d7c09ae79ec405541fb6676324912f03141161ef5c53c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1699658be7c64e345e61b73d1e621eecbfb1891c501753f52e3d348e749cf6fb6f4d31f5911041c43deee52d99b7fe961475813422a5e324571230e3895eb62eb7db9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16a22ce5e9ab31fcc263b8261fe62c53cffc466b5e80ef06921068182860c3f7962d9dd8ed86b9a8f28d1c44693e5a6430d3ba4212123eb14155ae9bb33a3e50e92b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ed3724cb5198327f431492694de9e96624c1ca80761f81f44bd1dee6b6c7402cf1dc71aa895061282ebb3908d38163b5a4cbb7c6970181f99151e8d2a03c9347d7a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aefbbc3824382b315aab33d7f850ad14e45d136f9e6d59196669b4e0c0c7709f650d01aa5b79206223e8aa621d4ba43f563a9eeb9ede4ef3e096e49fbf09ec92bf1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7f2c7a81d8a0b34266d59c5f64799b13593655ded176aebff4b676207713726370e3126f9dbdf5924466534abde3d16a6927747ba36af8508cc7ef004e6bcc6c8045;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4656637780711c63b743d3995658c583840dbc0fdbe387e16a18d8ef28e34defd366e202be11eadaf825002207cf0d1ff0465ada79c1ee7808f6cc7e9546dc2e394;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h92787d18b1172e0841346d689c088b98da78971ea2ced51cab623606c74dac7e2f4b6219776dfe4eda819cf480e6939398bae6c6e2df3bfe44e9206d8d8a9b274f1d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h191548d0a52f2dc88a75db0cd4e86a239111e133d9be65e203ec6cecf3eb2aeceb7db1130ba91ccc35fe3c576b8ec20cb9ec8f0fa39f3c5195c64312f3740df0ff84c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f925bcbfb88bbd6560051a0566b4c9dae3ee25819d87ac67231e31d4831636396f74f881f6b129ea1b70e6952269263f8868f1d622c39c7a4eed4e2ed10685a5e67a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haef36abf930c3f8acb9706eb5f42681e066a0b6cd2687919aa4c93d9baee7cc7e43e62fd3ab94e1952ed91a1e880cd3d4b7af9311d4e6ebd6a8e217b5e9d11b8d073;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf6cc50beeef16a1cb763b33897df30c9cf216761b3ea78b8126936e088a81d7afc0f42a401972e0a89b504da0d1deda7ca6737ff810cad0950de598984f4971f683a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175f9bfa710416481fa4ecd126756387b73c90ed394a9ceb2eebf4ed58e50f8ca0c29e4059baeee61ea5fad076799fdfd6b61ce5ec2ef201bf5a4368c7197bf8db69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h95805772e92ae9df8743c5c8e9e22f982a8999a49cf112f62936f68fe4516c799572a39306bffdd23f58c40d835d780c88c9c72468b90e6c085be47b676067116012;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcc847b877b6bddaa02be54d280e66664c5c3dda4c2a846a8e4c9a3a37a79c306d50e05b96df93c820f6979632737857d3be622bba8d14528a56de55694ef7ebc076;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fe5653aa2e426f1671afbdaec6cae8d8666f593edb644ac2c5316d22f222569e3ba7d62f32738e69858474333e232a31a70e19e37186ccca7459b797890f63cd2dde;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6abfb58ffca728855dfb5687b0e1faf87f3aaf373bd49a63157c74f435135df9d869cca81d7140c4a7b4250503e9a58b1d67ea719c4b7cc700da87bff355791bc2ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce7f410efa8b4cf1f29885b2f94936754e55ad25c906c17b6673035efd809d8a0d642a7795a4da5da3868e330109686211fe7c8c68b0e3acfeb472b70c3e3aa2a639;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f95b9bfb0f3dcf89753e94bf0c943c2887634a34c691211a11e4d46fa6446df61a8771e4b8df80dc1c60366144cd3ebb16262ce4c4ad65f0c03bcd39eb63eeca8de3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h56aa3918c16e89a9827e4c35c5f827c8eaff2a0ca94e226067f5699356309c46a72ad4df964a6f2e0b60982a85975251671d5fd5be1147e2f2812e71a711bdcf49e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3b010dec43c912fdb6c0da4eec929ccc3555d6c81fff670c292f4460340a736ec4bfed3144cb823771138360beb50341d95b8b50cd9a14bcdc55a0325fa63b1b747;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc3d26b3277bca1b0611b19fb62ff22f3404b9f0abd7b79048ed6121bc9deff7055600cc521444b77cc17509552e0f3b0d6e645ad3abb8bf01dc3ae750c1928790019;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17bce8f96c6412af42dded7a080b0ba52a0a28811d5551479b31665e7262ca714e23d20b870aeecc03079c64d830192553ddf1e0d6ea6ed529642929839e17338c8a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c79cd2376472c5f7e99848a9672377066a36fcf0a5af74f39463c30975155a72d87c5bd6e93197743a1d56daca77f35b8db224e78797face88a6570ccc8922b26ccf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb7bb2390f08c16d526bc748ae95de7352a70e9e63297f1fb709e67c6536ffec4fa780972196db6186dec482a48f10e1e4bd45d3848120eb425d61d09b1ba324a9ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h65a7296154bb75f49a413573a0d2f377cad8c5e876edf50382e16fd0cda1ec2328714f75bc13c9a70d446ce73b4b38dfa141cc356675e94a8aa5d3ea922a413e7171;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdecf67d6944cf3660914a8c4ae1ccf795c48995daee8a9968eba78b4657dd400e97c006d672673ed05d201dcdc907fce1596a0f706c47faa9139daff2ea192f4cae7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8e173f060d4e86bd37211a91382144cd91e9681bfd3386b1e1bf874e2cf4c4fe5aed296ae5162687994829fe10e5f34e73421d0915f8e19ad3be97c997e722783fc2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b84149156fd0c8c031b93ec99e017ab67898b4d3af8ff8dd01c955171913d382d3ec0f49db87983e29f3ae8b2aad6b20f511244dfa7c7feda3bb76e75ebe381f39c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103b1a48dd632cde25952d1df5c615dce6de58554f156ce2a1e4bd22dfddec08053e51463c5493866f8787bfd8537f3cad57c1d4d5589c5ad80ae1aa11c0439f68257;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2ea740a38b6a9a460ca1f83fcd895b809f43aa77823997dbbb5225d7f99708c1d95321d586f09a975217f9803862a3ac41e204463b3d0a0826385064c510a48e0eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16912cc33e745a5661c07b85c4f803c12516ab7bc4a02672f1ca565d44151ac78999045aa7de437e36bb798f372152be08f99c4b8c928a3c10db4db1b59549bef1bcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1df9078733ea180dca134fa0ef5900278df3a73eafa5644980b9263b089342af3a7dd126328810571fdf6580f201f381a34bba5d4acdf729b4aae4bc48882faf49117;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8b48d98795eae3e5f6da3af9415b986d044d3b19dd37234935aae7307aa312a95b22afddd99ddf6b8f7874c4ec90a138f4c6efaf7667a6f1148a30fe0426e51b7638;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a2e99d44135c5fb773163a0cf980e3a4e42c21ce1c08fbfc9e17e6596a90a6096d08ce76f30bcee08966dfd6cd01dac9608ed2e014d9f43df164fe9f8b0b54822bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1376cc441243447f192a26c621a44ba17465a166c302aa8d53917790a75ae398408608c8b36f19ab6f9798903fb521757f8ef5df0c8cbbf4fa2a26b61a76aa0262e41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1adfefbd7d3978db9a6e3b87be7956bc37bf826d1981775a88fee73a3d238f45d1abc3cb880b3f48ceb64564e22754102acb04e91b58e8f00532e5ba7852640070308;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b348708fff6e1be46d06539ce00251ef285c7d0a8d5084d3b7e8eb8d0ee02b825a304663dff77b55a55a10114adefd77719baa08f1947f6600fd80593120c7159e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15262d43d4e429dda913309419ebed5a84d699052ee466d0e2d3d8dc259efdf29eda180f4f47b9282b69f0cdeac4dd73e922d3473999da41a13f48daa796520b5d06f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h623b14a32be0004fc8c4a65aa91362d6f96a3b227c7c132207505dcc525f3fa62a6bf33de5c3760f7d0c05261b81710be4868ad92b65493cfce8ce2ad51ad08a1cca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10d81f888ce155ed379e9098c75a2701c4c101c14614021185b00f3fd4388fa6abd9862cb74fbc6318ee0bad719ecf678a23b9b1b5c4d741a6cb70bf50af15069fa3a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8a917e690c2fd0f2f316eab072ec91626003e6e7bde3c44c111e5692c0cd0185f2144f550461c9ab5d579e96e8cfc48be3d3e9f78edd25ed5fb286c93ff3ed2e5681;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb9cfbd802a71c05d66feef7d879bbad8607ac344e3618bf08a6fc3d4f868d0d09b63c6d7f882f9ac6a2c139ed159dfe615042248fbc7b32951449af774cc1394403d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf90574cf42ab3f7ea885a0027edafeb984b515f917b096ce82efb2ed95b336cddb3ce9835bc67729fc37daa5ab0160615c71f02a47189d64de169d33d0f4f609daa7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f348c0d7616796d57c101a15f6a1cf15ff2709fed320a98c268d7b6b01a72dcbd0aa73ba5cd7dcea92749e08b8dfba42c5e556bd316e1a181f54c23c1f568bac2a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9348bbab1171af020708a508a3f982cb3ff583345b7f0738e88bcf2d22e79965c059619dab79ece077eb0030cc6ef05f551ab90057acd924f8c5174c545f76f16c56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c0996742e97407272d1e4e0b57367fe3eaaf529cc6c252d8e332a9819beb35275feaade29a5de6483f8d75fcd4192f54300685b279c7e64516b8d4b902f50a96974e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hffa964e32bbbcbe866245a4f84bd45539849509e8ce62411c8d12cdff762690fa2eb292b5e412164cfd0fc862d642da132fc261fe1a82e53b7cfedde305a591a2ac2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6484f0dd8ffecfe1960d9ce13014acbd8be3e9c0ea9f5156e18805bb083a208c990aa6de846cbeb0f3a9cfe722f37764477a8439fa34c375ccfe1aeb4c8ccf5a4f91;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd1960d7c0089eba21f0f241376d7c48c98b41fbd7d789875712d315f04cbc5d78d4e424acc8a2007bb39b4c692b32535375a9c9892f6228f8bd4cad8ce888a2a68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5c1d352a051393a8c98bc5d69186fc0879248c2168697e52127e681fa41adc7f0216888d971bcc917ad44dfe5fafe6d06513e8e239be94ac17826b7242a6c83f5791;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b42bdc76b1a271e8c9b8c4a8d4b0c534bad42341ac461d4de1bfd3f6f5d3fd8954c0d6b97870ddd2bfb3c537f0bf7c16ef3874a9b83c7023e2cf69d4b25ca8dfc027;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3882548859de65239af5bb4159a70c3b85548574738ea1eff6d14a768e467d7424aff9a1bf9089b262b2bd2858ed1fd9ee3e14ef01c7636e3e1dc7dc54bd69b43ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h121173ccf3c9d87e44c93f58d5033024974abe8b8ee20e39b4e17753604113a4e71be0bd1335b5d4d7afb687ccd3b3f5e5c29dba19c27c690fb8b7c4b7ad482671506;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1911d6a7dc01f42ad72abe149b419397ae0147bfd0dcdcfcc680e96aec58287fd9bfa5e13b00f96cab57e0cc787bb099836cf9e53c0947c0d0e7829ae920dd9c63851;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c9bdb97471a138c5a9eee1fd81838a1eb2b99be14e05efa7b292d942d3862c0f2ca8bbc3c678049debea88063efef6fc7913c468fd76cff8c66f81dae1276463df2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c5a39c8c823065cf8199c887b4b2d0fc24fdd0d4d01c15ebc0346af18d2048a8e13503aa8d18539c00be8639495d1595ee6ae24237b81bffd3a71c2b580ef12675dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f4c08cf42163e5925d64f7e871e9a876396b9414b68721b6b9cc4ce85e6d313e1bb6497fb787e727763a524f2ec1214665ebede680f20f0a301563d0c276759825d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60a032188fec072cb69bbed3ae1556a4a72c03669f0e06bc1598ebb4531dae77bf38dbb8bc79df49c10390d024bac3683e3c89bef7813420780e0994eaa9fc02c5f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0be3cb638af1c6c7bd29759b75abed9794190c0a28e832877eb32dd4648d0187b53a7c3453ef97dacbdaffbd657a52d5da50f66d7c7c5f0439789ac12153a480ecd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h234b7b9a840212ae61cd5d272b0a27d5fde1dcd54b8d12ce2183f08866d668ccba71f0f215bc01c605e1d3d4cb4bebf16f02d9d2819c4f384e01212ff984fc384fca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1452109193f3fe6f70e17930e8cc00d3f817dddaf08a6d6603bb25e5c692f6e4e6fba6d69c0ba2ff0739accd15f14b2a0c8f8b20de790233407c6630c338d3e5db612;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12ee105fb92363d73e50d0f536817ae49934fc5ccb889e3a6411845109b5ed81664b7a5cc41ece13467e2b0fc426d636b32bbf459be367e09ca9a25c1cea4d975c891;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h150aa1379e1618399c5b58c4bf022b109371222e5ea49050569157ac16f6ab6c4bf8d3e8ddb874e8b4c9368588aacdcb9317f01a2aef490cd02533697f1e9fa57a400;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a1b11b891b2521d550373d99720e70c185a6d8abad4ae2c765ea2cf7bf77d7542d9edb3999ac534d98011d0834507f1d8dc7053755134e0c3536ebe9f1e8eba4005f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdafae8b7802dd2f3fdc0603fb491c489f4b3ea5cceb185e2f64eb58e03afaa48aa9bc7637e3c0768e5b2cfbb1c305acac9d0033aa358da549c97a7d15bb1d2f31527;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b1d30488d64724aa6e2d879401a9923480f319beabf4c7e77268deaeed9fd47ce635c6f738167e65873a23cb63fac647587f32b47e927634ec36558cba86f5e401ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5590f42eeb1fee608849ac9c8be7d04bb5550a9e1e4b3d8042beab70965b6cf8c90b78e82bb10dd2596f83abb159841a5c142b7f8751ac46f9e5c681ca3c0e7c9742;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h86f8d1c777d53337dfd810b29b0b12ab95fa2e3b91f042a0ad2dedbb61ff4303c856c811ff7a9d065f18276d28e4efc5789aeccf3525cf8589a6e7e20c58bb30e252;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h82d8a617c409994c60aa9f5ce61c289e3334514b0a7cbd4b4b78e3739c06ddea728216f2a25c57dce88f0cc840afb52a1cd6be410f5bf088f9b94ee6cfe53cf82f32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdb572e687d453b915f0db8a6e542458f9ed6c13cda8beae306f488132f1e10d28adac1995b5535d096b8ceda3a623309134ff5c44fb8b6b5fe60914d8ead973b9ee2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h114b013950dbabec8cff8d31d6a373c07dbd4b9d603ada6796ee2d77ca67b58845a66ac3a3312ce38231cae48de98fc3d9fb134c44c541923393c36da58004fae4b3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe7cc905a0eb9d538f292bf4bef6eaa7fb0160358a70bec28bc04d8a7fb9ba05ccf78b38f4f03945739c1e17cf86462576707550a9989e7c45c0568f17055133aa1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf511df8cb2194342dfa9f8b87fcca84aadc6ee27c8549b253e6d39c8fb008515808edced113cc3ec843dd5cf0403aeda567d417dc951ea3facc6f9344ec70213a49b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f8629a4caba04768c486f8e8c8cb17d1111474ba97552337afb6be5b0436a238b7503831955d77016b950b0cbd60d4d8604098e3faf101cb80bed7b436ed594eb99c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5195ce6284968c9996729a355fafa7439fdac7c20a2a35a99138dcf939e3229e18230b7ece387b0eae7a744173e2415f617b43eb2fcc20a72b764255958c27851e90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e0df2e795501e433ee5687d57091a7055bd8cedc648506846c42ca5b149feb6ecd77c4bc376632b2e060a0739439144d203a1b552447fee033da276ed6f121000e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c59a2b4579a5ad3105f9d6deccd08886b8f6f7f03f184ef0b4afe553bb38f480cf95d6711f540ecfa3899b53365e7c0bb7b317b109352b8f2ef96d26bf357c35bf6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1591fa28c61227c7ef28f5bc8d3da81666c63f2a84b0301fb93909d29b76e224b9c7fe5efdf5a086d64fa279d52b8bbefb5f5df81f5f402f0e2480d83301c75115eab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h124210c1febf306e069478e2ab671877ae2c7e96523da3680e40d2b1f91c72e933aec87d1e2b271b195aafe6e468df446c441cb642be80f30646a9baed119a271613f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12162fb607ecc88eb3fd6d590bfc9f21e2c0b38676b54972117814dd326287a1f81795414a3e100256b7aa970d0a06e08fc5e15f0d94b43ac801b7377dfdd8b859eb4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140fc75f33c523614e7c042eb5337f4961e7c576cadfce7f9cf368123681de76222cd10a20dfde0857d4c97680bd8f25713f3f8ac357e8241664dbcfb41a3c98a0b7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca7995a99385a1b37fa0d3f58290167a65c7f6e46406238da14fa19bb5e509f008e041374492ed0be75e9370f6e5ae7d55b9f493c2feb0d7d8ff6ac6bd110a82d49;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53ccf51866dc04633a009749371e366e4d2c6bee5d02748de62598b35ffbd3d9b2a12660980a836d03d500ba3641ec2ba53046e57c550f2094629012656c1d56f668;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbaa566ab8d18f94f2941f7e76dc8cc2fc243b39e10e0a62c33de81001f355155f02f627ba11a9a0c83f401e479313892d64a88456b91853210d1829281b5f82b163c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h164e5b1f08ed6723367877ecf0e79da90f87eb1d9cd90871e9f7756d7a73b48af2d391bce4f9b849197b5cac0e51add6f8cdf59627b37d6b53393936d825b43ee415c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0610083497184eb375cc0563ad7d72421f8bc4a3782f22bca941771bfb6b3828b344c72c133057c17c24f5abd9f1a409e535492df1fa6d72544d018161b8ee782f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fd19f4a00eaf4a4476351ac9e3f91b7df437c58c8c3a5834b8f3d02ee5e859992843320cdd22c180e56b3722cb988640a2da738a8d33ff863302678e3baf2da574ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19cc8dff7573e1201466701231e6e8b0520f784dfe3d7b76efe3e8272d02f36b1bbc55f4a643ae7555f1beacde884d892f91650b31e84a9b50b7ee994f3b0360b8160;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c1c0a176ee560953c1d641f3bf10e6669e62d5dcb9a33decbe3641f134b437e22f244d2c898d592dda7879969db9db0d3f86f137a18562394c296fb68b80470372d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6f56a6357aa4e45d51ba3464efdbc2842064dfffa7d187e7fc18ca87a5aeba19175df900c49f01290a4e5a80afe0873e508199c2ff5b3083dd3645db471248d80c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1204386a2a866a0eb18768ac0f7b26be74cc0d707870addb812f0bb4b1f7dc970333aaf9b1537a2bb49b21a85193fba90a2a0a7beacd09782dd07c3c69d7e93602dac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd198ac7982ebc0bb31a60bd889f80bdcc1aa258afc4c0f7abe4498aa4f2f324e7b3d46d267bbff3b5ba6276d39d747bed79649948a954dab889bcbbbc0313628793;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bfc4c98c65a898e0324b7d6f8d2b0c40e83db7c62f0c4d5714ecf2d539c0c6beb2f49bc725b4bc31808da4b1f58b9ed58aff1468ec3f44aefceac7f4809490d291ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4017fdd22be50ceffb61e3c990cc46eec8883302c53e66f0f94e98882b65d69a5f3e2575e2c1271af6b32f056bde93f673030eaef36f453c5e32b94e639f475433b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb3b484b080ce51b7611e44408fc7f419a5673446d2df143a87eaa5d91a30d1ee7c1c0acf7e8db01a512788c4955493310fc0825bb173aa1dec50d0f8bd9fe6e37102;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d90bce9563d7845646e11a97290d6fc9d3c2ac3b6d96d5283849c391547e1432412642ad00f9a6e003bc66221dcb68427b12d08c9eb65655b4d71bd2e01dcfd2cc8f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f61d7b0319dda81f5f4fd9d9795727acae16402c650f2bb774a071eaf1125402a0f9869a8faba9405db145c4759245ab988aca8e362341a86fb7eab6b098b5ea4499;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ceb21ff89b8ea8cd43a6eb0e416a72c42c55a687f19a7a9f82ae1dde40d6353bcbe4cb49d26c076d1c92ec6185e131b5fefb7020487904272fc1ffb1dac8a41eb89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14f7e706cc51d26c7d3ea58b1d42ad4a941282efbacc746d7d885c9e9223a2d1c66669b9a1ae938d835fda0f2d3ea4d2891a997d8b5ab01ddcbf1213d74293c7f5a0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1445fd317aafdda1f586c8703bdbae97f7229843c061eec914310697afa18ecfc51010af86e4e120fad551a74af14ed8602d82c56fa4b6af3c9c110b08945f89ef295;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101e1d36bc26e36847d69f746d3ced6c8d529caaa86e60a5e0da80a39e455f50b7b646c6bb496cef0ea3661968e9d4503430037b1c93d50744c0955b39c3323d33ac5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h76a4fd35f40b56f7e60cfb4d5ef17efb0231aaeb8fd3e4c4ea11d1522d3250ffdb41c1a0185e87fb680b6e75387b9461cf64396ef9b59307eef0560bb2e47cdd2355;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11de30a373e7530e6df2031910f0a57127655b4a6e166426cc474d0a300df70da73bca12783b1afd0efd5a4ab8e96ef70a77383f6a5e405d62e8685294e8447121d86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd664765c9fe8b56d5299d797d875545c743551769870378aa31e36e66b19d7554259c5c6d379234d563eb10d5525667d625e219f88b690fb81577ca7c76f04220068;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1651f449d0224a65be517b8ace5417f48912e8d0c16484df9a6e92646954fb179894ac2b195983b7b1dc43966c11f63704b5536f4f4def06e28298a5c25069535982;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18f69051230a4ea087a2386a33191f9dfce60fe804a0bffd46242cacb81de35eb5d14f55b47d91a01e6cb5b4808808338428c2c6444dea1c16e2dd99324829a7ee695;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc1b6f62ba1dbd626a7b53e655319409699c2efb65f78c6a4e899caaada295ef9b0bec7eda90103f02533d89fc44553776620a8497dccedec675dcbe34343f2c31b15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15bdf355a749d5df9e0617485afb13e7ec71488636d94be536fb9cac6917cb421fcce1942fe6eeed8c602af0898862315f147edc3ef6da1f3102cb1c98711f1aa2720;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a6f02dad2f41abb55c7b5146b359a3418120d402a762ac2bfce29399055008d096b342f67d7c2a8f3500923d247f31bf4f482f5f2b0e6b2d9bc3a427cc7c357831b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13277567cad99d7b4650b7ea6e12f05bce198391f68e0337a6a2bf788a130aa7f69d97bbf15d5fc6dcc5ed0effc05ea52ce535dd849ace4d4131d57697d3cad03d35d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15bf0262bac5172c346f84b145fc340fdbb58ac1365ab6b52ebb9476ae12b02a797e9feec03af03dd802e864ee8dba38c065eb7857f801fb251f326f655c64d2034c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e343e9007464a7955f1c6033047840488caff66eb4840fc3857b5daf78c67150bbf906dad729f8343b8eb757c284f66016afd5cd6aa42c92a73dffb58f5e66856f32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h940c1db2a802e2f1cbe8b02f5f0b411a10fe33b15b45bc46a9fdc55bda4c39df235cea2ba3218b8e05687d73d1d2f1dbae142622e11a7a0f50a1c4eb80c7c1445330;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa64a85650dd95447847b76005d84fd0213ce82091d04a986dc33e61b2f6b6d47c44bfe962ad3ca8be28943e15affdb17f8ab67de4266efc2ae7eb1e84c67b75fb8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h107c1f35a796b6058159829a697e97456ff26140c18a23b5b52f7ef79a0399b97f622a63be90453dac5f1092672f45f1d29909afdb0dd1a0bd6787e6ac81c437e81c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb4c3e32001fa16780945004189439b85b68d4c72f9013318bdb49f64f895fd34d7618e0a3298f72338a51449530553f7ee77b5f1f81e233edb12cb7f8f893b2e080;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hae6afd9665085ae74363e5266c35a0d9a0074647df6a4a994edbe3e96306fd0188b1b9a3cb6c27ecfc8ae4510c2d35d979302cee73294395ffc0bb74d60735d3356b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e5e7ed05019632cbe421649ef136aa8aa81e286460c7d1fa43c40c800c14054b8622d1ea5f9183680bcf2fd9b9d9fa22fdd1fff63edc1028a1204517549b91b9f32;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b81065044cf80c79111d9a394ff263332668bdd63009736c3d893d12a01dba3a6ba10d9105b47c16ccfbcfb8ef3bde617d95f62e42cb9e1ae60aaf09354b8f25a80e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2913ab6462660d4882998a77286f38258c0412e63649ce7e54de36c3ee90b5c7e4fcb91d900365d4b30fffd2658febe5f963a6f0307016dd6224eaef0d75e6686337;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h274f379e339bd2ef6aad364abe106c725e63f232f8ecbb71b885efac2c6d91e02c046fd229871a2e52f6bc52758d74befc710c270853b63b76b1482f0f2a6d47b696;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h298790efea30b27aad26f2112ae4541e05809e9df02e38b9d65350640fa4aa5520c9e2ab9b44b0dffbea7280d56943b7017b852912ff0410b0650d34b93d7bded9e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18d9dbb879c4a2d0e5b06a219e02737d45884fe4fcadca20528292fb32ec366ffc067f510312237bc777ad62095660ab0575c141159a46709374e8cf2311122ff1600;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h27fea8f6ee417766d990a80d5d1df15c6a998ad924d9000806ba6e38ff348aee1f47133f5a4dcd716c8ec1cabb701e67006f2092b6191ea32a7800043f7e0bbf1863;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11de987f99434b1a5749c41cd7c3a8496bb40f960398893a8af330e67d495c1c63861a26c5cc89f1d426fd9d3db6c6436a0ba7680211213b9f08624a552c39ba6b302;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h67181012186f0e4e92aedfa699d4431b23d0b08ddaf23a01feda54900c5ca9e5a58df51da8452a4dfd8bd6169e9cd7f7ceb7b40dd0fdd384824b2ab09378688df938;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd6b3f1bf5bdeacc3015675e42668569eb373249913b1faad5cb4b2c56bc96263c913fc80bffaf639ae40720fc501ff14041f626238e81dda57df4021253bc09b71c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c2e413d2ec119be80cd370c8afecd07845e759fc39637a34c15a03c77bf79f132b23d118c79284914ef6d5a4637f5888260542acfdb90b300530c3c8448229084a54;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a5324eedf1491b0efa1519e5ae3086732b5336000cf29ebf3445b5200787ad6918a313889c80aa1a7f1c6c05d9fbf2dc3cc6916c943daf006c4c7dd7778d9cd7867;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1746892a881cd9218a9dd2a8118b168f09a083971ea7d885fc73b028a54ee2ac560e56e9a88217915e3d477ab51de841a3c9b83f800b2315d39cae662118487f0d648;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d335cc652d5e156ceb088e2a5316d90cd3ef3d677b448deccb5706c0a1ad3f95fec1fe1568133aab44fb709d915315daaaf0341ccc41b47a1dcaed3eaf4eec596bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hafa7c5af8451345b35cd18faf1551499a7a158b8a8dc6832665b5e353a911f05cc339aac2c67d9ab5845df6fe4f7879d85fca88de7aba0a673866469310fe5db23aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ac84df01cb061cfab8e61ee5d923094de867b022db7f75dd8b538ecd5c82b4f535e960ab2d1abe23c56bec94d42f3b4cc5c5b6577cf2e197902e546bf0c55620c9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bb2fe3bc48fe0086187cdc360ec0a525bcc8ea926dbb30b5a092bbc2ebb2e9deff619f4dbff8dce5014918bdf0588238b0eca1a8e66db228ec27276e573303d45ba4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fefd8efe641c4fcc2625672b48c3f798c2f2438e3da63da0175bc642384202acd25f2bf0b64565f6e9acfe0bff91564cd2a29150f8d2c6627f0a9df16af9132289dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f9cc53ce04eed19f9bda61798426c9b0cd056a47d8b6c311cb3134642012339949223f61c16abd26b12f3f8aabe128343efed87d340c7d5e16f6a0c480e9d39ea6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h153bc8ad70c59a8d5f6f4574cf743ba36642b2517cb67d81d737870f102fb1a0445ab43484910c2c3da187427543ffc0af725b2cc3a76ea9c80699fc54f8cb3c67f40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1902853e5673114e10e54993ef7981cf0b5fc82cee0101b45577a4c1eea743bd4791d36320328c924f6bd3fa53794ea060a229bc39c8956d4f1823894e47824740839;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8fa48f4d9f080fa039d329be1aa04716599d3c3cfe086b0d83790128e8cf90b7fa8ff7a5ecc2cc84de85b5442b2bb5718d9ce1859d643effe2772221096171ae2c81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h51a85ccdc144254148f5887f26b02dc2198ffbe903715bb52f48c10a9526a9ee6ae840c4d6944404a6ebc03671d806bdca86bed2e386938b610362eec4f1e23b0464;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbb4c1c51fc12f5b59d7a1c08225b5bd77ae6b1c19c7ea7c104e3ddbced9e6ea8c7ba09c9e17f8589f0d0c511869dcc4c557d863c0cac767c1b9deb5eb078c1c16ae8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eb01826e72ffc18a9b767e4f3cb6f2decacbc0ce90de5fc605c496de140a17ebf84971603957f5b5c62ad9801136ca969ee22409a3b03207601ab7425f82f7311171;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19329149c18ce9863b6b07400b813124b3317bb74332b4e040fe4a3a225db2fa792ce93993dc69bba7323963d0b2b2cf7e6be971cc1438710df5b56065c5176ab1585;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5f369148c43d20718ae5aea1b289373dda6fe52dbc33ca63fae194b999170fe4e5f52dbcc066847d907ed7589a46b49be2a9878ad661a1e91ff2275138e281a24d12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h202704f7739aea9c5237442706d90b0cc2e7a8cfc9ec58158eb707ffc3eb08fc8827e9e91e45ab97f7504643156bb6188c7a249fbeabe6c73576c6cfcdf50e654e3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h415d224a8f3ea7b4ec3ada6884784dd8f79791aff492140966f529fdf93396d7c6efc7704fe9a40ac801601ae39024c76e59495171a77a7ce526bd90cb91671a57e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b193e1f72e336ad26bcc609b995e947f173e2ed8127a8548751aa36f940524edb67b6e893595efdf729b63e8779c9d16a9615714dd54e439bc17e601d71d68fa791d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17709f5fe3a71d9c726c46bd7af1e7efd7efd9f8a71ff69877ed2eed61c6a3309881e65ed9b0073555f9c03aad214bf6a129ee7a3709eb75de02c4dca1e6d0a10ad3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10539c18d7a6ebd26e5c30becb86ed4c3ca81e8fade7731418cbda0cd4b5f2e3a4c155f4d77054e52f1cea6a88f3801146e57138833d15f2ec1bf47d0ce9829111e28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1475598407d8c9ce6d9debcf0c9257b623498634333b896a42b3d27404efb29e5a511e0dede1a6fb97250fe760af9ae175fcd96c9fdf4296ca9d3ec0ac53428585850;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb71f1fcdeb7b0c53a3db75b1bf73f2f74fe1c42b123b3280d61e5d416d46aa5faef19d67cc382c5eb16e1cda6598d65828e7e3c524a100cd076edef5590f89270bb2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aea0ee8b2a3ea1dab4c8aa84767c386e75800b62e7e223e63e79dd583516338c10f3518d352b6558ac9fc402e57c0665e189571078b5c81552d5cc0fa57d02bde504;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a4b223bc11e94a31608f4aed39c0aca4d830711dd898e767e0de35fc011b33d5ebeaee18d0856ef75571cc86eaea12746533c3b09237324c781f4120992a2a659d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24c1fe65bc958956034509273132a46a13f4f6106eaa1f29b78f8852dcc3af5521172492eb632179755208ff7c8b825feb238923e249b478b82374e4edf087049224;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h167d38929d01f1e613508b60ab0468925e5cf730bb87bbe41191cba2713e3962a5bc4099bdff757ac079a1ca6a93c015dea07c83e58ce037d7d9be1ee92d6a4bbd2b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haed4f306f93d97486d6ccef1ec6d984fb43a2ca1e68aa1730d73387eb469ca274a8c11e7ae68de64f34a23c908fa83e0f17c6ddd4dd109b79dcde05091a48ca6e696;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14c4e143619a9189ba4b458ba9ed69ff4054e8a15149414d638665378e8f2d3ea22f1383848005eabd264c70004e47ae6c8a97f0ffbc0296dbb362c88775a675fa6c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ce6da456f5e7beb5c53e56a7d383bf0f3e18d599e6062957cf429688ef700880b1fc72d9e748f46522a7e74590ba90dafbf111ce417f6e6c7cdc3545c80bb2b73cd1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193993abfe420c88d41aeb35f95e38a5b2f5417da7423d8b5d55aad34167812f9b4f04b7d301b62102866f88bbc4c3a9d07bd110e5b7ece4ebf31dfadc4c1c25df7ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h978488e923012fe05cfe7229787a9bff382beb7c2c4ddfbd13c8632990c03be0abeb0eb16d0085f077a073b76807b7ad45474bbac22dd3431b63d2be8f3da6e15d20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h993b826602d3d374a02b45f0b4284de3314963e34ee5b258265c6ddf6da1aa924d7ed597ae5319dc7f73ee598bf4391f98de8d507b7da455240e399754b44e63211;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18ea839341fcabe9a0ebaf56f1845eeef784b9d8261d9b4d13667b9dfbef83e0c081257b6aa571f31b38a432f1a93eb6010fecfa7c75b50f349adb89d86e3d052d156;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19946394ebddda37b12a71cc0fb03760e6e4bbe5621ecc9a683dc2faaa007c10730d9f361dc1cf6f033f20daa44e2db282e9c86879038f4d92bab1122238eefacaa0a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e8f25895dfaa1da3d72af64a7f035731780708168e5c7809ba52767db9bbbbd19fb5af1849ad0061115f1c466a56901b87db7821c1426bca370b376f3935fb7f018;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fc0da8e0ed9ed3b626a9aee018be988647eb12e56b0041a58a6ac233f92b1b72eead2d37d0d0f1d3de82c938d1dd3762a7ea731b9daa9613871c2eaed3412ecb3264;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha88a076a6f10e0ef3f38789b06b04a2b72e06a3efd5390ec21686fb98c592d858da7f5f7fdcbed18245360f8b038ba93a0b3305ca81ba778aa22655ae855d37ac4be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b4e948deb15e2443924ab769e1f4033fce6bed2034b53c4d94a571a0aff0e5d27b67d5a43281f1d17cf563c7f1ea5d72431250863bb80c823cfe13ca370313eaa39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfac874905ebee866f3f0aa16331e789c476ecc7a424e12457d639bf7c83b02bbb2ceb888d3aa47aac881e0508e55ee9821444ed581e0571bf19ee002a1e8fd790c05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h22866e707b40334db486d52a8217b816ab0575079733b05cd8d132167ffe7567738cf2d651a647e57ec4b9d5d4498034d5b828e855ca13fbaaa2d61d068385312ec8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf81ec9386e858113c8e85f93df753afd4d6ff6045b2bf7107f817278df5f7e2131ede7e3da3c617c25f1307af482a7212733dac8cb76460e392c96586f0caf308e98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9fa086a1d0d178f3c63c5e94aee77c7b3b0d1c538d935e3fb5b0ebc58cececd89f27a61075dfbcb82ffe7c9c587de663c67fb95c3cfcfa19c6f411b9b6b26fd7164d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8d351fee77ca13355a08748e2d57ae4ed1298cac6f3657dca687513620272c9ce2eb9030212888734fe832bfc929c2386a5ab1e44b2e4f0fdfb9660376e65a30396;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb6561bba06dc71b0f58c92134662928b12bf66ea762b0267f38be60e2235671f35d570b4d2d5be1c8af5d71203fffc250282be1db954e3b40e63bb5d4955db2bc44;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e74f3946ae0c54cdc435394cf7e2405732775d91c3626dc7f19c9e920b742d047338f323ead17aee1564e8d2512f049c7557e0022ac90a274da5ddf7a456a28fe46d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf4103aa3bc0dc87f8f954985650c64863b4e41b748cf2659b62253832b430aad0d02aaebed156a2493d6f8f944cdedbc90f36a3c91ad154786f38758913c4c3b7446;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e3b96f47f0d5faa417e6b1c8791e65f17a7d3e310a1d74e9bea175512a27e55acd6fcc3ec23d31af486bb1bb3e44c110abcf3f95f70b2ab220b3d0c49530bbfe076d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h408ac4fbc00ce7d81c9949799b87c86904f7252a54d22af84fde504c906b7a87a3ee1ac3d0eef3713de0b751cd0ca4ddef5c0a3e1f72b15342b05e464caff634f9dc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18b4623eeeaeb1bccacce3d4cf8189f0e08558d7f614bb4dbc02417df54bfccfbe7a19292158ea5beb62fda7995c030177bbe1c4e75ad375232d3dbf44561a89fadf8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1613463987bd36ef1192ce42d3b284ae9eb3f2dc9f5a23d8bd6243445315c2e0b8e0859e6849980800aa4b23a60ef96bc4f1d978e0d5e433f3d80a3d48dc947db7acd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1632fd9ebcfd04a555b75bd698b6ab4484caab8211a258560265bbfe00f4d71089b33dd47fe6704f037fac8d48f257055af05dd42796e7eda54b97ff4c93113c18879;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2b2215629905d806ade9da167ec05f8306bc71e14b50f9a9f978b1ba7daf2a3dbdb7059bba34ad06fac1a348b27f54dac7f516349a17160d1de28ea01a5222f5f24a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1542e05fb12e6c2313a5dcfe8f84f2495f35d2829edffd4eb308a25494faaefa8cbc5e459d9355ea5bedfc94a4208ccbe72a7db1246b10c458e5439a03657ed79abc4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17f320961b1db34635fc8ae3b265a7bf399fd0fe315dfa97492837e7f6772d50812670c52fdc2faa32c5bb7cf475ee950f159d2aa9d46bde45c150e99544443a1288b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc688f2a9d638eb282a9debcc324d358ce937d38c88ea0e3ed485839a9e6ae76b2fd5dc2df33df3da6aecc9d4655996c4b1c8d8551a33c840e2f1f438df43dcec1fe5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5fcfa5a4d876a2a2c14c7188b153498c357296f13447e6f79a485293d86798fe126df7174d84e9f6c6c0a04d44e7fd273c1c4861f2337e0161849c4b55c09d12adeb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha761b08a2fd804f6b6a8587f9c1d341da70c20917f0ef2b09cf6ded56880ccb72a05d438d3960e48f51c6673a4ba664b6f97895e336de3d8fbe5faafd9ea30fee69a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12a8e5648a9979fe3bad969d4b39c3aaa3e457cc52f4c82c0c0cfcea11a20da915bfccea69e7a97ac5186234243968139bb4cabacb254636d7d355b1db912de0599a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14be49939646db8b1944b7293dd51c3da40f9779230da1e2c49dc202df8fad86ceafec334f897eeaf1e63ff35009f22050227b1fade09597c4d30eb374c1df2485028;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h536a2e4582e5823803529819377e152e7da83673ba44ff937c408613872ad04c895ff05384f035be86e29a25f9080325c5c685f335b3917e0289509728774229521e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h782a5208441837027a434c709e6c92349db8bda801ebfe1d2d5bbf2b6f524a34ff480270c6ae53ebb513f1f09776bb093a195681e6b210ae0aca84423c81f852b5c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h280f1299d4fbd7795407fcd42ea222de85b4b3a6946eaaca79471a056fb5fc7f75ac5c6d2f6796cc517583a02fe240391d1969ec6ad5c66fa64ac4b60a7c43895ac0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1832f545ef74c96d37f5629785711b34cf443f522b4357d4378a82f982cebe13b6bd82f7a054c284a570223bad2d014fb8637ed5f1b9b4a5fef4b3f74955b7621f5df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14748728e85b0ed04b38524e8b90d7287be3d7d7af25ec2670a2ce94708e0d2183922e8ff00afc486a31a8f36226a4f745eb494cdb6dc7053823f6897b9ae50befc7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a1cfa11647131cdc4a81b94f34c574b9c61f04526d9b30d099ac336a5b0701054c2c3682c6aaba51a4207fd957d842c49476950d175746229746f5617580a439960;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5504d06c7cd61af3beb770b4e0aa662176c2100e5fbf41fb139f0c8ec20b54a2bd3710fbf4c0baf339a73ba2381fdcdf59183ae875026d34755cd22055a6e5b7a90e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10eb6556086c4c7ae02d47417a3230411b45926a1f31ad6d25d90ebeeb2e7946e28d80833c8f386462c3dc49df7a393b76e0b73f3434b109b6199c0aed0f57f5cb7a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h109b323100058923cf162bd85eacc855d0e3bb434031b6fa38f3570bc30123b6c0e52d27f3db5c4f54ed59696521cccd3d416b8ee5aeb2d37a08ecd063ec3f7ca8210;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11d00dfe654644db9dd80a22d28525e1ac14dde0766c7264332a030a4b839bd6861b9dc78231135f0061d80714ecfcb7089e7db8d8e5d7eaab9b89e918b03d9819def;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dcde5c156a5e16633e2385cec2acfd4ad4c0048c5d839e95865f90a1da921a260b51a3256cbcf702e5af38a5764977ed347885a5ffe3c902268751b03f1f677fed63;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cfdc682930c0d0b8346b851a2f4b125636d3afb86133fdf1720426979be792134112c8f8bf0365d8c5d824e9e98ee9be1ce28ea58b00c2a98eb5af2d78cec0519f1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5f41f746465c5c845d1f4e9fb2810234e39556b398e8e86397acf30e3232e29314c3e703fa870f9245768a9cd67a901968ec7e5f0dcd32e29e326a43d43455074da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h372ddb4f654c1e9a1cb1b8cb76a0e251959d822c7391cede73dba78318c159b022c2d2d25918a4a3cdc09321cb9c7944d0b4201bbb47fcbf0560eaf0521263f462bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11be06c773075b8e7efcaeeb3e65b93de7c1b788a1391cb4fdc53f026baa25ae7887fa736283e81fa82152933fefd400943263726b385c6a2bb00716682d046ea0cb5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e4fda1f6f4cf492ab7364c9a705e6b494a17b82129e59f438db9c0e65b1c526a06de28f48b6122422fb6ea7000ceb2fcbb25aaae4417aa2d99393e4f715e009e140;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf2f38991e6492497d9c218351957d1020ad105afd3ca32c872bf25c045a8d14fe7fc5b81fe73cc9b5de0c9a39e021052e8bd131bb9f975ab32f56bc7adf91f32af90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a791077c4c07e1838da2b0a513327b55e27c97732dd9e752b435efaf93b99a55fa34329f48f66296b70f281f4ee9c0ae21d661b11a61831abd331e4bf1dc20bca11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e013789e9ef241203b8c576ba88035db12e3d5bba26c5f83ebcbd04e01df48a8b050b3092a1192c2c78eac33fe75a780d93d2eecf0d7583842994a4d0ed562a8c8fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1406014d7c671adbd5405c1b2e3e14a55f007bdd0854cf701982479f8ee8963989a5d73768f39adfbf0c2bc65bf52b3abbee0058155e31822be9b0455d60294cff76;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd38a9a66800a1c48a247b8d7bb782353a5927d3f3ca44ce9f7fc178a888f15b3852c480ed503cc11f54ace99d94330a57674e68c899de1f237316283794d2a22cdb2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c920481a028472e8f0c1cc5635f23c62661935fc7bf5b775eaa9900146887de9cd9722fe9c87680f076b11817c08ec937399d8963cc0d28558746d48bef811c5d261;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4cbaa3aaf01acbda3286770f689f6644694a6e4b7c252a0b2b68ecb3f550fc3d698d90a27ca253198bf55827f60379bf5d8d8b20b8d78c7f237fd6831181c1fb8dff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h297ea9f3404882d8210cf0f161f132a268c5fb59748f65156b764429f3d5afedc403828014cdb380fae9f28b0f536423046e8760a01c5d8fb889bb3301c5a1e77ec0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f89119ebcecee2a0caece63f136b4330016692f83067054541ac05064ac851a686ae03036d22e27e8dd116b2e87074e495b5ffd8f33a0ac2ed5040577e7b54d05c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7c4792a68fc89b943996596bdaf0f54d94e53f94cb343b43b73101e162ae9286c1912b45c22b545a34bfb033f14c7380c1a6d8573ed7320758d6a4904ed55ab4c7e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2aec35f5e468fd656b58df0a476a9e54710d0840139f0742872e36a6796071c6354145ff78cb9885e4640765135be332d13ea58e53a26cfd548e8e0086c52751c32b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d1a013b02c8b03a2d11ae8ffe6ebedbf9c23464b8989ef2f36a4e626de2c9570e971ba0646f6c45e33a56295662a3b9c4a7597b17b8633ea76c3e4551d709fcdd410;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hec09b5b839dcc881db75057b6efc52541c2ba9b9cf09feba09e1aa9b7a03999e4156722de7d45c7b7f3ae6d20e25ba35efa312895a5dd68ef439177319f954114e01;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h391c78106306f8ae66f25d290635ba19efce1ab988faf8fd27a0bd3db7380f6379f7e8822e16376bebe7540e999daed1c79a1b4b9575c02466e350fb221625f5af4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h194fcb180a982a7f8fbe93c3644cf4550f7701d93c2d6e57e0eab98724e0897fc0024a84e075e315ef997f0179f1eeb80ddd62d3dfebef537c75210054f6f68302988;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h795d7a511289d7fd159cad562273eb5b2cc62dbf12ef03ae8eccd4ff93afd5697ca1699951c6aec33197924976ec0909556426884916d0243fe5c0f379a72556f993;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9aa4a7c3a1580f225720ff35dfbfe382ca9ebedf24d63ceec314f8423b7d1efb1cb7c2db72d1554adf7a6070d5f0d4fdfe8118087a25bb57d87cb778d8ee7edbab3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16315a0fd207d95ab6095ce8cc8093de3fa767954339d3c803760b8195a9815ea35c748f053b2664c71deed80afb4b8cc916b8487ef3d3c2155e91aa48792db492d15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd48fdba4501e8ed7d731e51f45ed918dfb9cec2e9ec440b48920179b6b6805972a6928ca77f7906355a981d6e084e406af998bd2a2bd5a1b066bea4cb3d812ef8556;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdf784497be7353f9efe8778baacbc4d35c405d68f1626d3dd6bbfa39ee5bc6c0a7f831ac195d69c1e5e030a669ba0e023a7546d1fae05a117fb8b16793620987636c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e412711a7aa2388bd11db765fe7c0f76b2f3aecafe191c4e54d6cfe48eecfeee6d1bad0e82c8ddba43dcc07ef5158d4e84b2c233636f6898d7cbb02ead181a36e44c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9847aa06e82f017b69f8c9932012efb4dc0a76f9ec5de2af8bb079ca377f6afc88f42e237495c7914fe4146af4bfc97ae8961f634c5d8a666602aabbab1733bcfc39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e8e877d9a6991748afa900226e7736814014b1885c49ffae9ebb8f3e756fe187e5cd8df85012f461d4b2b3d7e85b254651822805344ace6ae713996a4f0d839ae3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd368f2ae224ca07fbbbf64cbcc45b9888705d672a47bb571456ccc88dac984d9f2083e801b2fb28178c21cb728040b97f7488944082e2570003a7c75736a82f04624;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he7c439cba0b4d32749ee4be31b2d6e510645468f7bf6daa4d1d139b28d651d4a5b4062cc7f26cf2345e513e3187d59bcaf4e82664e998668030306eca9aaa84ed49b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h117e3b5527f7f9af371e993ca39d116600c898349424f1b9daada7cde07e5b04f4ce0a8eb75b8cf7db1ed3568d72bbdbf8190fa66e96218215267efa3afe9aaeb1962;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1255576de71432a3e106137dfdf4725608f2d7906ace5ef8969a9d781e5d19bedff67a3564e304f266bc072d53fa3d8f3c2c2719728889b41b67acc23c906ef157d6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9ce1452596df518ad285b4c95532d6e0f295f13ec99c107b60b15bbf45a1bc092a63f7247d54f9c881407a169cef08f5245a69960a4e7b703cc3af4b02121c513cd6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14173657e75472694732a1dba455324462a196939bac0d8af24f9e70e297ddb4243afd2970ad7edc1fb92430c70b40bb680e5fbc66eef488397a8430a1b11c22cde8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h189b469953b1106166ba7ee6baf1f9e3faf241f9d0efd061eb311708a7a57e9fa0d9c285390315dda8bb2805a9bacbe09608c73b1f54af707677221dd8047bab4782f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdd93552597d8dc72acdc305d4e454d7bcb904c08251f04f806e0951e80e2a11c1320d514ab45596c3a23295543a638c63e2ba460ac7de2a362be327b571ce6449b18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdff7f5631b9143cdd6b88f97a4a8c2b39be045de668dbf7ac1977ad4ab2c1a4af99e91383c54067d8ee88a1a178e73446a50414155566e28863b71a8b505e2a08f61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h103708782352b3a3f36c04e911c5590864a487f088d1a5cc534a62a96e08150916b3aebe567a1e4e70d563e1aa1e58125c175c6dd7d0729aa2fa2205f74b46581abf9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1020a12d671b892fe0d8bff809d263952e96cc0d64c29ac73febdc7c23164c326570e32a818dfe154ecc0bc533962f913fdc7fafb571ecafc85cb9b64da76e7a6e9f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16931f8fb9c06d2a96eadc7b158a1a384af1a87590aecadeb1bc22d412ea793d74005e17c081893f208ac9f9a944be61f04f88b6a81e98abb6c6f72db2d624ab5df16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h691c17186e8259daa0fda1a64fe794daabd181cd6ad43d8cfaf7502214b0407e0fa4e48505995d61196a55524b7e4a3f3c7cec5e7e5722a531b6c541007a10030119;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b6599a0f54118b6a3a93c416cc611eda8b8844590d9049f8368d2f41d6c44f0ce3d94fe4af7090e30b1f4e14697796a978bb3d3b15250f0c626bf9d1f271268327bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h83da275b8c8812e6c826b3e357353485e4e56551391ecc0dd80fb5bb149ec396f73eabba3ac66fc6693352a9099cf362e8d994d75ceea5de3674af96daef4618c8b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bcf116a0f6082f43c62818dfaf3b9965e5bc6c7a61b886d16f58c6ae52732cf0dbd62e6a248d18f1270995ba489658be8b4af33a621237985e49ccf6548dc0c8fea3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc73fa1d746a60f035d43857e8e1454fb5e7bfeabb94055548d542d180cc1c1b2f118a9d8e2d4e720668aa7053750e5e7de535b93d4219cc953dfed04e76bcfc38a9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f2633602cc20b85e2f3dde15c45d5a2863a39a2e4f6fade7530eeb9603e58d1399d5f8897c76ac83e70d4242302652d67878e6de8081f8fd62573ca71a2d8a3e9d98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h113ba5ece2db2eaafbc2f4eba655798043558ad5b75170547422deac3aa29dbebaf68f885de5f10b3133f33ef81a5c59cb7f2dea0c72392fcc99d3e7216ea0ef2d5af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf86d786a69fd458814e46d0993041a6b181499d964ace03cc604aa64eec181e87525f3b235b12c0e5b62c5ca8533430337285ea1b03265c8227b68576b89f9dc6894;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16aeeaee8f4167319d9c699fa90fa47583ee1906a4b5db95006b6bffb8c8825f29a5379c37ca467ca10ad36d54345f15c201b5a6cf6f58c9df1fa677db0efc1db3fe9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h33fa2262b94032f012914b661a6bbee7efc93334f56f5dfdc49d6d37b32c749715d7e5739fd5487ddbe09c653284fd1c52cbdadceb71d67e37706f7d55dbf1491453;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb350fdf2d7484a59ea9cc522f48a06c79b9faf1a5c2aa12d1b0c598d45906d5fd048bf80d32f99000fe374e19d3f011e2c9b46b10600a1e630c5cf80eb3f7cb8954f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha6ed0b9f0a408eaa7c6580f023c42d57921f1729605de0043d66a2d46961b3e09fc6f507a1b6f9f41979ef0cd4f46999c3b7ceeed1d82e2bc54418a91a6d0acfb0de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha5eebca4b0dd4fb272f662e6b9216753cc5ad465d4f99c4d61601d29e6809d7be406ed61c104f6715f9956e5e64d3d4ea77f45565c146f2c53b42841c48daa8d1bd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h99ec6ed03d208d3cb43e94ec7ff82175cc75a57b40833699324f1d60cad82b946a01f225334c692002c1b2b7746fb99c33d9875a40eae3c347217b69dbc5631367f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10305a9e65dc3ad4900b273841de7f99936873934e7b070f8a71d7cb77fd258c5b236ad10dc1293f1c6716d78fc0d25aa0a0ae6add39b8e0c71000ebfc8dc21c3d4d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10b89a79670496aa57421d1227ff4a6611728d67ac2e38b1aeeebd54f1f827ebb864b751de6edd4b03b8439bba1a747aba0777343fa2fee33ba99408752c79108668b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hef69a522c725e680adae667a52fc93ddbbc51b255bc25a1a9e47b8797a7b38bb5cb3858e6f441a497c9de442dc4bb2aa8f546d7d4d1d3bad3e1c63dd6498f06b7b6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1798efb3f8cf0f7304ed6e246f9271b0bd7b8d3b0ecca98e1efc1bfe42aa98e99d36dd3dc0f5bbeb0d7347c2a600627ac95586920376cfca7a6cc4fb9d7b178e7149d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6fee6c9812db70079f7d31f05504514795bb95450ba7f48f8b1144df2efd90994dc881ded0f29bad19375b97d81091564aee8bf5dc07b8f09def23bebb2b2174148e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h115a0da86bdbd27a70f22a43638673ea03aa7329b505ca6e1f90d48ee41b3b5996d645a0c8dcac969de842da01f0928442c75cb750dc850266ef445f4343135c2214b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a81aeba6a586d999518b8351c44f964fa4e121e51534dc69cdce70aee5174ea16374014b3cea0cda294f07b12a71798d6b1383dfa4a7d0a603741afd7255e145908;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7716cb027f500692f006e164b308e6e900f63494dc199739f2b40dd18546d232cba43d362f23f2bf33a464344a2708bccaaa3c2a65a9d7362976e6e4cded9745649b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf6ac12fcf8596ab756251d277734e5178b49b67009cb0a143a2db04116e842a1581dfa2371cbd2bc2ddb31875a2bf946fb397e89919d44a45b2f95c3ed0e0d5bfcba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10054e671be5cd409bdcb6a87af6c04132188e49c603fb29773f83fe157b8e1b234167c44189eb7b034ba42439b06e248c2e8525fc295568dbd58e468075613ce9254;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15d8f37c27b77c68cc016b0343ed2399fd24f9188174e006f0154e80fea61d8007f8742cb2ca72e340bfc1c3f8ca5b3f4e90618b76307762f2a0c69595cc0d3ed614c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c88637d34979dbe35f3fd6dfb862cddf8e03107edb699d1ec93c6a8c38c5bb83e0407743cab0dc3c183d3445511c1a1591ddad6b80e8b77d20dfe46ff07d7fbede2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8f46132b57145121846e999fc2362d9c2f0925cc4830787475dc75280d7b1b920980e3e3c05b3a571e63ea84825bb5144502806bd9377ff068b1d43d2a6f070abe71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d277c9680950103fbbd041ea1d58336d861d5f24fb54136f1bb0697175624a98df2815fb4afbffd9b89bfdbeefb2b9e912f794a740d16fab908b334100841a2f24e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h719d6eefe8436f57da23d6b8075d8d0c7b1f6db329bd973f465d6877701a9fa5c878c14ffb093bcfe7ea0bc3edd61b3a22406da778a586974eed37b45c58b01e88bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h453b4364163600d783f86401f77b0f152abade92b64506f96ac6f493bcc86308b2d99fbf76bcc007610eac6685f7f03c2befb5bab31caceafd80384b8831723d2153;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1752501934b81d0173374ed86b666fdc26908f55ecd6a6b5624a86a18aef8d12e2b11c8555cc73b383d93066171fa55f8520f95713f790f73eac3d464d65d10b48696;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha453faaa59cab3924cf65489a67d2aa3f8c48bcf0ec03c14bcd01782a7a2bb421e1f64a85ed15e18719527f3b19fa364525bd29a3e8aa0f05ee5bae2cde3139a0e5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18e067919ed6f7322928abc9f60dc0a1359eb55353b9bd171e928e0957334e1c7256797070780bef6227383b17bf916387f1da02931bc0e99530317d54409a9468045;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc120cf3b06c521f54ade05cdd48f9e07f32944ced742cc71cf6a3f49bab7818b0996a359088f96f1ed519ef831392b5a0087ee6bae7b53ce6b3f9c8edc5677926529;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4af4a8bd147cf66dbb6c71ba78613baf897047dcec75b321119f8992f20b1f543f7dbda597ded9d9ed9f3a4274f550fe5719cf02744a664653f554f0dd124a84fbcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11ce78d0fe4a6e63a10eef180161f558df49a949ea704d12eee600b1d12ccceae8509c99440cc903e4c89603efb682f974666edda3427b6a9a36fff6cad2ab33662e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb47116ca0187f85ec9958eb79aab33e885c41f0c52cd93dd4d39d656a782cd47d5b834f192552b6bcfaa61419c02d0138ae67e58ca2615d3845826a7612db72155cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h529557628f80fb97a3cd2aee7a84cd29692ed57d59fe08f9121aad571d504d6c072486a6abf65ff67983008838e12928a6f5805900eff25cc8545f7789d1d0640ea7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7734df8b069c4487f28e784341f54caebe3e97e164a0db6f8f0e93e56a558ebfa858f704e6ce1c0be5dba80ab13cc9c493cf0d136839d0476f5d0f9a6b6c0b5307cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdbef41d78a47a868c68bf0d51957e4fa4f53c5412ceec3daae05b100b67954a743d2c5b005f8ec6b0543617171735a0774c253843ff76cc3b12696e57f6140beb69a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dd4de35a2bd69e4d4938706f688ba24e8c0ec4d05d9238e391d44e31f74c3c7557e38c880179cca22a5b51efdc252cc044d3510eb58a800e0db5f58092a4d397025;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19630930161ceaa2887c05ce4d824570d449442bd6b91bcac7e2afff0641af7140d8933d80badbe18424a26b3a3a8134461923c564de4f3d63f7deb1d17e58c35e31e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4717b56944e50bbf16ff49938cf694031132506b3c2c556ecca90143967a554f9f648eface5a8874fbc9b11b4780f11e3170a4be25b93be27f7ce3eaa339dc6571d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hffee85e622114646477d76dbd0af9e977bd985a924572d52faadafdbdb52426724156aadc47d2b9b9e9c3a3e22c4a95a0390b7f1228f89f2be3450e7072d65fe3ace;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf62cf9bf0f629518143e4456633499a475732bb20adf3c8a829e2694e9c92fc524fd684008dfeb1369f8399a0d40ee9c6d2fa109e299195d44cab0264060234be29a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2c8402135d4c3a3c264fe9fafebde5619e12d6c9f72291db59d45019ec698723d2735683b7d6a3fde2bf21cdda01eda63601dd4c2fc4aaa5035f5e5a13ad1e45eb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h131bb668605b6c989aa732004f504cb1d64503ec1028361f9b0c4099c76bb8df0de3a6a1421643153eec8029213a8cc73cb1c61ddfe90eb3df8ba9544bceab7e8a6b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ddbe4249c1f64735359e8525098ef45e23e3a4d9e7c24a285129ad6cc8c119eb1d7511d8e181850bdfc50fcd82470be24a16026fa0de89c9c3bb24c3446e8542692e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110e18eb7b0c3a44dc0000803ff3ec0855880870f57138437169107a41152d1541327b3ca8a8d30962cbbe5c63f4f534670cf198308e86597a81387ae13ceaa1767a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h196c43fb67507b42446658b8f6e15bfbb2bc4ff17040938ac710c6d737c7a78f75b30d04cd6f61c8da1df402251be780e57a7a509c5a978330dff8a2d0ce1cb6a8b64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17506b60013fcc3d55bddb24b1fd7c54eb8172ce1f08edcc53b6c736ba6ea6ca426f6d29e1b0b3c4a16e169204be0b6eef7be09f3d7a4c9b767f4608f5838d874bc05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b02477574dd27c52686c05adac757e0d3c10d179a8d27bf1337d84d18ea7837d461a8b152d53560fc7801ab3ac8d4830b91bfb94e0ba22190d3f901da71e5d78d29d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c5152466d430bd4471c5c168348f0ef92e09547cac3e6898f94b73017df257b15c83e9ad908c8a504fd1577fb27ef9f67388c6845d275e253f87656214efb3949a6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h179edd0bf304412c31967d60f8cab5afb7d7b0b1e1eb09efe4b06e97920a961c96042985c43b68d90c7a6394e6aa8d9f36fbeb6c8c82f261c521aa3ef4f787c3507fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15c3ff5cbd84975010d6ddd42a15db7830bb77e47668b07ceda1a61aa0b0c34081d86bae285f9d30acd2aa7fb531215a5a3cc858b33b4bf8f3dfbbcf2eb75ea9a0993;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4dcf57ed9deb1a8497a8b28531bc9f48571f2df591d3f1c9be1b678ddf54f511d125c1a6303cae9c36f76cea777a0ee314c6c7f35cd71a1611029441d2839be242e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf0f84cc62b1232a2a13de14874bfadabc2d6e1bad93a977c9cec9d8816f67e816f9652e478aaff613dbb7c011a7b4ed05ac9b2d881ad14f6db5cf0a2ce1386d7d9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14001d159b07bd359f8168b72bd06a47d926214e6ab60f9b187aa4dafbf72450c509af02e5a15e6ec36eaed66f7cea92259f9abed2a2b62843a5d2ed4f3341d6f41c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7a3dcc73ee7faf34e4b79dd27040601947d5329d1564c30bed296ed746c757c060e99428e0bab989b815692dceb4423ad45982cd8dc3d51de487589e916cc41ad1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a9224512a1ffd0cf182cc5fda93ab8be62825fbfd14c008c4d785ffff76b9013244657ac02d753d9a60887d05246f55d1ccae034f2f57601ff3c89e4e30c5e2a22a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19e8f4d4842554900eab5e7b1f3697051eea40c126868d734154ecdb5a723eaa8a20efb4634355537a055ed0ad4e2ee6496677f829ab826ef1103dabc621ac001ef5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h111e96c28803a8df90e73ff4a121596d6c941c09c190664fccb92d0a6f9fcbc4081049e8ee75dd7ea1799b599e503200270b2cd05a256e0c9a719973b74f4c3600e24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h198b83718cc32b1299ad51ab1b92f542c468a5834be4166ffaa97775e9664aaaa162b7864d0128cdd050f72c581fa9d9806d75e76645149ef5e38019d6dd0b0758514;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hceeb00190335bbd90fc57f7d1f3a4c9f32c2d00c8085e95246a4a92d4ed35ebdc74161a125d49807c3f97449fd839ad2f297a87505f4d0d7b0eb547c9ef98bdd1431;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1606b04e8389849e0c1ce8fa37beb76f315d4a879fc6c544cfdb429fd31abc487da413890b3faa59c89fae895e83a9f6695aeaa4ed918f59e36ef45cb4902f6325d24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h60e2ae623dfea67546d54f113c25b691df0b582806ead2f76fd76005ac35c312a9b00fa37c027a9144babf9aafcc3d83a093d222917e659b503ae5ab4ff9d6fa7f79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140757e56ba01448e464f45370db8cea4abb5db4d70efee10ef6978703495ccb2dd15bb627aa3344dab944e1f12594fb0d41adb99194063d4b261f846320324f541bd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f6102d016a47803151776d9b958e85ca571c78043e84aa25729c6b881d4e2158007258cd2625bc13f82f6125df8ecc5b8c4e0d07775da92ef658649f4f186feb82da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d2a4db1269893c256e4f884976190df47a0fb4e3c5148258eef1a2c117bc6d67786f76165a1a972dea80ad2a06006d98dfe67da4e0ec61073e6e89119661d2eefdd3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4a9ca69a22392422b8871eb874ec7331ccd486e614ce5f0e5a10d284ab1bd42540f0f0ae289dc8592c5ce984555285529d47a70e70469e86f30c9b5aa88f77c49a21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ad3107fe29c72f9346b5759c9450d578f7c84ac7ac9ead1cbc11f2c71a0d181a23f37a5b9193ee99e662b2e1a87fba49142629d8183c7b9fbc0f3772402a0c59329;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb01ae77c8d83bd384d99da54f74b19c613a7ba151293e7e020aba8960f794ecc636b119ae62d5b4439e39f2a5734b58a3629f6c5d36cc5288ecb667b35bc14fbe1f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17ba642041e057db6f58ed26bb94be88bcb41410967fd77a82d3b5520f2d7c7c44c989b1c9974b97a4a0127a2ba9965c981c35a658d6d3dfc0138fda68a6753b3036c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e162bc7b7bc21e1d0acb7f80417e82d2f7bf6a5dbc1c425540ffdab7809412913a540dab0a6df82fbe270d417faf9c865697de2feb854692beace43ea270013b729;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h163be49f2555df21f1aaeb1fd67ad936c09f1f52a4010882085a9a61c714bc1cf60d42eb9d32376a21b0f0556ef2a7c517a03985e19423011759cfca6b380afefb388;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha0a2fa623d3982bb617a955d2a2ce718665a289ec44065def0e11a22f6cb0be03a9a49033a7303ba5b83d2c8c10ad52f94a1c78684c79fda29fb37eb9603cb878c4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h909fc15de6f119699e8d55f7d26de0f654d2c6e34d1e103c57cf8e601b411b670725da646922754b5002cd1bd9866dbf925ba37c85d3dd8c55ea59d6e847beefa3c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc108083cc835fe12f0be50908ea831b5c465eb2984324d1704acd17b59425f702a1c648a830853555e2e09c4729615cd2f0e60da61c26486b4c2440341643d228fc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f91ef3b86f8819d1be0c47a749e5650ace8b1456c6ba74d38098ab732e324d4047d7386fbb18547a34958be4b1bde6e25d64ab3998786ce8a4e7d74c914f4e9eb912;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc2bfd2f430e91c5d1f56fe1ba4a3e28c10569ac1a94212e578cc71f3f7f8b261778fa4e0e2b20e9c05e79833437950b8d41a70f0841e5a9279b54478ffb3e0271ba8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f241417b55f084ea6693adbeadeea6e92dda43f6486b52ffdd6d7633bf751903ecc0127d9fadb74889254b492fd4bab22d50eb7e15ef879da17c90ab9b8c93df13f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1115cf3f8c4d0afec2769aea2553304016314056f17c8cf96bd975017003b0967080f63f80fc6ea741804eaa6247ddc3647e2a867ab0c425233438a8fcacd08f70c45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h127ffdae385cd81719eaed81d2375295e149189444c017a0ac597f3c2a6364552016b5b7dae9e220518b8ea501495ada2fbdf9c11426ef3851a59555d2e0eaf839807;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a5c96b639088d5d929f26f7192ca8bf25c733973fb500c72ff94a90c311ac5ebb20499281a060edd215c10cc460c4486efe63033f88d058fe14e94a1e7f539d3e5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h765f4d03221391a8c094125c9258b35e9459df7bfdcd430deb17e7f614a1a1546ee495b180a6dccb2c9afdf6c91d712a1d9c8cbc9bcd84a54409f63ebca6ce5269c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d751106c4ea14e0ca40471f7a320cab841717148c36506106679035dc6861dbb0d91b8338fe8b73bec650c70e4d569f0ef1af52e85fe3a49df62459028897e69d37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17408488f67d6f4ac879e8c12bfceca45889f01c5bcc62697b4478e9b0f0e351905ea1e37e74aa25b67f14d05aca1b6193494702644126c98cbaf183303b88b728dec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11d812335ca6611ccae2db13249dfc08bb91f3e3a55b7be979428507bd653b7cd44f049e8dfe75348983623fdf2708dfdccd935d7b285bf0ae764404e6bb3773b9d56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3ff646a7acc662b6a44279b5e0da1e966ad4d2eb52bd769112c15301327309254494efb37462144bde918beb7453a5637ae3f67ddcc9744b4f4af2f7e11f34885dca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a5da112601d6e703fd3fba2625e14dd7f84fa434299571e1ff1ea6b5d0e4a5f80f0d8d3651f190d925829dfb60ef4b0a7b334f210d47b8c22ca430d0b05bf664cf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdbdeae437a047f3b0471f9d62dbdd528eb918fd29f4baf2ea5cb7b809d4527d72aa745eda591b08157992ab42a1a249849232ed6f1aff4c7ad296f530c76797df3fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13e1d1fbd4f6fc5171c13557da514824eb17ef803e0cf2464ddc958d41d7dd906346f81ceeb4cc445cc2d5584949d1d14be7fa3fa243f1c77935573e4a78bd03bf139;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9ee51e7b5fd5b8030ec5abb2ddd4f3f06bd0ebdec53a4845441eff0d56c4fe0a65a65200247b7ddfd3c1665da2e40c262ff1070feb0af32dbf708551e40c5df04f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h456384e3ac25cc16cc45285b3a16d1feb44a8bedcc5fa5d92f761caacb1cf9f6c85f77a03a324f5b0964a7a6be2bb4d2f906ba0982dac7316b9db1415763e526e196;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d7bff6e63bdd65904a0c398ab24988142ac903519a7b8d85ca81261b5d20ea576fe2aeff589a39236aa3c56efaa50253fefad69bbf08298fe392d292f205389c5330;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h234db7a028469187566f87aa0a22a9f12a932feba513f6b6ff6fa5a6ffd6b6d6af41465249524a8d3ef5f321e3a2e626fb9e00652f48bd3e9b4db1b2b54e27b43a60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h48fb5d1b927c20186755e5afc3a1e8ed39b45bc9ec2938c333802f09b751a80fbef15b812a4a56612bd8063474858ea9b08318dd05a15d6949f2ebf8c227ffb03c87;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a1af507657f941e7c35507f4ba74f109ae1db481643d2a7f82d196ba1ebd3efacf6e778171d3b97b5f66076164de42d112198114c1faeb1f86e3f20492c663fc854f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h159b1a80ac4f8a1579a9384c834f4d3a8c192e5e50553a6a0ab5b83d86cd0ad5013e1c86744a3e5381c24268b546fffb7ff53b3af531b12a55165d9fdeeb9d13007d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha24fa9fdb1229d2c78f2beae7c9ca7264de70208ca77a00fa025e33000673db3d5257b1b3f4eabeda562efda42206b3215c3903ceb39bb24a1124f27689d61cf0fb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf0a76cf47f27dd52f9c005054edd3d76d052d78e94680f9d8897f7bee4179247bd1de07f41811b67b80d7149dd5f6cf5422f575b02f6dccbc371124f1ecce0b6423;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a0c48cb97498df62fec25ea56dfea70ae5a7e02e6b4bdc651ae2b9bb54fdf599e7454ae1dc5d6bd25ce38d9c9cd94ca442986420a1793ec10350110d232adb4ab42a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe31ac536c0c31f1d26391ce80378de85052794cb0c0dd09c0e6f7e2b76bab5ba284a7cc53db816ff4099f437e167fa53d712e178b6eacf6113ad183415cec8f9f3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h355eb08ed89bb381661cce7c7e1dd35b2336f4c5d0fbdc47dec067c985e10758cf84680047f197c5977d7f31d4184aafeb24fefb49633f418b3391272a0216cdc33a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd1bbaf23dc412aede8f8c1c741087273a245d2aa70a795b9d270d322088fd5bfb66c60624f7bd832edbd87eaaa95adbb77c2f33c0acc75fd660cd88bd2f439e0b753;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hab5699118368d6e3853d819fbcdff8eb1d73821d7388a5592d03c10236f1ecec4ff8342e8fe536263ea05dadf3144344dc24078cbed6ee9cc065fc0e1f0201e9509a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3eb9bea08de3ac327aa5472c368cf93d552550e1a97d85579a29568f88e6ca724df5a675c1bca577478cf181389db7ee125d14f498ca1c3f74fd54adfcd82ee689d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e24d25d767feb8723a4eae3b068f74dd38dcaca288cd74744a7e1caf07fbfc8d181ff886a482fd27cfc506d566acc82b48601684957ded094acb94406dcfd8b3b73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1659a9750f434250c924bfeb37f42f8c5e738d7f13066e2c154b36bc59e1366f80404d4bf0dc8b908e84ca2660002b944910ca74d25e8d51e24e6e2a10984d5496ce0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h185b08a49fe8d5b89d910dd93e85816b1de39c92c62f4c6325c9cf588dac29dff58d866a9bea105d6021e82ee5173b8ffa072cc1e7b0c23face2b645ffa1d64195f67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1840270bc9b52db356df1b80b6173c9781a6a7c44af665c550fb7edd40744041a1b842fc3c47cca7b7499bed5de6a102c7e80722f6890371099e6daa30e9fb336ede3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9a9c0905af445f5c55a770a7c345b42dd5b48b5fa2d3a49ecd6c5f4f2796b9410d4f182a2dc9e3936a40c8609d949476c1524d035c5b150d4d4577c9bdd09d0759ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heea066136320b8c60cb424ce2933781cc79b553095d3cf3cbb5ab4a22d72d16f4a51a3156bc76d8fb0b00cee73b2922835db56c4757c5e5a150a7bd3dff8e580e363;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb38008096852110e5ad0a78e4b9687761a9f19663a4eb2147f9f2959f32e7a25144ecab4a0aea4d9a57b0cb46bba90465c591cf21b5ad09aaedf6badddd9efac7c94;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9fe0d40debc55651677793b3e2701c8800dd868a063d029e2d22396955b01a504fc8d3f9bed0cee3f2de7daa53ce5608430a8812f76648c896cf485a74f8138d8539;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h166d035a418092e4b208983c84294baa439ff8f9d53faa47830f2851d6b70c24e42d6fb5dcf8ef229cf376403ddad97ceb60774ea841bbb569e323e63cd00b9ebcccc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb8f41bdc8e300404d61c7d9900182b89b7cfecf84549c4ed5f83bef9f5ac2c0c56b12b6e5b12b4866671ce1149761b5c539fb502d0d7684d2687be983e05cc6f6063;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h96f1dd93534fed2901909578d557e46e29f156b08a383b5bd9187c2bca6da39332cf450d12e8f8f01ee559891411854c99de68b4c6efcb982815ac571479fe7a46d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h159357cc2db611d2985c13f8f818b4767ef9790f5ce58de3b7f17211f540468fd252189288d8b2690adfccc489bca1f1184bb92ee79cb0e3cd409665789b7555678ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2610a80f593f838449d3206376f77eadf6e2dcdc8f7d1b6b5e20f352b3dd9ae194d98c847d49f289cd272ce25988688c7cd32d6ea0ed6b36d596aea372429fb306f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb2104f1d5194e266f1dd53a56b75de7beb1ed3b024ec18eb1d5c347b3ad5898ac3a1a110ba07d9bd323db2457798c73e1df3ddc4b8449b9fe041f7f4ec20a53503b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h68950af615ae852a9b1ec1f70ed8b842264e83c16145fd97b8aa5108e27615f5384047f09b6a4ad2d6bc5dd75fb57415e7d27a18f631299307b258807fd9976fd2ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ad9f7b04b91c7ae38fb106917810a6f5f32d4434f15e20c0fae0b154591d4f72385f90ee373319794c97d270a9f9938ed3a0e8c7eeb46b05210aec0d084a9827a9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1827bd66267f98bd25c1e6aae971df9756c54f06cd531d4fffab09b75ed29b9a2b69ab83b3cd85f221c6b80601984ec9fdfb2eeddbe8fee54592183e1390b12bd3813;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4799488a60150c728daa798d259942b2694665f2f5a49f2e61f2c4838f8e7f27d43625808cdaac09d46f12c0717fc766a58c1e2ba05def123d2cff9b4254a52d1880;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15ed246f65f3eb7d35cc05fd1c8beae058da942a0bd082d9d6a09c48a118d15af3f9b59a9c2a622c32fcd94948e5beb4145ce7651f17b2c065e774d0b85c27ba213e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h24a3c0c3c2178acec3ecec1fb98932798fd51b8884620cad208cca7255a99ae1cc192d3f5ac791acedba94eda5a899ebcc017bd4fb9b441bb2603d3bc52e0ec36351;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1aade7f5ddc3adcdc63cce1ecb24940033f5148757266d2a7c5f59b97931b1dad4e4c9794e63ef7bdfa0d3200cbb165dd8de06d7b46feaee9a6a6c10a1cdcc47ed2f1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1014e96391f131e48ae1029e026e4b2ed75ee465796d3c2ec1102d59d0a0010e6b3a61ea46ba5df7d963dc3b10b7d675a3f76a2e82cb88a321089fd022f64e895069c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b947bfc2341f5e38e1feab4c3ce59f178c8ec541e16f4e83342f236613be34ca0edfc08c24b73e342cb739b5fbe63a24a53615887b0e1706159eea135c8b484ed81b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b8681b308556904154dd2063460ff1ef13816da2c52fd26d81d959db9b19d75d44b2655b95fe21682c54277e75be64316ced6fc5c47cc4b0d64c2ce50bb25783b71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7aebd2429ac15e7202f0de690a16318369b7bc77f708f47ef6ab447023b13b1c148fe41e842bccf288735f055e72db3ef0605f0b4a592b34f3fa1e927f0b29bf8db5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'haafa22f182e8087f3879077d109fe4b4030c50f8bd2a13479bfa72ca51d66528d65f2f7917cf489e617ea8ee91276ae7e7ad3fa45dd9056295ab81d032b66abe5f61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd054fa67dcf48ec6c2b8acfe99a01dad735dfb47ff039bd01cff6e413975b2e43b28bdc04bbc6d33c340b2b214f14e1ac10edcb331419d2b14d29938d34875f3453a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1694edc339315a2f0e684ce9d04bfe54bc2faf9170c3b9348a23271fca533e0b6b6dca51fb8b1c05d8ac8647093907da109e3b2929c7cc77916d58f864c4b5520a66f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf05e2b33c68a6c24b1d0a8cfa0a5dcc709cc810c2f17037f3a2f9a31e6b477bc7a1258c1ab4f47bb81b6c918f54c13df6eedc4b377c76c38f06f05ed76bbfed55f7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12bc0a8f09ddc7c6d783b593888266df225182d1436d9bbfa0c6bc15b78fdcbbb651790b83ebfac65e866ee164ca51d9429be0987eff3234bfed3b72d512247733003;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7bad5a3874efeaf6d3c31899aeda38d56961981e7132ed0c78c6ade041bc21769770eb26348e3a266cbc6643c06c3265e3589ea916e5b1578a71543eb95cd27887fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h63dd34b013c1eb58fbe4eaff343b05317a48f8f662d3c9fda6c09f5160b6268e5839cde98f5e81eb4e82685b6bb1875e6c4d0deb8a3e3989836fabf48e86d17aa626;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf396f0a3f6b5e2967d5942c3278900ff1b248f53a292ae2db02f70910fbbc4439249f1d33abdf22251e873854e2c44d39ca677d63031507ca4efe7024743af00cb1a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc28f0d85ebfdb9ebd9202a63a4d9b34943e8c5d75943740778a42bce010072e8240876686f484dff7a02e4be5ebb86ae360f2321e6cec76d805ad0d769e85c6a3c92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b33e9d6a3c8052b6b7e63d82f250c1e0673c113f952acbd0073c5336b263466928390112b431e6c2f89a61be9761798ef5866df6fc9c0329dc36104c83b9e9225bdf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h845656b3f57470d1c856d60672b77f7c48a99141f15573a5e31d7cf3302d49ad7c4198326bd1c2ece40b8731684e740d0ac5418f028109af502f54f6b3e39e1ec999;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c618c3c64888d4e7903f027cfc57fc08ac7a564280f1e4f40e18adcc4c0bb7d6de83cafe98026d10f1b3340d5a9ab5b8ac240835b1e5a40e6c64e2887ad2f903e3fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf0048b61c4293febc91aa508871fac3460f0bb56d9d1159e207899d0672b29fb7af609519c1b6471a1116465eabf949d748c891732175e3b0e07a252a9ea2abfdfc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcee265ccdf898839c069838002f11e172d410e7d18aeb7a0956a76612117c5352dc531cc84777119acf1c1d630773fb8ca1014691ace305e03b7ca7ba21bd5468732;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1de4428abe472690f2dede366dce44b47d56a6f5c4ea766369eef1c9d0246d051423eebaa450aebb8f01c617cd10173cc13755c22295862c4279583a961edcd1ed2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h196d6f239cd729f9bf0e3dfbe3206c57d662b3df50e2d911b50fd516626d94b23fba15e0fac77b11b826433a5f3f4a035339e7a08c8f7c896f2799853a30867d9fe2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he9f463b2a2f6236dcf0647f62dbbdb7adf8d8af8d0c931da40b89a77e6fd48caee1d15d63dfab40097836ae1ea84af122a6f824fce5eb00223392c036a15e523bf80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c77bfb72a20fd9ceff382c95f34193bec0e41287c9ffc26fd666d07d970ec256c22cab7a1fd7c52406f49840616625ddb5e1f0afa53afe82bdacd407999cf68475e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h365d83d53e38bfb8c4e8c770c136ff99da0d7872068fdf2f6328f115e252a8838cb384182aeffa9c00f487bd030dc3f8ad16e0d674209335ed48438c095270026c8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3bbc31837616588810aac2ef78ff68e368206fff498208b70a715630ce971c4391bf5489dc58ba4bb5ae91557910a242d583ce85c7149db92e59ba75c061496a113e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h99f9528bbbae59218db34f83f9c4fae3b670d7e4f7520998bd93aacd48b6dfabaecbee54fac4cf27a0af2a9672912e4f99a6c784dfdd08012138415471c9244917cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h26e048347d109c047917c43a1592d233eb175a2a9014683941e05a64f61b71fad1f142d451324eef2f23e605de23161ed9ef84011854670b36d8732f9e77bceb1d57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13bceb430f73b0edd24877dfb5ba96fba01c5e3e685c6b85fe28809b89407d5434658161b38efd9d1a40e76de2dc0cbf50cc17e6053926d6890d8ff6b5928b374e74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1336db12443d381223d6ec72e37d24942e7e3ecb69828d2207bae10dc62d50eaff96afc11d8c6b8f6aee43b897b347dd4f20a1819304021fd247a77b55e696a3524e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa8787ede45e4b39b7c193c9eaf8e1cec9fc0f1daf0a196ebdbd77e4d03525b8048f1d7de4be873b3921655273125e4caca6e8df902a0e8ebc5b8d0e8d1ad1a0fa6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a41efe4bdf2d7599ca2a802593b4b1e02dadf84287b8312baebf595441876489e298fd135d583329f1d26163e807c73cfe41206d42cb50140dbe87a39fc3e9ed31c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h61d97bbbc0889c9bbebdac43dcbebb71e133c93e78ec06f55ecfef0af87d0f917a0c02a5e5cdc82b777852bffa42d618484d476361b60f06be59efe43370b2e6f412;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3a79f761bca7fa7ae60edb886aa0bade6de0404586e91d20e6e4cc5f6ecc5e101508ca674f3365aa7e4d0138746bce4ea2e27dc82d0ee24a35331d2dc4842e22cfa2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f7ffc2505abc1c3d2b9e30e010afe6d1817f8ddfd4550539c4515472e36a6c0d8b1b4738cbfcd79a2ce4e8ff06768a958f2fcdd0498114ac79e4a16c75dba8a554b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h79832cc9d6df2bd91a6e74182da57cc3e45dff3b74f6660cb489fc80ec20fd12d644e482ecc4f12ec6fa36d78ed1ae8fde233363d5b1f39c53c90d9bd59962c01f9c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ff5844840fe6b4d771e1962eb5bc8d07fa0f9c5046925b8dc96315c1c437ae02b6395f124457f4e52d106b878808fc1dfd4b715ff16af226dd2bfa446d1b6eb502f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h21356f337de6d5b51dc3b7b81b5bba38caab3eaf352bb26c098306747d7e84ba93c0a6ca1c1de7513509c3d27ac1d80fd727b3d82301d4c3b53fdc2cfa45e1cf714c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h92b3fa2159ad279316e5fefcbc5aec58136f4cd207ea6cbe5dad8c1c1aea8c8fe8c0f6a7330ff79d48c7838869f57dacb799326673bc41544e8178aec7231c2d5fce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb822bce3749ead09b7f7d097967bad9adab3737127b2f16c0ef9e1848dd19c48d8f6d30b92e69588f4a55bb37601189981886d4505ae1aa268cad9eda4e9b55f1dd6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea7d53528930ff15ebdc3f19d7432802eb539a30b722513926d367767d564d6d7dc9c15db194453b6f287b8c6ccd13b22695d27a6a5bbbfc59dfb7f82458379fe18d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5a7b1992fcc95d7077a29a22c1162c19d55bcbefd21f0756ffdaee50aeeea54b6cf680f7127ce2ff0fb81656cc187c185a5dc8c8a9da79983da146c805bd5e370d24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h138f749f122c1b561125b3794a8cada5959f6c52e8aaa4e0696c5428d7d0e8e0326bd8f4672e18c90a44ddbb8d9342fedfab074e6eca3f07c32822e6feb520071fcf5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h74e7ecf09cd0484424a4bd450dbf78bb60a752cb84c65e961b73363e68c0dd0bfc2a675cdf48a078efe90b78eab9a46f98c28bda9a1abbd7bc90223ef842f4dd9784;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h70b90c234789da03f90484f4eb458a8a8192290905fa99138303365841a7ba60bf3898d256a1c60f7f46a6fb632b2456ba47d7e17a3834d2a9d606dc9d841a847d7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e53634029429e50002c80d566f7097f22297285b30b0dbbeb9e7b18b9c43bc5b4a927e80703da576df7310af27795f63f053d172393f34530fe9a68aad63629665db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15705e051df2e184759cdd1432abfef1cf297707fed17049f92765021e2d552b4ec15fe9a30025785774aff3da3e5f303951492dd688394045bb5cc827dafa3005dcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b7800787cfe5ecae7dfe8968d1eb158412202d759620a3dd4586c73a3895a78d953a358546d44b5a5ec4b7702f340079983102b9aed0513bd08608e7d07dd335dfe5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c403ee2420e87c1c7bb8c29687299089bc3585a541e03a3276655da76c7af1169fdfb4ac0bd35f7aec6ede44de631cef8f97339639764404bbbdd927f4c4f49a2461;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h12cc2e3978b7e8246af0f3f3c3cf46cf489dfd176887961380ee7bdfdae1eb08df7e96595bf476798acabfdce37e969ac2b892888e56e6dcaa25da359166cf2f5a007;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c2bcfcd22314498f17bd72113669cfe6c314c6f3d9e1c2aaa25f0c8b52c61506d24e1eeb9ee24c18ab1eb400ee9692591ae68672eebceceaef5fe8606e9e94e00d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbf2bb6e34eb06b8c95aac2af63606b5b2af4a62ffd79b6d2e405c7a2f7df8fadd78069a80d22467c5762e935e969101d6d84fcbee039deaf5461fcef1ad1b838beeb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h805923f3fa52bd4e651f90854ba1683119328bee6bbb75412084ff51baa0c737096458a050ac33d6f751371d2f59a6e0426edd8a5ebee34f8b601dafcdeccff6cc4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d22c7b1c6b1a29fcdf926cf43ea70df56f6aa5a04962d5b3f974ac6d27bc58390d4b2fea6a57331f7653c53e1a5a30c97f1c30309e941f391a3d8a751f629697535;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb80961d949f4da0feba6e9f43d2ba0011a87638bec44be37e6210df69d20e65b807622bfca11b70a7d72373c6e546af293c55d1c92b693ae6db3fc40cf986b0fa2a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc36824be8ee2051b3ad913d97908dff76c7a18c49565cfda291c9ff096fa4b27a488b6db785daa4707c7a2ed763bd9376bdc59ef06200560f78b557369061a8bca62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15f6453dbb11436714f8bfcd7ed04613d9c90f627ce8415fbe62c3a3c3bf94d5a029401c2984f3c4d855550e446ffab63f20c0920beb4641535edeb6d4e105cd811be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3d32df0754c589a7eaccd9797c9164b363d729b8698436152eec0c964eb986b22e224a8218ac95f20f6c3ae4c2d2d763a82889173048e095c3b6ef03ab861f9e384;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b2a79840c7f7ea7fcc7467f4574b53bb6ea297fa79ac9582c013e2bd7eea3c8c75c0c98ffac8a1b7530413a4b6f8b7a453b6229b98f4ebcb69406ecb006ff5605ca0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9b81e56515e7da0136427db4887c13d7c404492a9635dbd7f2e672792ae3276a42bfda7cda593840a70e9140f624552ee527a50761182e035f39e2252c2edfe9c77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2bb38839d9c8c049f0fd49af01703abe16bc997fab0a74db56b8c3c4f3372b7f86ec900ca5d5292a95df6d5fc2cbf6aa3a80b11e89d6196a4c676571a85e1143f245;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he8a2676558ef23224a1b0bd6d677e4f6ddffa3acbe01277ceabfc1b657336ec893be57d676ddcc459ead258799a0f375f87847489a398c123eb9d7a839c0f98d8eb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17810fe1517e098ef1b339eb0f58023abb585bc5f5fd5124268d8923ec573c7bc75a8553b408457f09a20ef3d4aa6087ed6b2dab633093ad6d00629f09af7c148d9d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d588e62f0ba9fbce680f787e0bd75872108d66c3176dac593aaffaedae05bc9db1eb1b7e4e113b9b67d2b6adaacb4acda53d469c0341766f1a3590134872d662e113;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c1c2f67fa8021231c9fff2ef05a328bd5537bce6fdcd30e8ca93d89a0f7e9e49cef65f43dc85a01620d6c4ace1ac966129dbb3c0d41bf1d58a59481ce0e0546a7c0d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h906d3955e926837876154844b749ee4719a7ec8f406fcb4ef16e580e553c62d6c57d10aa1c50f9233c9a4b3225510b61a294471d74ce2cc40dec86a4326adf31a664;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf37ba73c621a340cc768ff6bfada698ab03fe63d5d11ffb58d2348a70bc3f81cdb510b828e8588f2f5f2712629941617998e50bed4821b19058a1db1bebd0585e85b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc5b821ab840a02a91a21adc2003b03536e934417f616c481bc202fd2fbdb789682c84976a47989681929f565d616d92c9b74e4fafdfa6a880a7cbc2ccde1628b7c2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1cf9dacf8d17f55c48f2e48635963c36e038c3ff9a156a4d64afac98baf0a21329eb688d25e69f29dc9082d3a91e4b0542680e72f67ddb652f76c1fbbc21df22ac7e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2cf7f1870c153878cc794842aaa83bc8827d1d4483157e1575bf496e664588a1035a1f6c6ffae4ae22903ee6d0c6a34d8256096f89229c41fe16dba5fb21568f32f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7df4e70f49c2ee4d553eedd4fc0bb3572223248bcf6c2e292b54efddecd0be7977e482514a9464ed133bf279f8324fae075749af88e51fa0aa7b2113e3948f282f89;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3f38e9bfde5d8bc227b980f9d47f0cf0afc3379a3bce8029686bb4597ade68f9d498e815e0f92013d8b8a4d9354d3a179b6c0047dacf1c377de83e9e15e17d8cb10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151244f49832c3683d1348d645f8823cb69fe2d6261903968931ae1f669c4e33c13149e1d09841db2af02eece7252a41c03b18ff2210c27408eaf2ad0856d48c671f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he704b4791f3c4c8efabd5328647b1ab13a2f823b334e41cb685fa6f997e56b779345ad1cb761db1ef5bbaac713eed82810022ebfe4f30b474d8ace6a4a94ecfa1352;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he433db318ba7f9dc8d438147fce8b4eac0304460b3d0ec49e94a4af14830ff43806266de71be5082127d83f6569ad4aa841aca454e95900b53fa3b95f459becbbe7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h456cdd1ecc43d4d86654c2a0de1ea4382e465a4147702dac3b85a3c18a9cef2ad7ce06b11bcdb5fbaf7977264d644568ac12c8b6eb8f87d8f1c9d609432ff4d0e1b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19251021b5be96b263b2b497ca159669771c8359a60e47baaa9086297f808dcf10c422f9796f2760ba5acad110d76d5ae9e8de95157287f9f400f4f4e348307b5074a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdc6d0decd507eccaab9ca7b77042a663125cf4c4cc7fd20b3dc665e56a8b007e02974ae7d1ca21305da08f3b72974720e9afc9b9fe8d9e075a6f0d253aaa0c014bc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c7828c1e1ce2194c604c1dbf4223ef3d920a8b8dc0397173b21e634fb0a73f6da8bd90d92f9a813a2109afce4ec1dc93296fe407566f7c6d672c92520f9879bae78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2eed5a9aefdbfd7df2b9eab4f7d383747e3ed2a69b8b2925769429602c9ba475c49c7d643d69a71486ce7c3f657ac382bc9f78d26a4f7937c34e2428702af641ebb0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13f80dfd26bac759849fd9c6498737c2c71d552df5d1d7ecd039650bedce18db1ca54264b478eace77b43545f96f08298b244b0c6ee68a010ce24bc0ca85b49d3b8a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h126e0594122e6a3b99b4dddef4f857b631ae0ffeb25ee064e3867951f9f374847cc855915c9f2ac9c646e641c69c261ac569b76eaf1103ffcbd95d2372d362f033b46;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1524e7257f130fb356c034f962f0cbcd319c7d52162c82cee74b6365ee3f8c2fa279832934382ee31ffa554bf649b4a02d42a0d79a4498bdbeb6baa4252aaa1f163fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbecd296ba17ebafba264b923dea08f0ccfb608251429fde88f5dab64fe3618a85802aca2d853b620017622a6f09b297835143dde085df6ef952ee1351a197b3c516;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f7cd4f290fcaae70a198f99ecc42e3de2194b9f1414325e4552f81fcae906afdb444c78b586176250fdeb1726f4d176c6fe2a5c403bd238837bdc710e8651ca8af5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1998bd6dc02563641d6cf828e075b8606faa88a3dcd3674269d2ebd72c9b1b1f5f9e22d16e3df0623533201cbc45bf6ecb589a0c6b957806a7f96a15c9bbc4a2e9117;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h181451ae11ba093a779938ba9a23437c1b54207fa9c0b9b4b6c6227a92071daaaff95e508b012621e8cd94539c9af267d680274f519fd067467689c7aadc797423ea7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd70558150f282f92af90a43e9dc9c31419dadfccab5f4920075a04086310b86f4594dfb950f6ece6596c90a67be5506370a1603bdea2ac7febd724702f8751a25cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fbdbd89a0ea87be5dc300f24ce879b174bcaf32f6453a1a4d4c0df3a48cc5696906a388cc72f08b487a741b443c373f192c63ccdb3c96c1f02017bc43a65d8d73f58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h193ef485d636054b7590d8f1c0657a144f0e79f5887ef086ab15f4a21d981a0bfeee3db76bc86bac899ccd7e673e4052cb3b37c7f0f6b1c810063779e1bf9badb3c69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1afe8fbcb2588a83416c25248e2983f43d819206d47541aa617b31d6ef499cc6e045d387c35ab5bd6a17fc51642c60499219a5b4570067999d602b2a3907f630e68d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4bbf7a662c1982c01369a5f18be0a9f85ba4a12eebdb0fe97b3d74588aa35737dc30a1b83d53c7880569d277f858ea1beab2fb2db71d8f4ba6970e99fc9f15deed7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f823a84274072c1a3ff4b5667e958140cfbcb0a512b5dc83888c7b6bebf740db3043152b85005ab1e1362e2db5057b44e7a0c52a3039129a14141954eacccfd896d1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hefef350bd374feb0d74bc3c3e615794d5f45aac65bf29281685881e0fcba730530a660e9db37e494de8e89d518f638f479dee69556bb838e5fd466f7b8a20d6fe9e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6b28611a1118a710308ebf3af83ffa5d98e10f8f5951c11b67507fbde581d61e9f09ed0c651198926fb5eee0767334a25930e99692cbce99ca683524c3c78906963;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a6467b50d9d31633049b87fe7d90494eb1871d264ae0d7483c67747d643ce469b360018ee83b55a6da07c08dae36d3553abf34383190890e93d3a2eb24d813ce242a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h178360998b2b853ca1f7f7fc358cdd6ded3551f89d9077a3757a1005dbb7cb6eed938811e1b0ca98adce6ab3cbe8f81353da740f48576b5c30d9a85524ff2594fd8e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14a4ca93d157fabddcb2263d0eef869a58dd3bec7b77d7f42739252c1d8d9f23a226e2e489ad3077ad2c61884232dd05b6aea6d8ceae873e16e70cddf41e2738ba4c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d3d76f0e7c7ab2435c99c25f55317a9e0c2ed59aa9a4f8c2a23c3893569592bbabe8301b709477158bfa25faa8c4a6a51fe5bd4b6209c160a60a9faa62f8d75759e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13d235e19d38e888a5f251deb35857b8aecdc1582bbcd19abdaea1421f82d80b7c939b80550a696a72777c31e358a66dd185f43715e08db4206ad419a6b0918608a95;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h89a0a7533eb81287b7afa40884a9e5f2466935331c151f6095c0a84cf88cfa02168304359d36a4ea0a7c6b8c34b4e715642df37aec1737677c8db33e879564db9459;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f746f6a98d5eec1aa81db7d6a4b5e6c2d7625470c05de9a5054923d0a2f6b1a478f26fdcd7db22ca5e3b47f7945be7bdd8d88be2e77f5de91b449f83216177ceb1fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17c92e6bef936565f6fcc9e96981c15467905374a1f57660e5ac757f092654a1bc7f0d2211507266626bae21942df44817ebb9e49662533e5f42f2dc0a669e67be4a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc0a718769323ac6878cac4ef5b1eaa1e88516b4c183b1e0a03edb787d72c98699b3910883c8586644d2fb2a2e75f318863d383ccc290a1860ca4f2fc1f5af4ad504b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6d1e1c290c6f3272a78a2f3edcafae93d06cca6a6e6d066fa68082e18adf44deed81ab879c36656f3c56522e0765f441ef9aa27e3bc5b6b881536eb1ad3e23ff4d43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h996544edd22b837dddcf70d87cf22842d12412a8b76ddb8645d2b97dfed8708e283958f90df52bcfbcd0ea5201029e2aa052e438e9bad011f10530482d250a705f64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18bc86f9cae59c00edc849b869700387341f08e48e86f4828c77b2f6296ca836b29d2ad84455efd3dbecbc8f8381bc07fa8a55e81ccaf64213aaff9943fccf6212fc5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ebd96bfcfc81c62e24277514ced1da9f66f0119ee828878b9682cf7294b740580ede52e91b2b4c8e507903bebafb4318bb7de00421776a816c1c239fe66f9f4b7761;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1485066bc50b01b4106152c0c6a1f42eed301a683a7d32aceb808cec92708e007eed14540b91d2960c8bce78a2f4ccac469d0a9f09013cd610199ef6ce15db608079e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9cdb77da342ed85f8e6fe47c4bba8ec144e3cfbf80f6ffbb4b91b18d2aa17a88c3c4e6f51c5e85588ec91de4721068c4642c637ed38572546adf2d037366b2bd8b51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17d28dc7a1ff6beee7acaec8e90e153384f28d62b4d86632e1da9be1d724a624fccdee1d864b315414e5d354c44a7cea41041ba7cee99f21ffbd86f6369ab95c76d9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16c8531760e3b5236fe27d132973365ec28b0e401fea5d735cb195166cf3b17cf68085be6c0f2b6a951e3f3c0c1d7f63b71fbb007e1eae4f591cfdfdfdd7e8b17550c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf8d6889b90bdcbfb07cb19ea186d8b26aba56aadbac48b333e2c1bdb9f01e19c0d93d4cddcdc1a6146f13a688842cdc4ce40d7bb7f134b0fea3c4b82eaa87f02e41b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d95f40027fa3cd1e37c0708c443d28c16ed477bacfb570d1826d37a4c7e3d518c8d7507a1ec2f6808c7ea0fe350a28b3f01237c6cf0cf9e5518b48d5efc0fe47c56;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e527ad8a7f814ffedacadca728c273757ce2cf99a0797e00607569a1e7a15533057e7bda2e5e91cbe5ad752d2451260907cb673b47824e298f38b8244d0f48b592e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4469f4d8a52b5075c11813768c0d2d89d281bb5cac6aab5a4862c9263835b976f64fb26735dcd075da66119f7e774f99e0d9044e4bf7e5e9fc153fdc830b9a2f43c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h18a98af571ecc22e6d4e13180dd33892df38faffff28bf60704ac36bfdbaaebb97cd568d36dc1a6932dfc95bd7144dddbbce28d59c923509dedfb0f62f1b16cb05cff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ab34fce1e65cd7df3c95f5ff93f3447a53c83c9b7ebaeab50cb2af07a6d9f7d7172b6a1aea4c18a0919507a6359bd927202a6768c8c615d60ac53a1bd8e31a37220;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h144cbf516efb982ec23113cee7e9e4a945e72d5c5439f7c7a67123b71a6974d9e5bf8d6844f3bfc1239727ada848f49fcdce44cabd0e0c987532fc7a301822657ceec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a8c9509c19c6e74cfa8cddbb2bafcb5f4bcfb883054ae2992bf9560d0d819f699dc893eb8bb5319b8c2141d0ebf997a2ad6b20927b6f09536e994ec419210f30e0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1612725bf16031dbd874e196d617a33bab06ab0a4928605ea4dfba3734c8c74715be76140ff922c207d8117c3f560661989f8f7ec78b9011c12382524aede82ff4aca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha75e1805a63014e72908c7a05291239463a2a1f03744d853e141fd930541ce694c7dd599b8f8adb16ebf4054ecf34112c4b7388efbdcea243bef376bb0c00586612f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19854f525fb485152c61561d545e713f3f9b61de66b4852b20b279bf54582284b3ca5894d0da869c7b321be4533d3bf5b6827f9329cd9c886c3b29c0a4e3b1ec25e9a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heb1808425e7b58ba80a451acd92adf39069b236c0baefc35a41a2f73c149a361f1bcd7d01705502538d4af895bf6261ac20da981bd7fd54b7cdc7c5054e9315b7a6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10c4866966121da35ac4dda47316b077d2ef5bb27b90264da12d9779d33cf877ac3d04295dcdac07340485582fa3cbb7212a4e20284289b68e9877b112009b26541ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9fde87a459fa60e8856862572c3fe622dcd4d6c389dabfd544b59f1ab7e2642e4cb817c0b70f85a89c26a2c6b1c26599992cfbc55bf3444682cee0116babbb2e4a2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7074fc0f1b1587c7302c6494eb503032c38ca8de4ce5677c4e153c3fd6f6cedb12bf0a1746f7222e526b10e3dfdd30e1a096da6e63aff2c850d1e0664aafd0aeb534;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf6c40dba3f41edaf24fded0cfccb3cbbccd7b21524f32791d935cd0ee6bf44794e00b1b15e3f51b6f69b5e177dc0d292174cae077c0bbd6ae13cd8ae19fcaec3419;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e6d6a4c2012ff272f270b9b8a8d5843600287f074b98f0414c1a3765f81aaee5cce54745601000064574307b905416ebc9ad96c0fbd3dbda944415c518281fcc2fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf29bbb67d6dca505748a45f603365db24b381976f1bb87f807a7c52b5efd63cf70b9ec6d23f93c66aad6a57ba9a5d710dceca5d57bb4925360062036cc39d79a585d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h555fc524627a6dd318384f3a418ae724ccb3323fdd83f38822bd506c4efeb79239bfcfa38123d95add06760c891b5eb01bc79513c234ddcc80dcb8e898b512b0e6f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he435aa50aa2560cc6b75eae44c29a1cda49379da63a277f23568b91e1bc6545befaedf6e75f5267d5d19425c0d7ba12daad10a070d6b6027f1359e31eb53b2be78b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ff85039dd7731b2e182a8da85d30650d0374beda48bb369c3cbc4008b79526a8546aae184aecf3c54075bb4e7ddc2903238b8abef76be0a7a9c0be053ee0877a6cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3c901c6e9c89c87a8585c5aef9f4d97da5cb0423f28549de6d3be3c37d36ef99313eaa789a59075063af1bc994f278a60b088f0fdf46e8b80a085b5445f09afeeee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13626cb8185cb9e703967f206ac7603b70a0891ec4dcafd13c4785eaf962231ccafa611230858d144b50effe21020d81ad2ab815128dd8fe74cf55e5648bf920c9331;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7e6036af93d0c7fcb68bd0c86fd1cea47d0e725d92be31dbb0d7c6407a199c2554e4996b9f7fbb9b89895c845bd5d50901484dfd8f45bfb379175211863bba671838;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c1198a6ebe4cb486c50cdb58b328842dfa511a7feffa26161170eeaafb74a962c1bfa0d339780920134a4dbe954bcd4e0624b4e1d369794f71a20084de31f3dc4a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8854c59703d05a3e009a70ff392ebd3d0a5597fdc09d7253ce3a763a5de51b0c3a8890b1d1e119dd4447438ef3ec9cf69a8a1791470e37438f8603e195d5cb1651aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heea6be7b9ca0c143cf338a723c94316ee0a83297b7f6e961943cee11483a5b02f2da015310a768a8a4432b647ef143b8e665028ba889b3be8e119a95b32cab4de4b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h220cf395f3012d76e8df69417b7f626cc6a64dcdf4a12fc926e8fc7c730fe1f8e13a50ddd529be357bc257a9b5e086b791a8c8765448868b208e97da53b7007cb780;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcfb570f2eb0c8956a6bf4f7846fd701f0755adf8250196fce0e086922ad27e964db0ffe8bb00d24afc62568bf26aea4059fdfe457bab7be8d71f33af21c83c6b4056;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f0084d00a88557071d2a3bb2a7c77d8cc0b2732b336953de6a311cd08d0719b209f7280287bf556c8ddf4af95ce47f52cc353432bb5355bfd1d57fad907ca871d47b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h702d685bd3f592603b9c9a08ba331a21d336c917d692d196f066ef4f8c87c3cc61d0ac707ce32f236ef8353344bbacca1d0207da6688e843d4419bffb029f7f7e5b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h157cef073c305f5f7445c53550cb742337cf393c453b696da7c1fc5bad2aab9852dfa7ef72de4fb7c04714c4f68fb9a67796029aaa225ca373aef758592e8f70005d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14ddfda13994d862a8e985aabf725c05ac09e55c6ba313f2b17ffac3b3117f0fa8e6c75a17e6622cf20b304bcd95aecb90d6479aae5938add93edc5462df51cdfd36b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b9c92c2154e2ab02467746e772de173edd618c8916a6069c77ce267655fa8d6ab136cde3c71bfc6367d53a22a1eab5a5c5328855b883d28fda6fe9b168262d22a56b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h13a90e91a3474cf19ff1efa94c4d175af025b324a02d88d5cc2306efa01c4051060daf10bafc058399ee78edd3f1a68a7b56c8f7856630423179e320b80f5461db753;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11f91e0a7757f4accf09cd7d19f92b546454277f35f7ffd0f259f7787052540702c2b1c193ac1965d00fe8778cea24c2f0e745490ce604d6a514ca10a27ba3136ebfd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h110f10d581195986d902e562f48dd204e8aff0ba89feb5a5250d842192198a59f9c6f1dd397b5956336722ddee714668a3442f7477855d23cac2b4bd83a964f407cc4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5ae6c97a29114896a7590e45e34a3bb176795c0ff930e14cd0b97f27cb28310948a69a3570b5400756a7818ff1bdfda0c04a09e8d5e1458c1389fe280ea21d9573c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1711936cb5d75b5d6467fc3ad333b41c1a51fb787fddd5065a7e9863909372f26822cf214464c6a8806c87a14d7aad450025da820544cbadb97eb95cc3c4a0bc9356b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h62d83fd12753936fb1d825f71dccf51c22e30b2acdc1730107f6be73bd0f05c334889c109055fd6de001b91ea924386aa0b3d7098e44c0280ed8c8fa114a7e1e15c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ef8ea2ad0aaedfa0ce5c620089a321a2b8944403605ddcc8819b47817e62b0109ba3f25625318c1a0acbf7ce4b0ef70f915b9246beabb624699a93b0a4ba6e27bb2b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b1f1b2be2d7608f9146e55f56d11722fa6a3753eae46af7e28ee316585586ffdefc4b0ca2a95d29682b0ec13a2681234f6ff30618a3547449ff3ae3a18206d4ca435;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1eda1c9aa40ca6dcf11fb50e6839c4bd79ab4c903bf33fa2444249e216ee1aaff391421c9e00d131be771231fda1a451dfff94483b6b5287c62ed96bffde544bee380;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5cb964cc2ac718e5841693d6f5b15a7dc9bb177ac7064ca1b2e6dbfc281e76d3f567355dc8a2acbeb56ec27a51e7c4f024322040b30b834ec7e62357093b9531ef5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1314967838e80bb264fe6e6d4dd91cf5647c074458c18ceb958417a9cb02ab7937c86c1d33a548cc314755cb0af582c757d1e55837d88cb328ecbe260a999c82c4187;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5d4b40c6482f24865bbc30313698c3be91e74aab69a1095e2d15ccf463aafc9fcb1fd46caa0d524c9b48fb10b472f57ffa100f4b333b010343c1d61b239f58823884;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16110543bd0f31fc03a500bf23a92ce94963523c6d44ee3673b3d7909eb41e8ce0578791aa9830fc0824e31525baba76b3dc58c73ba7f3b2aea2764f93bba5b6f899c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ca9d0393683c43370896c5132ac33ba0d36b45f34911d6d2b0047a6c6ce41318ebef109039dc97d7a956658138bb5ba8487ea32d757da1ee0ce56a9ea30291abe8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11d8723d7e680c2511df3d2f38ca109862c676e3deb8b25edfd66ae4f5e3507b773097fb0a39559d4c73c5a81dd8e746cde008db951d51146f5c880095e31bc6c90be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fb20bda66fd7230a817294c618033ee173bec9847c2161ad1882d1d229c4d0e2ca7af13fac3307ddc5fe364983f46c6237c9892a13738324484d6533d1ab55c8065b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10da6cd806a3997d24099094429132a545637f71b8c200ab8fe6484c77fd1fcfcc5eff5773180627d1cfd123a773d721d36e3ed7d9efadb504f7c2c135be726b5d644;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8c9a34d48c6f5cf97680421419f99a85583d2203b6cbe878f527d8f7097bcbe5480ae2fcc7d219be72d732b8ce3abbf43c47c8caa7f1c7fc433cbde65c80880189cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175f47be4570656cf7e8d9e6138b57c040d0e52ae0a407c0756c0dc4bf527126b2a71f1c485a2b45696baf41ee2ef8387dbc627333c6bb3a672085925c2eebbfd65d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4daa8c5ab6a000d0186e92869e08aa1a2675aabc64591c961705af38e038b625fe28bbdf78ecd6d17a9ba911e5ffdbb33e7ee90bfeeb3378c1d2a803b2c5aca868ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc91648a8945b38817c169b55c96ac4ddddfe04e102d1ff3f0cef5a79435d5d2f97187df63b71dec5820ade570d3e0baeb90a73652c23cdaaf49323a532aab0ce751a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ad5d037b600c1331f6d03365e697d676e2d052beafda573ecf4321c3a92869dd4116ed7e50d4c9bd38532d287cb001679c57bd81409b7d7e0f6898ad3747d7cbbfd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14514c90dddc5056029c65cb5c1dc53f12c9e727ad084aa52fc442a60664d431e53261011eb706fe60a68400e225c336241ade3942aca8d2eed2c816133c5b5958be6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h584110c0c5f05f8d004d59c1121f2fd3faaa97ae75d7a7824ec7eaa06ef898814765be863c0576ae04bfe48f7b6eb484939ca52652e01116fd2903ec609851e54fc7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hf3ed2ef7ee4c216c8e9e5968bee6b8381e1d9f525946830d2441dc3c0c7567eff04de41286b7b4ac565791e4b6096b03521e00e7c3f86610c3f74633cd21529fd7ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10636c773eb2214f6d2e858386e096ddaa996a6b254d5177ab804d8c2d11ab22110a7ba195c0241178a7a40943d789742dd57d0bdebc9fa9c4fa3f332ae32493427a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1035e2c463849cd3d736464770e60d1d1670e06e79c54296fc67c36ee37c30d14ea704d0f225751f7a85ccc98dd3cce86bab3882b57f971dce0e9e6d5c26cf3b0b04a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1987ea368b4fbdd15621b8eb38793bd16614167165c70f47f576ed592b590e7612656ab0910942c95a7bacfed6b29a4c5a88ae918f8cdbb96a344528e28674b9c5b0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h6ff458e473984d6d3feed467b3096b1a76ac40ce94d9f24aa5a880069244aeb591fc2ccfaa78d2f8bd54fd65da57265cc82e801d8e515cd943a642058ec19b88fc79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he45b4fb3c3f42ec7d42df96a7f5d2cb4001ac0a90cc4fa477fca55b1ca3a8e0b365fd31819c5c0c9491ab9dd12a2a2161adcd121072381965b5ba22ff5f6fc01f7f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1da4f5f58a98717017734d50cc65a9bee0c7584436eb0fdd54fa6341c0a77dc8f6effc79ff100d917bc2df16c0952800934bf5dca21dc4a73c29540a59a09dcf34f6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e5ed58f1dd73467b058dfb23297f8736bd92daf03d298bf5dcbe05fb389c1f6c4755f9ede9258625a5197412330a2e1e943fab19f3b7c072fd5b92083852a3f8b0d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ea234595e2978ff1def30a186807df49544f3b4cfc7cd5a3a3e90b7b2d123722d95eace8aa5da840e465c2c7ef265521820801480ef424f823b9d84ccef1cc717085;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5512f56fa414ceb214e2a1cef590aac1ac6a2af18f3ffdf5c66ce56829b80430640004703ddcd9d64dfb1cbd003716d52d23f13601b07372251fa52b7b751fed6e7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfcf4e0d1274089f42cf0268a2870e77efbc1616e0b687bba64498f4e1393decb4f615c3d2334122dfee6cbc4028a1f6f0695fac785424a85517ff7702d6591f443d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h600b882538bca0e64cbe2912c9b7b10a0e0991de29ab35935275cecc9f878702ea044b6cc43a7341ce27c0c434bdd727507831be38a16a653d19b039cfa973728328;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9f769ee4dc034d686d376720f92c98e6034bdb99383db77defa5f412e2f774c673286c1492a28049154c66fb3d6cf532943d8ed98e0ac4fbc50ae4fdda31d4e8d268;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h17692fa29803f1adae6e57a4a393306938dc555102e5c35ec7ab2e1dc7745b62a044b7346f7391b421a4c450f84935050d3edac6c4f3b9561f506b0b8bf52faaa7459;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3a8b01592267056ac6a4086c0bf715de07d29bf994504df005d3128120c47d00c6daff568e8c4f20ac3a2315435cb6e768e2b3f20f4fdf53c61d3531d10f9bfa939;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h891e9170553800db05b8e32226fa401f159a11e981fd70ce30ebe5b073d5e777d6ae910ad7d72cc55d35623d3eed87746f25db51f0d612857bfe1f7e2d8d3f7df608;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcd754b6bae3d64494ac98ceb2e85399fb9a18346a81cd6a20925e0bfb42aeead462c8c0f68e96af499a57a74d0458d2e267cd6b886607c2c00a31d2b3eb0dc5d13f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h419f591cd5c577bc370d21ad6255a928f57a8d211b04e4dd27e9f6348acd256528b50f8afb555f2e743e7ce60c93bd41c3caf0e3082087d13da58627732a0ad32d0b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1447f703a37c53558f41902f8e72df6aaf65c60da30ce264a0ba523bd09fd0dd9efe1453acb2bdff5b0b88c24295af87e6f15e5f5792278a4941caa2540608c544fd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hcb8c2d651d3fc1f678392290389566b62a53372c3167946f3a2490cc6bc43ef0ab5f3b7a8dd6c76d4d0042140c101b349c6eee130627407017c41b80cb2edf56895b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10963a34a93f7aa58d25e39444faa7b82e1155ee506ae560409254e368cd3e51168c578e0980c2cf4484e844121c9069900540b1a4ca04e3d06f2816ac5f7769623e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e6f3c40a7e70f27c1fd9a8c96c0c4e09a0fcb314b51c58754f57470b21f835b3e367bfb664b33d9f2f520af8ebbc9cb35655b9fe96da304efb49e0889dda6e58772d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h81eda71d19998479322569132ab7c7c94a5eedc774795dd0ee581aa1eb3b9f58f1af199afe0cadd15b1c884438ea0ce8b4df2f003d7a913660ba469d1dcde23bf0ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfefccec5ef4312e1f80ac5723f739e968cd062cd2230ad3f4a6e46d9726fea06885e350a434a02608b37fd48e52dbd55c11223b3df4758f704f55c58acbabdaad71f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h44b557fc756bd0607599fda59a35d0c189f52ebc742357cd0484c4a580bedc2e1816e1aca3e5be4f61bcc3339105abf3700302e0251905dfe825275795b404d0d455;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e099c52cffe9470a0167e3bc8071c9daaa50a64927235143cf1e6d44defbff0004b19cbe05b8263530ff1679235b28537c7fa5f934220a0ca2c3405f2b45102862b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1711d157a03ffa56ab9b243c313e67998cf7e4dc2da7e9cba8b9d5d1ec4f6ef87b4ad844ec13da92d6d444ebc1e05acef4cb7876f83692e4993e79709c71f7f9ba4a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h156d00f132c5045640c47881cb72818a7d0e0a22312b009828ca07f5afcea20be9457abba131fa3193160670331d74b33d57e26f9b25a5f41578364730df1f24b80c7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32386aeb6e09f44f361147624e1730edb73f6e7a5fcacc330cb47937ceb5517e427e334239a571511a5111498f54304220026e75cb61951b4b3dd971f8e516bda41f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1261cb3cbb74ad5af465ccdb802fe9e136f4eb7512ee411ae72cee950782639341ddcdc47ae6ca7cf47c401cbae45850ff94654db981966492dcb9990d2eafe56744f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h146ae180e8ed0dae0bc7344565bf68b5da16b9ecaab8c61ca01206ae097ee340dfbec0f48275c3ba822e22f57140d8d9f9ac94473868010b9978e3fe68e39da749fb5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h32fdb4c6f7eb7df788a1c2c2aaea7061ef317474a51046718fc6489c9113316425ace842195223b280b2d599e895712f41eae0205ac4133fe94c995ba35cbf1625ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he3c7d864df674acadc8896ab3e70f045daa5183b8a64c41cbdb035aab02bee0bd708fe505c71cd8e7c4d70f6054da94e3afd544460e1aaf40c2cf08a4aafc5377775;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h174f26bb61333aeab80ade312e62af6dc03c35f88063468c11d45275c204cd247db3e5d8d0a0c3d71a8cb11f0cb30f948a393b44fdc965239f5695b569a925c810f7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108c15c1d64e354ca8a1224be473242921e65fde4bce0155a488d52993f2e5f198fbba7ccdf5e22d1ac9acc97ee5b99019898090f92c99f547f800a6831e7a16f4dac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16ea2f426e8fa3dff302710b9e385a975511072f3fcd587367de2db11a1c2bd737405fcba108669840ae7951127f54e640b1b777d7afa2bb3003b882d200f92ebb42f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a413a2c1475504b2ab12aa739e0193782af6b550901d825b618d4bcb3bbb46bcd1501e1985f91764082cb2b02f1d40a5d46e45adcb31cb113fd223823384ef78bd8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd3d3585b4bc67a9d1ad56d7977798cdc40d23a232c91823bfbf4149e0e7ee653530313e4357ac97b3e0037486218dd5cf6b0ff335bd60b3a6a12907807d58a7bd43b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d3ed60ccaf77ccce8e87f094225d4619c5404fc73cd6ee930733e35cb4dbf0aee6553a99efc634605e28c610b8e520b411b9682fc2101a6e7316183518432b7f2bfb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b20cb3a944fe476f89f7efc4da52a96ca6a6e43f364efb9197972bbe34d9f302dc7a5603aa994dd5175054d9d282f711e680d53d8535593611f12e12662050c6d7ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1bd97e12a5640fb77acc2c7821c5ceb9cd15f10efef9d139c758351a76b75bcd65a9d87b0555b9307398894e935601bb74d720af26b440e270deba5ebcdba019dad86;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h53f7302da476c569c7774b10643f66aa4522efbf6712a25330c877f4ebc8ba90c8d315a372b1f7750d7bc1fd5f79cde4d79e660de75c776d4aae02cd144a3f488faf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h54baf4c1ea014e4f693e0c8c655b83c7b3ec60d104f024cfcc6edaae150b3a083279cf3e05dbe20b489b20f669df5a09f775ba7f20b8f1ef31a4df6640b771e02b11;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15b435793afd29681d3328d21e00e5ddc8fc76e0b430d917babd7f0f55cad51005816d1a802a833dc07431b13d07edcab40c4840b5ccdac1119266003139dc23b7c00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e1853cec84ef4b053a64232f0fdacb19941f91d06dac3855ba9965b7774e841356cc43a16c0e1f3ee8dc76e15bc3cbc00a6443dd88db146b588df650458cd38f0cca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he1eedd14e91565f01f553081c747a3543889fe0a1764984e3bcb61a8e249b50ef24a52c81a5ed0c6df1d8ca164faacdab930a6e0b40a8a402d9edd8e92bf842bcad1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c3481c6fb4dd5daa6037049a671f6668ebf511bebc828ae6d985d7ff2c7d2e9a7fe884c361befa8ca8ca8a65b821f8712776d1f84fb664ecb3f23170721576101371;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'he74286077fc846fa16c523529aae83b0b43c088cb1969a7c6ea0dfb62410d4eca7e236c5b84174cc71ff8186f5c206a33ac6b6f038f2c484963845225b1c4d90776b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfe941b73732bd2372079bf520ec8ff9591b58e13e92ba6bc53d3f36c69a1c9add71283f7f2cbcbebacbec74f151484004e765aff6f6d84bf7540ffac72dd8cd71ca2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10f9910353ea8bc9ca805a1dcc3b635eba40429f661e044390f12daabcae143e4c5c3552dbecfff7a8ad0887dc9e229eeb40d26ac144f4486eba3f1ec7395841af4b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c6909971f3afc17a6b41081c379e124a0131a98dbe76879e42efb1cb806dc4c2a7f51d2413dc02e7c9b20d4e45072ccd6aa815eaff7275b4979167a215304ba2ce81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd7b79a0c9f8369e0498c02cdd3eb5a201ca0227c0b03a1c52ac4a158a1d49dcbf237d9f14c7f5249ba75953d04fd73abbcc507ebc8923a81976020ad9bcf8e71667d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d12d1b05e803a0c82239ff0e07ba1ac095dac414f5f4dc4515d3cbb820ab768c7998348c085789da4a3293b767cf980f378035e6686117849476e3981bfe76614498;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h111083ff278943b2b897e2672a073c6a9b437b109ef8a98940567bb44ffef2f0badf302ed57b802674834c34ec7868b9c8a6d3abc6c7b18845e0555b0c4990da39bbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h49171331b0dc53ae5e2f134d4f02bc159fb0173f66cbd5ec720c10c705ad16d48adc3c8608feaeaf1d135b8043fc56b3b67244d258858a1a5663ce47900d113ffe96;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3c7b8993a0e0764dcc11985e5b34d9e58a40e11c49cd6dd95c9062798047eb3c88fdc892f224463fd5b5f51885a7768ad804ec36375e03e1165b57fcdd0a7f6d7218;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b0c4e170a1054b8219902e6a55f7429a1bcd071d1c6ab2f1ad994340523e5b6b4bca70ddaa739b0d628566d3c2f556ef35c9bf26ec886b312be0dc7527fcf1457aad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10a03f66a7d8a6e84edaacf9462052b289cb1325bb9a0df13475823d5da15364871eb749a6cfaebb0bc8afb8f5e57e3ae8caaeaa94e726ed77cf89be714c14b9c7816;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h19a8a94589bfa293266a97463d95708d65f3b7f40c1c61737fe230411be5e4fecb4dd8035e09bc39755053c7a421779a863c7dcf0d2a4283f3662746cbb31e2b282ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h9666293110aeb402c96eab47c96a3140659ee21af0b5ef43777aea70bcf96ec90a83f21cc0945810376af49ca96991d84348a827cf6a298b451c78a89ef9bced7850;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hdfaec13bfed8470113a553a48cbd5b6fde659bdbb42d2bcb975dad36a50b168112d39cc62b6b1d4e1b119a3ebf33d55ac6e8f17d39b66e7c0af5527ad77f7120a98c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1ff79c4e98e4481f73fdca59cff3c782fc1315a57364367edea30e8516713037b70dcc916b4059fd6b4c7f1b4c9d66d5241dcb19fc6724638491c21413c43f9bb60b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edc9de6a3289618d5d4179f9987926f23f21ad4ce7d64b42d254e0c8d1c282d77e4d5968ec2e0beda814de1c5e3345025e163fbfdafac873676018ae316da446595c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h112b5476458416c00eb91fcb77d4ffb4b8d16620760da0db2453cf30551e18ad138cc7b569247467d9f04a1e8e0a55095390459f3922fb37b5e398225778fa2cc65af;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hd8b31d1ca96311422d18f6dc1fa404068182b964a5de566cce17f84d38b20ffb7fbefa2bb34d84ae27183130a1827986a971f96fca69697fc42ebefdd9a48cee5899;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc66827b030fbcfcf3fe2941d9faa6f0684fd5a1858c346d089a870a6662ef12a0c498c7a23395bb6eaa7dfe9af9024be6b55bc44174aee8e778934a8f6dce89a361f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7eb9062b084a020e2c6fa9c1bc3e3a8b20d81e820f74cf68cf15d72be037aaa683b3fb9474d6241406b15ad49b4bd5efdaee1b7f41c5832298c609d95a6ada442080;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h4e3a1ebec5e84817b0fc9ea1699595303e2b54447823350d3c0136f2016e37fcdff6e02855199236638dbb89fa73dc9a1476e8c0195dfac73fd45391494afa131896;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hced81a6fee53700df6aa6e774bb3aa019e9e00b363e17e62626f0562fc196808891a27053d1d77717b301fd2d80e0dbf9094f7961adbe79351e9df8a48cbbe86a518;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c8523c0deb8d54e179971bcb91f583556c4baf8d33e0a0301feecaedc0340fa6f70b6fe95e40c2ff77a4ce59330a67897f22b4a3e40691e52d95c7ca96461ebc843a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7fab4ed6b4746d8b30180d67dd0648f4ad7e150846542858774c27a8f18c805ba0825879022143870b9e5ed204fdd47f1b11ef83dda39c998664b865169349534e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h3432841b07f3a92248ec6a3aeb5ad14e1bfe9d67667a9729e801aaec8c7984be793d769aa9121e2b7504799854b2f0b1e12f068ae51f2e13eb486ad7bd35e453b3a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h58f378f28dd4357fb6078bd2c2127f6736878b6a11c54aa497faea86afe3a13d389f68193fa2f2d15c1c5800077d7cba65bdbc7ec1cc8c95fae76c4658ec309312a0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hca7c4f92518ce0e7f00434effb01de91111d06bd2224e99405e84587dbfa5143f0ac3ca3b33ef711ca089af7cbaa92b84319ee6574d0b0740a5c0818e9a6268f96a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f31ba5427e35e0bf5768456205cf0c24aec43af5ce2345ab059a17128a51f431c0afd8661dc562c9b15c54ffc5cc67d1a6e6bfe8392798bb55f1e0352e5a20c45905;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1147aff448e6705b32ba81bcb3b927a1b8e5f11cae8abdfa861a34754b252ce09eab332ccbbf6d56df35833413e37e020f8a419037d8a31b8b984d270436f83b91f7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h66845e50414a4d9f2fd9f86e062b433560484c24026142b85784542491aadfc8632819eb68cbf9f9efb220c4891ce905c971770f544f4e558f7032fdcda10c52f117;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h15810222a31dd2d221da59a721484c8bdfd9de5cc4f996e97d6c7235e3e8dccf8d34329ca1e75be1e2d82e2edad81b6a9bc30306334445779f018fe1dd503061369c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f343c688660e49b31c5f6c10948b4217fc6c3f09e6bff04b89e6f593d0312ec23f2dc383006513531aa82ddaacaf24fe84bd3cca49684849ca6d68af5ec20150e662;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfc27c57a0c41e7cdf614e9839972a03a28ee2cc1f48b0c01747b856f4ecd915d2089cba725e1ce77b57e60186221248c19f4b0529b0d71be9b2bb40317617ad176b1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbca4e8f7b5901d2456c6b7ddc54000cdb23df164539ad1228beb61a49743610c82df236670c4a2ad49ccac38ca9452ad2c69a2b7f054c140e183a1a08c7c58c0bc74;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h132d5603c9c353c3fe15f968ba942c0acea76a98ad13d80502a81dc3a1f8edb945355cb52136a084e32006800a874d8449258febe9bb27127c59daf672d29f52e0666;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h175a29ae5e7b258b92a029f11b087305a1a8d930932662b1af80584c675534bec26cbf6a16d27fb5434685decce85c475c7419eb62e549cf8a629274c358b5fc8f74e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e0d3e84f738ce6d697bb4f796ed6a70e2b1d0d1ffa4dd107785fc37020721cf16d0050c255f1b754eef4e983dc65f9eb4186608e32303789527b322754c246f4503c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11e523cdd3dffb4e4f3fdc29f307fbc9a22c4f09edf2355326f816665ba9f238606b787f3afee23ca1caebb92805cb9b2e4f9786cd3fb30d31dfea0531bb11ccbd9d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1fff663e517742f817e216a3ccddbaddb2f53b06d0eceb670b278fb560370adab53380c1d0129aa4cdd258132c5374ee44e6980a5073c0571082189f623027e89e766;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h5e450f1d8f221c5d2500b4cd579df2c3358948aa4e348263380d8490d3562a567ffaa818c6e0ca573960e9b36a7b3f111cf4faf14225efa1285847744eeb8795a2f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a1fb944216eca5f3f518e1aa2f4ec9fad1a35cc774fa53a633c33fe3913de3eca60e9c6a3a61b8576ed1ff31e8042371ba38b303e95dca0aea54c9c50d28ed13607;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h989bbd95b4980dac1d79c5dec7184978c72e96f6a261e873b34dab6432ccd8cf7aec8ecb8339756865e7e3bc3aa219d9175e7af8f97ff1072d84147c72b00e5de42b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc6cc1700a30193443e7fa3451d4094bda6fc1ba67c8762b796eecdc83294efdd06c64d98cf52ffd025706f6ebcee34e3324cee660c511d0ebc09eb6471e46cb7d6f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a97f1b9bf46574b3c450f0ff2c57c6f79ab8e1a0e6c93ce71238643ec3d74b8601bcfa31e7440b9bfe8f8e45e61903a118373d94190f546754de70f0e152edb7165;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16e891fc753c0416f1add83a508a316f0b5d4c93385e791ff32a96e127fff4444099fafa02c15ce4f9295bea26b14cdab8a6dab66c0d97bbbd148d5b3364cd280880b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d14f0ac65aae348f386d646a0c3b0a45ac4630a68475cd3af68f4609bc1a8a5ea05f41a9c6594fb7f86809f19954164ad1f39585c4b7656524745a6ae832f133eb37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h108b82321e7b277dbda1e2a687220f38ae4b1595fa1373cc76c25bed2586b79417468e835be9d769948727c3757c91b6cc85b4cd5351243d6b07f59b1201d28f0485f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbe8fd311fbf06aa4bbd813d66eff46b5ca2c6cdd9e8eb259803b410479fe0592e149b14a2d6ec79047fdbffea961414c05e1e3b27e25f0be4ef1ed6dbdea6a88e8f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h807abc379a55d4ea54302dead28bdfa351c83910a5a851849d10dbcf1ff1cfc20e1fb2fba9fbe858f389e5d556cbab2a363bf8b8027e6d23daa4abf605543451a1f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h128a2e0da95bb00eb892365e26ec1f2f434466f7d4053175a17efc817150989aca24145fb627d7ddb69af8fefe98e47a896093f209fb937ce672b1d87b2a571cdc528;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1664774a7b7afa4fcf569f0680ba3fccd74e78279a6705c3fc117dfacb54a3c5401eb3aa51a6dcdbd83f0683ca307ad91db8cb0fe78bcf15ed4d51a3368e417031bfa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h2c724517fc2bbcdec67b0356a5320ee345d26d581d3312c0f90907bbfdea1e74b572a98ffc7f5e51d60950900fc3280d3176a08a72e4654cc51fd033c8c5ee2824b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h8ba6264653a3bf65d2d8808376318de9de665383a4de482b877b86e219e9a2fe0ea4275cce6ff5465ea77e4a6e84b90616f8bebc6ac0854273a9acdb58f326c48ba5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1934c12ddcf8a076504f683dac38410aee101a48a173ca1e790f10a6732b6766b83a6cc03f7a38343d9521052984def987a395209fddae8a72aa027462b5168debd18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1dafe1496d1b982e02b5e9c5472453ab2316be1bdd2af701bb35a17306ae5caaed6651b8599ccd69a94d28b93257d999723f114f250cad3b0cf7326def8b4613eb8e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11a89512717a3c574ae75f6b68bf4fa20a329265d6d55b047c7ee782832cacd200b7df8453fc6e6640c332f8d9358bb916664bab56aaf8e3b917348e253694e7136c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hce79f828fb54a1c0ed281321ec94d965174a02b5c2111f83deb1c14fd89c7f0bd32f37481e6a18b219455d1b02d970361201d5a56b87b2adda37f890cc1e72609a9a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1e9f35487094a45c61caebffa79b6797b62abfb0ea9e8acd938b3cd52edb8c7f86d478b5069608abca39a4634a9123b30bb9e614d4d19d39b668613ff1f80a2e3bf9d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h16dcbca3f37d826fb7a06596c67250e3b13770e5ceea2ba47c2685decc3bd6d9eb1ba815c2017b655e96b2b0add5ef187f84db5c74390e38f8c0b8edd82cb57f0466e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hfa0d9d7a2765a709910338a45e39ab0844c2bed07a9739cb339bbad4dd17dbaa618d53578939cd975226a9a017d6af5808034238e096867ac96e67a155d0464635fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1edb3f7e3c84f132d20fbb778d9ec46ae8a3275b505ba8309a9b282d80f689d5fdd7eed652773aeaa27d7416dcdc56af2a335ae65810aff1714340fa67662bbe8889f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h133c0e626d1dc881c8ac6a57ed8eae8efd4fe8dd658153529537007108e6bac0bfa966f840bf2363ef2532cc6e254d24b76a513516442b2388c8b45e1bba12d06ede5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h39b646efc2f1b22fa4a358cf8bb928113b0f21dab55defffeb8378db704160c56bab2a9a12e6ac5702f18856affae5f8e0ebd6510fddb0f96481b4b3e9cb1c624967;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1409cc65067868160a888915702ae2393bd640f46cb6953cd45dd07c23234ac2f4b59e1ec50f582b47ad6dc798b52385fc5d605fc1e8576a8fbf0a9bb96b2c2b8b2d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1d47cb95b174b7cd3d1e8bf6ff7ae68bc88dbd2a632cc4b2eec526dd7e0613f709f0b25035428021c16ce26c0885f433478eaef21d0e20cba7176125af25d9da67d79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h88b2ad0a86cc5d691432ca0289a4c6921d361453a7ea8791d1407ac508db65d5ba8bd5e625c7d5f1377085361df89e7c9b18c82ad49117883edcbf33ef78369defc4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'heaf8ac58a456bf297224b8680f544cb0ecf06b9164d1020bfc865e240c51ca452ba3371f3f269f4ce94bd7ada139add6bb90bd0531bf464ee0dd571152c58f0ae37c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h195c28415925c0d06576c0e97245615d7079400fbf3bcf4c1ba67daf289f219cec33698ef897d28e6fb2ac8dab9b7c7444a21741d9fe1e3f252b1355e7e21d5b4c00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1b18118fd2432babf81db0fb19326a25dca7dc090498725c4095bcd9a1b3c88c97ebe18b2b5e325156544044b94a3ca03ef65d14345f8c766d35f29b35702c21c2bb0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h101af4043903f97201fada5a03a25e403898eaaabac4c41a3339775cc5281b62ed0f30a65735c834a7bf063dae7bd1a78b84ebb5b4da3636ab04401fd30c1d8812749;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f3a7364bedb7104335f6d5d5bc3801d16896cfdfff3c7830c71a959e40e17380cbf4fd31f93f2cefea3bbab4361bc6ac5f41d64d6942925d455b405f1675cf35da7a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb42767a817ce3fb2d8780064315c216b17d4549c14905f622010a4a05d850d72732fffc8054a30c24151891d3518e7622599b459314cbfd9bf16a289631741606c58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h151970ab78ba7754f8ce94b4b6d6b676f7e814bd67cfd6940ebc79229bbb66d51b51dfe9859a4b9002dba1c4ffca4eb369c6aab4e70893b9d11706bee899efd33639b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hb6fdaa35d1afd3e3312948825fe70f50f6217f601d5acd7ae8254a2618e3f2cb169c3ba79ae1fcc4215e1ddca6fac8797217401d58fec48fd0ac7e55e03cafc0c31e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hc731cff1159a7758317535d9a6333033acd713a1d0743f65ba758653b4afc470c409ee68041a5ff6faa32bf0d5f6676ce55e6ba5c1f78a19bcb48fa0466674b928e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h10714bbae45f13bc15007ad84b8f874d302c0b26fe8c0e6f29a0926f8b223c68b2ef1e6a0f6bc00bff5f7d0176afad70fd3ab4a2c1859141241f21cb6159f2356814e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1c35e7eef9e562cda624fffae3686e98349a1a77ed545d614f5045d1b6f3e5144de1a1d922477e382f00b3a9f1e2bab1dcedf08058e76d9b3924e805afaf197fbfbb6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h7a9c75e3bac7fdf4b42a4e1f017aacc436cf9caed22a682fd131c2b16bd4759db0bec38c0d397932f2f756972a8ad472088a37c91972a109e2bfb5ffba3512fc1315;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11619d8c8a3d286722aee26a35c9450566d2bba904b9462e4c39608ac906ebecdde73e40dc4e055e921246ac755e8efa2877add4ca9aa2749d03f983722ef7da1eec4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1f786bad0b647e950af31f4cefd6667b5b4569cc77bfd62502c2c13aa0d37de8bab1cbfd042a0e2849ef163461fbe71f841780787f450bd7b6e901f9d8ded7e0c74e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1a347905e3c709a9f0b7b31a34260c34d646359edf6dc85f5aeaba50bb29528447944d1b07ae591acf0cd7d326159ecfb8eced70f936c716cd1c7b331b86ab2b6e0be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h774fca45e880a4ff3a18602481b96831ae7726fb7c21577a998d78331cf3c3b85520fab24f4ea5eb45696db36315861f90232382f658c937717946312435d468c83c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h11efc360ce8dacab5538ec471a840b1b9750ae95020c6037ce67f548a3e929e1a90c10ba984f6b2d57bb60e36b951dda2fcbc400681e50cad9890b57b5a6d94e7087a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h148efef09f7b82fc1c36d94b1a36c8179bb1cd2a781f2bce5fa5265cec621b3dc0ee70eb371d92f67ab25e9b419c824d762b587e3249f1e21e28024582803fed1afa4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h1490310da06e3aac7d8e149f0a7750e05610745d5b825c7fd66e23561d4032c3ae83a724f1eeecaaefe6f465c2da26a123763588eef6fe8c0ed3133c061f6ed45fcf8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'hbcdc86453b6230ffca77946505c789c4a5cf4edbe6ce5c4148c603d3ad9be9dfa32f7f9cd9d75f8bfd5bd5c40634c9bd3d415d15f55d09ad33572cb2ce94087a3f13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h192b2a5b0bf4c0e95041defc7f9fc7ee9d2b91ef413c939268f6d3f946f9e210ec44e9fa86f3143a60e23e24ecd9871a188e270be911e70880b429bc2bba71ceeaaef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h85c9843dec73ce01eafce0cddec2b8663b62abb2009f4168b5e8b187d4c92106caa37c1ab6f1ae8a38a22e9561b205adfd4e163182d3d48582c5096c7eca20e3ece0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h742db5a1ebbe18cf8d226e5782ee6242453f27c043acfc7f34ea9bfb9fd7d606a9fc9b3a19fe77eed9de4333ad1316b18379ac055e11c42050d763407c6be5a5b3c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h14fcdd9690dea6c203ad924188e1640a2e81021904948ca4979ba8c9fdcc835db272b666a61f4596e434b5a5f2e6cd6ed93a88f67bb0880779dfa1e2550c48a09127e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'h140c29b94233fde93fd7df16ab9f7e9a48b6c0c3a229f767c0efe0507197bc6fa39de9390b712b1755cdbeeda049fcc388fa79c54e4611b76100bbe5bb50ba82a53c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 529'ha77d1adf3e9e1f2e89eb1b17fbe190a42e5a422d71ba79b65b211431aed6699a8cddd27cdf6d8fb119433308f42232a1117da764432d48094a42608e237500231afa;
        #1
        $finish();
    end
endmodule
