module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    compressor2_1_16_16 compressor2_1_16_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
        src12 <= 16'h0;
        src13 <= 16'h0;
        src14 <= 16'h0;
        src15 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor2_1_16_16(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19)
    );
    rowadder2_1_20 rowadder2_1inst(
        .src0({comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst0({dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      input wire [15:0] src12,
      input wire [15:0] src13,
      input wire [15:0] src14,
      input wire [15:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [15:0] stage0_12;
   wire [15:0] stage0_13;
   wire [15:0] stage0_14;
   wire [15:0] stage0_15;
   wire [11:0] stage1_0;
   wire [8:0] stage1_1;
   wire [11:0] stage1_2;
   wire [8:0] stage1_3;
   wire [5:0] stage1_4;
   wire [5:0] stage1_5;
   wire [5:0] stage1_6;
   wire [13:0] stage1_7;
   wire [5:0] stage1_8;
   wire [9:0] stage1_9;
   wire [5:0] stage1_10;
   wire [8:0] stage1_11;
   wire [6:0] stage1_12;
   wire [6:0] stage1_13;
   wire [12:0] stage1_14;
   wire [7:0] stage1_15;
   wire [2:0] stage1_16;
   wire [1:0] stage1_17;
   wire [1:0] stage2_0;
   wire [5:0] stage2_1;
   wire [2:0] stage2_2;
   wire [5:0] stage2_3;
   wire [3:0] stage2_4;
   wire [2:0] stage2_5;
   wire [1:0] stage2_6;
   wire [4:0] stage2_7;
   wire [3:0] stage2_8;
   wire [6:0] stage2_9;
   wire [1:0] stage2_10;
   wire [5:0] stage2_11;
   wire [4:0] stage2_12;
   wire [1:0] stage2_13;
   wire [3:0] stage2_14;
   wire [3:0] stage2_15;
   wire [3:0] stage2_16;
   wire [1:0] stage2_17;
   wire [1:0] stage2_18;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [0:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [1:0] stage3_13;
   wire [1:0] stage3_14;
   wire [1:0] stage3_15;
   wire [1:0] stage3_16;
   wire [1:0] stage3_17;
   wire [1:0] stage3_18;
   wire [0:0] stage3_19;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;
   assign dst16 = stage3_16;
   assign dst17 = stage3_17;
   assign dst18 = stage3_18;
   assign dst19 = stage3_19;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[0],stage1_3[1],stage1_2[1],stage1_1[1]}
   );
   gpc606_5 gpc2 (
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[1],stage1_4[1],stage1_3[2],stage1_2[2]}
   );
   gpc615_5 gpc3 (
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10]},
      {stage0_4[6]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[2],stage1_4[2],stage1_3[3]}
   );
   gpc1343_5 gpc4 (
      {stage0_4[7], stage0_4[8], stage0_4[9]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9]},
      {stage0_6[0], stage0_6[1], stage0_6[2]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[3],stage1_4[3]}
   );
   gpc615_5 gpc5 (
      {stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14]},
      {stage0_5[10]},
      {stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7], stage0_6[8]},
      {stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[4],stage1_4[4]}
   );
   gpc1325_5 gpc6 (
      {stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15]},
      {stage0_6[9], stage0_6[10]},
      {stage0_7[1], stage0_7[2], stage0_7[3]},
      {stage0_8[0]},
      {stage1_9[0],stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[5]}
   );
   gpc615_5 gpc7 (
      {stage0_6[11], stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15]},
      {stage0_7[4]},
      {stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5], stage0_8[6]},
      {stage1_10[0],stage1_9[1],stage1_8[3],stage1_7[4],stage1_6[5]}
   );
   gpc1343_5 gpc8 (
      {stage0_7[5], stage0_7[6], stage0_7[7]},
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10]},
      {stage0_9[0], stage0_9[1], stage0_9[2]},
      {stage0_10[0]},
      {stage1_11[0],stage1_10[1],stage1_9[2],stage1_8[4],stage1_7[5]}
   );
   gpc1415_5 gpc9 (
      {stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_9[3]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[1],stage1_10[2],stage1_9[3],stage1_8[5]}
   );
   gpc2135_5 gpc10 (
      {stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage0_10[5], stage0_10[6], stage0_10[7]},
      {stage0_11[1]},
      {stage0_12[0], stage0_12[1]},
      {stage1_13[0],stage1_12[1],stage1_11[2],stage1_10[3],stage1_9[4]}
   );
   gpc623_5 gpc11 (
      {stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_10[8], stage0_10[9]},
      {stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7]},
      {stage1_13[1],stage1_12[2],stage1_11[3],stage1_10[4],stage1_9[5]}
   );
   gpc606_5 gpc12 (
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5], stage0_12[6], stage0_12[7]},
      {stage1_14[0],stage1_13[2],stage1_12[3],stage1_11[4],stage1_10[5]}
   );
   gpc615_5 gpc13 (
      {stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage0_12[8]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[1],stage1_13[3],stage1_12[4],stage1_11[5]}
   );
   gpc606_5 gpc14 (
      {stage0_12[9], stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13], stage0_12[14]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[2],stage1_13[4],stage1_12[5]}
   );
   gpc615_5 gpc15 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10]},
      {stage0_14[6]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[1],stage1_15[2],stage1_14[3],stage1_13[5]}
   );
   gpc615_5 gpc16 (
      {stage0_13[11], stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15]},
      {stage0_14[7]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[2],stage1_15[3],stage1_14[4],stage1_13[6]}
   );
   gpc1_1 gpc17 (
      {stage0_0[5]},
      {stage1_0[1]}
   );
   gpc1_1 gpc18 (
      {stage0_0[6]},
      {stage1_0[2]}
   );
   gpc1_1 gpc19 (
      {stage0_0[7]},
      {stage1_0[3]}
   );
   gpc1_1 gpc20 (
      {stage0_0[8]},
      {stage1_0[4]}
   );
   gpc1_1 gpc21 (
      {stage0_0[9]},
      {stage1_0[5]}
   );
   gpc1_1 gpc22 (
      {stage0_0[10]},
      {stage1_0[6]}
   );
   gpc1_1 gpc23 (
      {stage0_0[11]},
      {stage1_0[7]}
   );
   gpc1_1 gpc24 (
      {stage0_0[12]},
      {stage1_0[8]}
   );
   gpc1_1 gpc25 (
      {stage0_0[13]},
      {stage1_0[9]}
   );
   gpc1_1 gpc26 (
      {stage0_0[14]},
      {stage1_0[10]}
   );
   gpc1_1 gpc27 (
      {stage0_0[15]},
      {stage1_0[11]}
   );
   gpc1_1 gpc28 (
      {stage0_1[9]},
      {stage1_1[2]}
   );
   gpc1_1 gpc29 (
      {stage0_1[10]},
      {stage1_1[3]}
   );
   gpc1_1 gpc30 (
      {stage0_1[11]},
      {stage1_1[4]}
   );
   gpc1_1 gpc31 (
      {stage0_1[12]},
      {stage1_1[5]}
   );
   gpc1_1 gpc32 (
      {stage0_1[13]},
      {stage1_1[6]}
   );
   gpc1_1 gpc33 (
      {stage0_1[14]},
      {stage1_1[7]}
   );
   gpc1_1 gpc34 (
      {stage0_1[15]},
      {stage1_1[8]}
   );
   gpc1_1 gpc35 (
      {stage0_2[7]},
      {stage1_2[3]}
   );
   gpc1_1 gpc36 (
      {stage0_2[8]},
      {stage1_2[4]}
   );
   gpc1_1 gpc37 (
      {stage0_2[9]},
      {stage1_2[5]}
   );
   gpc1_1 gpc38 (
      {stage0_2[10]},
      {stage1_2[6]}
   );
   gpc1_1 gpc39 (
      {stage0_2[11]},
      {stage1_2[7]}
   );
   gpc1_1 gpc40 (
      {stage0_2[12]},
      {stage1_2[8]}
   );
   gpc1_1 gpc41 (
      {stage0_2[13]},
      {stage1_2[9]}
   );
   gpc1_1 gpc42 (
      {stage0_2[14]},
      {stage1_2[10]}
   );
   gpc1_1 gpc43 (
      {stage0_2[15]},
      {stage1_2[11]}
   );
   gpc1_1 gpc44 (
      {stage0_3[11]},
      {stage1_3[4]}
   );
   gpc1_1 gpc45 (
      {stage0_3[12]},
      {stage1_3[5]}
   );
   gpc1_1 gpc46 (
      {stage0_3[13]},
      {stage1_3[6]}
   );
   gpc1_1 gpc47 (
      {stage0_3[14]},
      {stage1_3[7]}
   );
   gpc1_1 gpc48 (
      {stage0_3[15]},
      {stage1_3[8]}
   );
   gpc1_1 gpc49 (
      {stage0_4[15]},
      {stage1_4[5]}
   );
   gpc1_1 gpc50 (
      {stage0_7[8]},
      {stage1_7[6]}
   );
   gpc1_1 gpc51 (
      {stage0_7[9]},
      {stage1_7[7]}
   );
   gpc1_1 gpc52 (
      {stage0_7[10]},
      {stage1_7[8]}
   );
   gpc1_1 gpc53 (
      {stage0_7[11]},
      {stage1_7[9]}
   );
   gpc1_1 gpc54 (
      {stage0_7[12]},
      {stage1_7[10]}
   );
   gpc1_1 gpc55 (
      {stage0_7[13]},
      {stage1_7[11]}
   );
   gpc1_1 gpc56 (
      {stage0_7[14]},
      {stage1_7[12]}
   );
   gpc1_1 gpc57 (
      {stage0_7[15]},
      {stage1_7[13]}
   );
   gpc1_1 gpc58 (
      {stage0_9[12]},
      {stage1_9[6]}
   );
   gpc1_1 gpc59 (
      {stage0_9[13]},
      {stage1_9[7]}
   );
   gpc1_1 gpc60 (
      {stage0_9[14]},
      {stage1_9[8]}
   );
   gpc1_1 gpc61 (
      {stage0_9[15]},
      {stage1_9[9]}
   );
   gpc1_1 gpc62 (
      {stage0_11[13]},
      {stage1_11[6]}
   );
   gpc1_1 gpc63 (
      {stage0_11[14]},
      {stage1_11[7]}
   );
   gpc1_1 gpc64 (
      {stage0_11[15]},
      {stage1_11[8]}
   );
   gpc1_1 gpc65 (
      {stage0_12[15]},
      {stage1_12[6]}
   );
   gpc1_1 gpc66 (
      {stage0_14[8]},
      {stage1_14[5]}
   );
   gpc1_1 gpc67 (
      {stage0_14[9]},
      {stage1_14[6]}
   );
   gpc1_1 gpc68 (
      {stage0_14[10]},
      {stage1_14[7]}
   );
   gpc1_1 gpc69 (
      {stage0_14[11]},
      {stage1_14[8]}
   );
   gpc1_1 gpc70 (
      {stage0_14[12]},
      {stage1_14[9]}
   );
   gpc1_1 gpc71 (
      {stage0_14[13]},
      {stage1_14[10]}
   );
   gpc1_1 gpc72 (
      {stage0_14[14]},
      {stage1_14[11]}
   );
   gpc1_1 gpc73 (
      {stage0_14[15]},
      {stage1_14[12]}
   );
   gpc1_1 gpc74 (
      {stage0_15[12]},
      {stage1_15[4]}
   );
   gpc1_1 gpc75 (
      {stage0_15[13]},
      {stage1_15[5]}
   );
   gpc1_1 gpc76 (
      {stage0_15[14]},
      {stage1_15[6]}
   );
   gpc1_1 gpc77 (
      {stage0_15[15]},
      {stage1_15[7]}
   );
   gpc606_5 gpc78 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc79 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc80 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc81 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[1],stage2_4[3]}
   );
   gpc606_5 gpc82 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[2]}
   );
   gpc606_5 gpc83 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[2]}
   );
   gpc606_5 gpc84 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[1],stage2_9[2],stage2_8[3]}
   );
   gpc606_5 gpc85 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[0],stage2_12[1],stage2_11[2]}
   );
   gpc615_5 gpc86 (
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4]},
      {stage1_13[6]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[1],stage2_13[1],stage2_12[2]}
   );
   gpc2135_5 gpc87 (
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10]},
      {stage1_15[0], stage1_15[1], stage1_15[2]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1]},
      {stage2_18[0],stage2_17[0],stage2_16[1],stage2_15[2],stage2_14[2]}
   );
   gpc1163_5 gpc88 (
      {stage1_14[11], stage1_14[12], 1'b0},
      {stage1_15[3], stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7], 1'b0},
      {stage1_16[1]},
      {1'b0},
      {stage2_18[1],stage2_17[1],stage2_16[2],stage2_15[3],stage2_14[3]}
   );
   gpc1_1 gpc89 (
      {stage1_1[6]},
      {stage2_1[3]}
   );
   gpc1_1 gpc90 (
      {stage1_1[7]},
      {stage2_1[4]}
   );
   gpc1_1 gpc91 (
      {stage1_1[8]},
      {stage2_1[5]}
   );
   gpc1_1 gpc92 (
      {stage1_3[6]},
      {stage2_3[3]}
   );
   gpc1_1 gpc93 (
      {stage1_3[7]},
      {stage2_3[4]}
   );
   gpc1_1 gpc94 (
      {stage1_3[8]},
      {stage2_3[5]}
   );
   gpc1_1 gpc95 (
      {stage1_7[12]},
      {stage2_7[3]}
   );
   gpc1_1 gpc96 (
      {stage1_7[13]},
      {stage2_7[4]}
   );
   gpc1_1 gpc97 (
      {stage1_9[6]},
      {stage2_9[3]}
   );
   gpc1_1 gpc98 (
      {stage1_9[7]},
      {stage2_9[4]}
   );
   gpc1_1 gpc99 (
      {stage1_9[8]},
      {stage2_9[5]}
   );
   gpc1_1 gpc100 (
      {stage1_9[9]},
      {stage2_9[6]}
   );
   gpc1_1 gpc101 (
      {stage1_11[6]},
      {stage2_11[3]}
   );
   gpc1_1 gpc102 (
      {stage1_11[7]},
      {stage2_11[4]}
   );
   gpc1_1 gpc103 (
      {stage1_11[8]},
      {stage2_11[5]}
   );
   gpc1_1 gpc104 (
      {stage1_12[5]},
      {stage2_12[3]}
   );
   gpc1_1 gpc105 (
      {stage1_12[6]},
      {stage2_12[4]}
   );
   gpc1_1 gpc106 (
      {stage1_16[2]},
      {stage2_16[3]}
   );
   gpc2135_5 gpc107 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4]},
      {stage2_2[0], stage2_2[1], stage2_2[2]},
      {stage2_3[0]},
      {stage2_4[0], stage2_4[1]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc1325_5 gpc108 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[2], stage2_4[3]},
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc2135_5 gpc109 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0]},
      {stage2_10[0], stage2_10[1]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[1]}
   );
   gpc606_5 gpc110 (
      {stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1]}
   );
   gpc1325_5 gpc111 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4]},
      {stage2_13[0], stage2_13[1]},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[1],stage3_12[1]}
   );
   gpc1163_5 gpc112 (
      {stage2_15[1], stage2_15[2], stage2_15[3]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], 1'b0, 1'b0},
      {stage2_17[0]},
      {stage2_18[0]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[1]}
   );
   gpc1_1 gpc113 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc114 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc115 (
      {stage2_1[5]},
      {stage3_1[1]}
   );
   gpc1_1 gpc116 (
      {stage2_6[1]},
      {stage3_6[1]}
   );
   gpc1_1 gpc117 (
      {stage2_8[3]},
      {stage3_8[1]}
   );
   gpc1_1 gpc118 (
      {stage2_14[3]},
      {stage3_14[1]}
   );
   gpc1_1 gpc119 (
      {stage2_17[1]},
      {stage3_17[1]}
   );
   gpc1_1 gpc120 (
      {stage2_18[1]},
      {stage3_18[1]}
   );
endmodule
module rowadder2_1_20(input [19:0] src0, input [19:0] src1, output [20:0] dst0);
    wire [19:0] gene;
    wire [19:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_17_gene (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(gene[17])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_17_prop (
        .I0(src0[17]),
        .I1(src1[17]),
        .O(prop[17])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_18_gene (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(gene[18])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_18_prop (
        .I0(src0[18]),
        .I1(src1[18]),
        .O(prop[18])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_19_gene (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(gene[19])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_19_prop (
        .I0(src0[19]),
        .I1(src1[19]),
        .O(prop[19])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI(gene[19:16]),
        .S(prop[19:16])
    );
    assign dst0 = {carryout[19], out[19:0]};
endmodule


module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor2_1_16_16 compressor2_1_16_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5033fc979927d48c1a3e6b09844e6fd52a08c310e97dd271437a9fcbe5bea775;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h239244496bce11398eeab1938ffc4a29694cf9de2e18e8178347ad8884723aeb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8522c40a75d87067d6c3a0d420c27f7ffdab1b29fd3e3a6a7c2fa1220bbec76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6437f27a8380881375a964a48aebcf9c8071d204fc098a5bfb48477385f0a05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he09de47b7cbce124fe17213149e7d34c577da709917f120b9acbfc328bb033c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h950edb9ebfcb91eac959ac346622aaf40549c4c659bb2f945974eb388ae478c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7dda9c5d7124c6efdae7c5a4ac404c7afa73b2841bf3eed7c9253aa6c6c0c00;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h697d7e1100a0b24ea8567efd422b40a88a696ca99a6e48b477ea11857e5d4777;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1dce738e0e20e29215075b164170a7004d43224fbc6f722967c346e3cc4994d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6290c8681f2c29a2bf172e41c924171d4cab2c22c9fd05794d33b5e1dbfa8db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcee86fefb1963da8d02699f4fd30397ee44db4729d9412447c500baf98ecf8c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha82e80cd404a46be6c5af612e29818b2fcc9d839daa3f9ff2fbbc768d10be86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71aa569dd09e18272cd3549cef51a295fa0db60bc2d46abdd461ba396b811789;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6d6ab659f64043d8d2d42e160f0b2c217e21f203e18b6bb3d748aa9aadb81a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc270f76c6ba1df298481adef6460a0d97091788a8ce7e5398fd35c5536746e1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd02c70ad7f3a2bbe073b5dc7df29f0c8fa0632903c67a11d6732545a2c289b65;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47f39f267be4505c61faa0a50eae2277782ed6a4498b9ecc39f8b53d8b43cef4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8fdeab6e5abd9b0d350c265ef739e1744cafcb6e9b186b18b8b70fe295371c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9208a52799cbf443dbb0335f525626602a7f362d96653a0972998647d8021808;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21faffc90be022fe3d3ca5999f05fbeeb96a9345caa953b4e9a38f9f0c1263ed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bbcb6d2e78148f95649798880d6e72812f2686da4cef16e895fa8b9fecabc7b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6a1c85b61d2b1345b60839caecc69bd3d6c0076cf79539a5417ede961354bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a86b8499e01041f104d168924032eb4ab2a8fa51cfa7e6a9a975fa93980f260;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87d2be2a883b65d6a1c7029f2702f5a0bc0cf7a4d8a3d1af30534031f81f8710;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37e62432ee966d2989833ebc3a2726ec7bce37fa6786c8119be7dc233fa44d28;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1e84a0410c84bbc98f6484911447dee24cc9846a08fcb607994a6aa352858d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b5bc576a27962b69434604eea575085f242486b3170ad58e344bdebe5ca8014;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5efb1825c4066e3ea8607a30b08c9ab0cefcb448c63f8753aaf1b91969d54cf3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h670820c9a0cbfca2f1b69ea0e54b3ffca244388a6df5cbd3b3686297a6e25473;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17ac52776de10d88b89ac04744b2831e5558cfcc0ee2c130872427d7910d6a09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9df7133f9a96055f09786ec472bff696fa6bc92d8d5e93a126775a803d771cbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac93248fc3b553c09364bc44b81caed1d96908d3eefa217bd220f9a2091b6cef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h314fc7b760c2d68446493280d318a7f3b536eecaf37aa9c2fd7ff122057165ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5a0336396a8cca882dfedfba625cbea6da998c29fc3a2ddd73e5e6f464616f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5c1202d3d1ec3ddef0c0ea2884ee841a96e6c0b977635425ce23c587c0a09b48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4928e64b7e1adbc93c3a17aeff02dec3e19113c134329d970e98e55a4d4bab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82df2e6508f59c2ca9fe48460913ba4a42eb80b2b31060b644341f3af8237f30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9464bd9b321908f4be6de3fdc9ed35f9f65baa656720766b9b8b7df9b829cfa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52f60add29059ac7d5b3ddee9eee99317683ce6a5d2b435f2001494f91603a9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e80e536fba73b4c23151b28feb2b6862371cbb31dd95cf373cef9fc52935fea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6134b5d8d8ecd16d172630e6ce863c96ca0dae70038dedf5e96993d3e7d1500;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h830384b468779510152aab24223c788956858a18434759874110d2099db3f681;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6dae495bf8d9e2b6069ed260e59618bb8ac1c580f5b322e88792b3d88d0bdc66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h290418951cfc0eb052e24663c3133b0b8fd06b750a02418982f6f3ca90162aa0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3fd8d91c890a16b490ff1c44d5b7cad7a5528bd95e8d47a8a89a2bf67ce5c814;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he53f4b15fca5a2a345c12bf3b9ffbffb21b9938675a03b9cee360b28eb9aefa8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84b2d768c80d5f659f7b4d743a0f9d14ff31a576d5b9ff49f0c36e90ada70e0a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd780a8b1dd356a03b6be3fd61afd8ebe32d1f2e701f17f2545451765084ac960;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdebb96f26c49e6d8dc70acee0c7f24179ed7ff0324efdb9ed8e41522491540c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e2cc21b91576dcd7508220132fdc36a769b2fcfa406e42b364bb4c08024f3a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e65b4fddbe43f143e7143ae5c06c599e71e97b1c8b47bfa66ebeb14b18ad003;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha33eb7db63957dfafbb6eefd52bf7d7454022da6dcc54c5588ddce34ba2c9aea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7bffec3fcac68af28d7e29dd0f8621eccefd1d92f558ba6ace52a0d869e4b38;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf6be74a4c835dbfa24395c25413f7277701684410d8ea27cc379b20d7e62ad7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12bbe15ee2b24f8270340eb8365919ae2d48b7136d827fb0d0f9d46c329525c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h961cf88fac63d8ae0ed706764540a5bb22fa3a128431c11f1e7f0a20a5e986f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff7baa8f6548205b629b15015ff7ac6fbe14f2e5494cdc129d46b2eec11b2a47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9275d669753e697c430ac7baf30186e590a3f45aa0f87e347e55c27740a50ea8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c33222edbe3ce91bb4b2c20e9e78ccfaab5e5ac46db92715a5a8b0dc5ef75e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61ce59789ab7ea3c70483aa222acc8ef53ec67900d623ce7f34a881342b550e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h339e0fa5f8bba92f21633aaade453f02e73ccdeed8c1a8bd0154900395f288a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha67aed619b49ebbc2d0386dbf0d8cf930d964bcd87b9540554b4a07c4492d1d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7c43ba6bb3aad22ec3dc6948211fe0152a7f28ac95dae53443b713bad9a5b6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbfd002390d8a6cfbb4c092aeee645bcb3316cfab8eaeaba8beaa32825d6c36ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ba7f8393e743639e53bb85c4a675d33cfe6eb267e10c515cdfab6dccb1c2971;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1a52c5509230e836cf2319d49f8fac7eaf6efe8d3980d7d023985c56f192ca6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe4a0859b4a936899af822132ea6bd9811eec52f6fecbb5606d23f3f82e1c1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4113abdcb3b22673abd92f1a27f24962d8bd2ae837721fd07dd752d6bf78c7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8eb2af7c45aef1968ced61777cf78ee30b9fd56a1ae4ce72344650f65e346664;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha85907b522a6cc637140d39891b6a140a8dcd8eba00f937f5f82781896e600d7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3cadcc683c2a29e1106e1907c9ff9785a599e4230ad65e6bbcda8d300ac70b2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59c8ed99f8502d8d8277b1cec2918e337d8aa3510508a3bea5cdd3b666dce7a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32a8a0a17a2be3ca1269470205f00a6d8b87536b3982de64cf219c5a2c9269be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb94dcdd206fdf9acd14cf866b531a6ab1431dd7a1e95a80b8ea80173449cdd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbe39f22adfd6fdbe4bba43f4f90fc958594ac034579472ea1eae618830c7ad0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haea1630b1b1faf32e6eec3ac146b1f253a6b20246bdc98463a842cc8af4fa721;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6175aa3970c60e4bfc0155f63733498bdf14cf6b65c6b1407272098428342f0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8567c44b4965b2a794ab93add71d26511a41e939bbd145afa5d2e00b28639adb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b7bfdbda3b91bbcf296b0b2d6608bcb5e4137b9ff2f366c0db8f899f9f33e9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc511b2d0df21cfb69153cd3b96f5b4e381ab58e2b982172405e318e0c107f0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac0a0635e48ed67251d1a240c43c0429760b42eb9e030bbbdbab32f6b7cb4627;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc670b79ba2898154bb09a0585bc92dfc24df25f1935eaad1010f687ede726ebd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd9fd7be4d4705f476a844da12679d9e81b298fee98aead117ea90bfc57e39a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ef63fb458364b93b24a5b3a4b5e594f275cd64c92376eaa1765521c57223b5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5cf189d694652d93f31a8258c1c6fca865bd06c75676e7e597cc624347a0337;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74e9a49242f05658fb12e35e7e792208468de8001ae37c686dffb93f8c3ff534;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h200ec3306b7a59ff1b03e036516ca81ebb5564de0f34440844f8ed19b873a3de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e0c9038ec6b6a42a83fd7f4f49d11bcc4040f88d8174e52d208761c75c445e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21275d5e434b73b62b2df3056ed3fe1ea00422beb8e57a7479138abede962939;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h48eef577d6e7d4983552bae86360bd8169a77de84c6a0c3919062aa49bfe41c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ac25b62c1eb7e24343eb81f1b1de2518259491c798aafe6a7f3b701fb0539e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdef6a715bc22baf747935dffdff99dbf6e70e943337b2f052605bff82438d579;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda8edd11caf1637b024882707b459649f151ab01331ade19a8b3a18a519326ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc7a003d5ec7214268c2705cf9e8ab7d8dd8e192ee23a330040f874d4dadb6511;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b01cad91f726b8ac2dbffef45e1f2d0e0d60ef973a6619ea5c4c90a4bee023;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93358258a5ed6d1a9f4e105812263906f7aa794e067dedca5f146fb8a2a86e6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4e3a8240778f1a1d2cc4fa4f7d2297933db9220e3028f6c285672642a44df15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2cd3428c4993b0917755300ea38f35a118571e31e2edf093a2f4d80be6579b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8dea9b8f68d79acc27db5ad38ec32dc5cb2fe7b8071db7484bd5f5a73a199203;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56f1075535c09c5b072dde96964665e01ddd6d9b2fb19aef227f8afb968dab26;
        #1
        $finish();
    end
endmodule
