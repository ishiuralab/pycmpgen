module testbench();
    reg [23:0] src0;
    reg [23:0] src1;
    reg [23:0] src2;
    reg [23:0] src3;
    reg [23:0] src4;
    reg [23:0] src5;
    reg [23:0] src6;
    reg [23:0] src7;
    reg [23:0] src8;
    reg [23:0] src9;
    reg [23:0] src10;
    reg [23:0] src11;
    reg [23:0] src12;
    reg [23:0] src13;
    reg [23:0] src14;
    reg [23:0] src15;
    reg [23:0] src16;
    reg [23:0] src17;
    reg [23:0] src18;
    reg [23:0] src19;
    reg [23:0] src20;
    reg [23:0] src21;
    reg [23:0] src22;
    reg [23:0] src23;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [28:0] srcsum;
    wire [28:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2714937292f34d8c599ecf4fca3970ab6271375799e81390d1c6fa98b5c4abf348935d96f12a47de77855b3e9e76c744d2365bc6a660d125d428b43c64bec948b07b02bcf2af24fd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0a94f33ffe2e740c00dd26af91284727e8a03b7888ef973b7ff975486aca2ace49690ea40e4ccb378a15c35c6cfba399110cbe08bacb7efb89c781d05f031cd566c2baaa2197135;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c06ef5e434e36b4d06f84d120bfc2e819505e853e5da4bb8258d367779fd980013bae3a1b82ef52f244712c5feaf89ec48151f98190149326942f30c2f2b4ac45a7d07560b6f7c9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h795888efa3a15921c64ebef0973277812cdf9f15a5d86c1e7c3438dc8d0359444b7ce55d7dea66490c8ed5e115515078d501b03624561139902a509d84b829c49e6a45c115d67aa1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73a0a1920c25eaf677ce99e0d1f80a75b95d9726b2c96b210d5f0c423a40e2d8b7a62d24dcaa1f794a5beca0df54ca069588651665f19340310b2d0e3c94c51c95a25e009ce0d4ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f0f0950effa474e35e34a33d5a1027bac5cff8d6057d5afaedbd0a7e1d189356a85849e8a385be4f6c1acaad6fb47f307d9aaa84d24f2bb46f2d13de139ff24e471471c354ea358;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1d4ef34cd058e56113a5ec5368969ebb1b2471322cbd9f394c7bacd1cc75473038b7b65df517e473f26bb04138fa27a1095941e904cc2e7945052619dcfd583873ee7cfc9e73000;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h748ec94ab16cb0005cb1e42476e589a6fd5e024f8b04251d7b184c93d1cc3c8feb421c1dc69875b5abf3b856c5e3e15662a72fb50282264f98bea7dbee3a327b16322fed32a09b0d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3081e196ab377262665b0dd47ba86e8a7e8796ad5851a816b0ed2633392f6b396e6a176bd0e0149b0f9a3165add88bd01ee5b3cf5b4a675a649b7781382142e8acac23a2e8751ec4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac5d4f88b9ef6aa64cde742a8d00277ae948735c37d2a3917a3c2ea65dbd7c5858237b2f7d74e8577a8a4cdc04bc3e76156e4b6e355d496c0bf8bf5e03cd816060e04f50611548f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h443257c2ac766c573e9fbde920e8cd20693a91a92e7aacce44c38b5214c6add649d1885d70ab81ad61ecc748962fc14692a18d5d6adec78d4b793dd47f6001ae91e2ecd63d6d152e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf0e4ae41a7d0fa9db75eaacd00b440ae5fb04015907443110306b715be0921771906ff89331e99b12058cfe71668cafc8a8091434a5dfae7eba6ae86be932e2917fe802bc30789a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78e6975f565eb50e1170f6a58be368dd523ed27dcaacab061df8322a65848bcecc0dd06a6c11b027a86000bcadd908557558cec0834fce5d0807d4ff0176243e0ce144039a7395e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9549c2631a01a198cd2aa5c3f09e645bf75e46609f3854269ae394dca51dd0a9617551e9777e3858bfa2b263957a2bd58d3cac2c8a8605c43d819feb94fd8d778821232d80d491e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e2aa3c3a64d62d3f57e265155bc588625e393dda5a6daae972a2b41af4c651f75deaddfdf7abc8f3b0f243082da7279c3c7ef2a8fe678285212f0fce35b1992f3966170d3bf3ff4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h573bc7fc36f437695edd22741ad01c679f1e19bb52a0dde65117e46277795e535c25df1916ab475e245c4175cf003c81947c14e1631f91fbee6299114da767998d1aa1ec9083d900;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7072f0f48727df0a035cd7e146f2baa7c0f2d58e1e68760e3dbb40b13f6758ca687db848c5e65ffda3997771d4286448ac7740e209d7eec9aafded98c3a3ef2aa4f822bba18351f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c63cbce82b860c733783150767baae79f5afa207ea8c3b1fd6b8d02b3c5990a25674924584597d7694138cfe43a9e7afda3d05f1cc1d28920971d19b5dae0da60468750c01f6ced;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec30d0cb7a0f6fad52059ae81f428471fdcd8cc5339c95922a484ea490608def3a12c88c1d0463dc0a0b700149bbc4d910530677eb5521556588b40a5e3983dbf71f0bff769a0e04;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19d845a9db60ea7188a525ed6307c292edaf85e1bc071105c8cbd0734c25deb85771a322e97589ac2f91aa35f94d74ef039a77a33b232083b03f5c22ed41bb61f5cb67256f8a3178;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heff7f0906dff1e4a290e7605413c1e8a089027d8c25f57ac652de4268e5097eb41773947d4bc28c03f04aff5cd08127e906506947d7dfa38ae1589efc3ec9dc87127e9935b87ce8c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he37f1d032c6b532ba5cb2ce6cc431fe16ddc2393da44455ef060d467c85800e97d1102fb636dc90d7c88cfa36e3c81be67214f1fcf85e849d607a0f7be9e8644dd8384d6da0f5dc8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h369b5039ca79be70cc34ba51b3e17e97b0ca55eb9d9268a4df23b771e04c83d6c9f5c28a24e8b27172495f5a90a24fb1c77584ae9ebb9538abf1b3a0563aba6a994f0d57f99b3c98;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ba0ea14b05fc13d344c52a0ca6ae67062c7c5b95af43d6485036c30bb0e7999bdbdb7218aadeb70326e6b83265026eb293a29a617d176115d39bebb5d4ef454573ed643f6ddee0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8bef672eb0ee8248266e9639b78e9f23c0b1daa95aab9759ad406cc7a61325323472d80f6a2c1d9b661e856a5e62273a96eb01bd32ab68b4d0ceb694535d95212ffaa48888611ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3828e7682dcc1e91358721f30a4621ed9027a2b1b4806f99af4ff51cfaa08f43c8e3cb2fe8ea8e3f199be388789d6c37c967867c67b068256d2ecc999df0ede7592ec4b7d7cfa9d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha88c38c43012cf8150290e393138354d3542dfc1e9944006b1dbb25b04d328b90d3957d9336fddefcc712f250f5a5c45611e43b1d8a34d29846408947e51fe5ff4803c486bf7d192;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haba0fe8775d0a14d6e8fcb6bf75bbd6a889fca60f1129fab5735b564199c8b804deae73c48f8ed780ed15e5f2c42b573ca9b5c92dbdc476ce86c0ab69f8fc39bf7db237c6bbc7d0a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ccd0da2c17c409e2062b9269a896ce4034272d1853fc647ded6e7ada3afa36f6d13f39d164508e391420aedc47337fd11917f3a41f26e9d66d4c7046f0f0e079908557069b2cd33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36a1fbed677ce3649f35ff1e629a7793659c2767fd52d7a045b9b77b9644ef80c85daef49742b19ed1f59f9d71777e565b6ff9d893db6e66026ab33aa093c93c09206c42d0895fb8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e563075e0b2afbb7f3ca7cf5c5367bcbc9da13cfd38cc92c479cb4b2bf0eed06c52a5c4b12a9a8a760a159295e3d47efc41760a6cfea99513d6431c93daf7c052801c105741a6d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hacd046f24852efe23ee357479e52e665095a2bc92915c80fa5d6d054f68fde4857f7e1d16750ec407b45f8ecfc2d0ab21c1031efd9f91cee576b7dde6e91106c6e52aaaf34224ec4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2d8c42faaef5bc5393ba5124f8dbf7a6303fb7f57412c570e8fec95771fd78db880f075f10ad5e7d2ad62dd12e57f824090c3c746c159b406437935122b172815617ae938f63109;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55a8416d3e4ee20e35d7f1c767b2bd76f03310003aa2adba00f3c86c72f13e06e5c2084ae8fe140afdb10b755d4ad64df4d4b17f1e9cc3610a61444a1c1199d360e543fd6fcdd734;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34669b34dea0f1cdadbd815ca92645576432c7e15c6e909b5bc48b58d65c21820e99da10e8fdd3c635af40e9d3a7f926f922778d2fe5cd64a2ff3bbe3344440485b47e0d3640892c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ab157124633bcff4d7479fcf2170b74d48ad6df5840526e163094b623cc080eed25a4e4209b3288b7d92ceb05fbb88d82578d1d931a3b9b702c2309ad40e037889b0f2afc3e6f8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf86aee52fc65356a26c06d5da62c1f74d307b9d0aeb36229d69924670120252a748f641466edc4e42f79fd249873570b1aab837c58334b26358a68588ec85b41d050d75b79597806;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d20b1ecac4a9e2ebe41ea8cb5be4779f6306d6f7e011ad0159dc0a58a23a0a0eb9bfbf6469bb0ff8dc9e5c7ea27dfc0289bc8e0b69fb5d60c9fa1a3fbc8696c5c21f9c50f48b135;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66a5dbdbe9ccdffbe9d0250fb57729caf7e529f582b7b9b96c5ad0ab31864e2396ad7b8b8b5b719c0d19b782a77b9dd4f431b97bf46b46d8ddd1f0192359fa767f3d1fda4de38a01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc7e37638ff82d27866d8d5121637468a671c0979f060b7dbc13cc8a9d735e3047c6f1088183a31dd3e5c2481136a7bd3bc55c9df93a980a04f430739cc0c28dfc1f40c8e420e887;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6c4cacf50a2e59da07bccd7e69af9c55f47f99e23d247e68d24e031f2a598b2e24821569c0a270aa16e56a0588d2034be801ea58475b0fe809798dafe40401ea83c4ef7fe464905;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc99c103959e1fa05e336f332ecb1bb6b46c6485156454684ea6e2eda210e361237dea4224dac3eafa70196329014528a87a10dfa016aa917920fa2c819128045090687d3e754362;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3795644a2ac6b1eb4d218ef3024e1da5b8e560bb3fb62ea036f6ff9d56433a190234a7c5b1ce9a9ce579f7e30d2afe952c5e7bb12b0aa9e70bf4ace90a3952e1c51d5c40291eb0fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85e0300d961456feaa408f47d07348a30ea3b29a92a8fb3be6c4e78a763dcfa725e32ad5cadb9ac1b2048c755a55a0943824df444afb38ae016cbb50ef12af68d88db71c1735027e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5758784133e5963f8d438fe6077a25dabc56ec05cf10bbaa00d55b938e3658a96b27ef7c5af15b00464ae6b59d912d641bd2bce1d936e94befaeeb743d21310e14be8be22c86eebc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4aee8787edb23aa05c3fee636f6b59254c60602e8d5b885d6136ede7fca3258c7064b03ccebceb63f144f16eb915907c7548cc6a3cdcee5a06e8d60235cab9bf54db5a549655b8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdda63d1fa1093b2c4e5426b4e2344ff266c7cc272b64b60d1f144d3675044e51d6b01440dd40dc2ca31fb8d93980a21781e24ba44802d1623f0455435609415047fe0a8c2d2eb5ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79945b918c4c9ba37a840eb365cc296a531d39872e8271896e9868ac70ed46dc9bc1571ffaff20baeea6811b22c11ade8671ea57f292fd2b0d3c44cee972d9314295091ed6bc5e71;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4caca6085707daafedd0ceecb943ec85c378ca50dee6c72771aa93945647edb3803319675c9af79a913e99dbf646776bea23b1dc0bad57ed9065901aa0eefdebde295f696a2e12ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c07217c45480785b503d97d00577ed21dd48046a1aacbd2864911c2a79703c689c01ec0e07edaf26fa6f8754d798c769b2c84a756bfb1680165e4a70914b17a5f12ed68bbd8a877;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h656a89d200a07fc99d423b22e13b75da01479ab099f5570ebcaf3c8b5d449ceb926f0ba3af8ee544c0a83f87c694a0df8547882e0c184390f4f85ebbde5005d7ea1ad51e59f10988;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18eadfdd115441da180d5c91a85d7c9773d3570debcc375d55b55375c781d9437bf02c8f3cde7db9132c020ba2c9c843b4aef5cd821682f54ccc173c77e4e65bb8b3bc33c1262650;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3388fff4d8cb4ffd47780fd875195f19a4d96ff5301009e75dccbf464c35f01c0338122c126dbcbc3cbd7f1f619e3b705347f03874e325d2512cf47ddb7f1d2fa49706253657b636;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3193bfa814aae06263c6106c242d8e57a3722f50472bd647f96e8e28720915a6e626184265e0b9b3b8ceefcb28f00fbb2b107df3ef1c20c6be2901567c2d62fcd71fe37a6664b1e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hef72e47a6efafdf638f952439a70eb154d4e04853a668cd747b5662840a07bee404fdf4474267aa3ad551787550c1d86aec021309bb7569ee21f90fff6ed0f46aa897397c1c4fb27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h204aede6f28f59a58c64a1c7d07a4d3c80a206649afd555a391d92fc00aa41069a7b91bb1fdad1e357919fff8f14603617f1e39969b8e93c73e05f3296556af5f12ef3f17b41c038;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h231ab6ea9278035318c73379a23245133a8e2b289aed44e89e2504b5f216bcd6c4892940ec8c81ae32486f06563bb295f8c7695ad76ef3aa8bd292d7fd916b22592d40eadc445e44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbcaf3c304b0af2ccc12e7f6e0c751b686625434792a04a7d45a04572cc915c60dfc9ff6ee7f4d5d077e1d6880a0feae0caa0b22bcea5dd551790726c55fa780573a7bc9d852f7df7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7449c24a1c8af07edfd5f07a51a94f146806725cfdfc7716ff7b5e62f92548dbee5b714d541876cc75159fa0c8f77359a76a9cc1c2ec310b9fb610c213c32ad683f073a30e7286a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c84c869493bf0960c0563388c17c7704273871baba326127d5cd028729f6f9a54f476367f9311e53e48d399703c204a2b6eabf03d88c510c899ad39a2d841567f95c9d5d15533f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41b84e81f020009524e4719b2e57be845cf0cd317c434cd50e19f7271740ad94434b0687e0a90efe775d08b12a563c163ac4c5bb4980c9af015d6bea33d129b5f61ed1c8a17752d7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fd7728b34b391204b4b4a27ed8348cd7b0aed5370059f5c62f367d015efa58cb5b97fabd5b8971fd1ce9b63b59c13cf4d1264c9c48aac4c00358286815626612d3ff10a6dbef5d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7eb5adcde5179acc0e6c7d8f50891a981a416726ecb1c036f57dc5e21171b55ddc070e863c10e873544b27207bb1c10e29d3ecdf75737b8644ea5387e523d2055340d0946f59d09;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c2541d50afa3b05530eebdc44bf87717f3c5fa4e0cedbea358df783e7ab828eee169c9778a57bc822839cc42bb40b4d7d8a093d937654eb756048217933b8707845e649126c250c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a53c31679b1642da55b5c3196c3a10e53a15020c03f4584c8b907f8ed2e5b4082a5e816d1e5ece1e7a845dde560aa75792f7afe7f258976cf23b38618f3f4151bb60a74149367b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h663e18791b4e112b1882506db948d7441dcc3377ca0fca24c1734bfd1ec85787a32e02e753717a2c9ec0fa9087f351694b7f9bffdac5d0ecc42728a200fcaab636e4a7be9c27329b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he387311c3703c1eddc77026a689af1c3d91568dfa4ce3821ac482ec14953edd4ce1566e62007015481ee427d4484e60383e42d04e1d87ade02265d747ca7ba2b8713b2d1b181c1b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc75f2d65b3a0821410cc7a203b9bc2b84c1d51970fd507b60a48c843c15c33a92a80abc881873168da5a49b599fbe08f3d77247ab70fc12dac40d84d8cd7e8424005ee559239c8f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82391d9f3baf4f1aaa43625dc50af0e83b4a8347c454c25e0fb50ffc51c0c52b90fa74529b01f5ace4e0ece0ad0d1e393d6d881857c5ab549e2b3aefb2dcf6b22d73cc89701480b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haaaf676836f2d16f65d9a16a6bab917a5e5ddfc7d2a3f4b7e2a332d78781b8c1e6c7326a27f414ed3e8ac95e26d08d865b0a9c1405a681c1fdca69afda6821c8015feb789052cc22;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b390c16c77c5c5e91c71ff7e5b6c7e3284c7602368a710d2435b8a91b011d1ad14e3d51bbc54d9f0466c6ea12aac3ed723dfb81c84ce176a42db32356aeea53e09d74173aa4d590;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5b873e1bb60780f9431d6c6f8c5a0e214b3fdb2e00f3565ca6292d28b8834ebfaaa2ac0589685adaef1bbcf07ab9b532885d6d947910360a60a98b9fd83388df082dd854b6d01c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56972295cb3a675cfa08287c02173bcd0f330534cbc76ce0d5f64d0d5dbd71c196412653cd1c41912a55d7a09de1ed64cec1c1fd805dd59887ec00978e9a8c760fe69b63c5ce40de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h962adb1adf5e67d51bbffdc1c8e207ebe7da1236bf8db68b49fef90ac6ffde6e4ca7c7cbc8f283d60b2de1cb685aa6f96d0538730025d7281e428a0f674760a2da12c6f15235da09;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63d605161ede1663be9f353981e44a67903ba23c73f55200794e0cc5ba23a37d2bf6bb917dd9e8faae668afd2b18e8665720d64605d568b2ddce6bd9833e34ca73560cdd7cd96c6a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56d2cf91905d0fbc4a3f3fe6d16a67723f9ce1a9e6f6e6ffbf23229f3d42f98520274199f2859757938617d28bfbe9cee2e988ad1d34205ee2e32e57b1f38354fdc151183873f02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h329311134e702ad1582aa753ce829e5efaa70bd2d24d5c739f2528561e3deeb5b0aa73b0584308d088b6b406972832e7d5602c34431fb1cddebf9a0008230cbb0788814b636f40a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91b168c4dfe62e49ee31079155a73b9d2b56f0ccd72f8df90bdc388c5eb519c993e03a7739280710653b8aa503dcda2c8a87ecef2b06446929cb710ad6718718893b4d29449e2207;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa145881fb109fcd7c8c1bd224060fa4e04e25ba4190048c5d63db975fe4f9dab459087b3f2c1bc0e771e2737515afbb0b8bb30c05032cbc78bbafe2b79f87100584c7db7575344d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40bdd86c850908abd90d3d5f4728c996453f4a706cb2a746024f62686097f61b7e6c840288eb93b2b0b0e5f8a4a31267a332cb89f3327b0464d6d640621080e297db113cf16f8d9e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47b876c42b89391818ff949c24d8732d517e2e03777ffb9aff395e514e4570d94d9461bee9129c7dd81fda06da5e2360f73832d2d4e1c1ea079e297a21b7915750f980bfb38ca986;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95899d224fc0949ead06737c158a1292d6fb9901f288ce6b9faa3adaa805ba38dd1354e34ea1253649eb5467da0ffdbb00dd3a73a3f093689bd4a6341ee28ab9a4ebb5f126adc0f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33318918045de806bb60ae9cbd84fbd88429c9fc27c6198512c6566610fdd9df85f3dba7309fcc942757494925c08487bfa9d91035999bfe73173f3790e6e700c550b355e7c7bbd6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91e0b26f55a553981635644cb6f948d430a1325fd6a4825b140e2ffcbe1e603c0f0e7939ca004a3ff9144895d2b78cd544da23ec7b9a0e4c2dfacfccfde24a8f6ddb25047564b2e9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c9a115d4756329516943f31e34bc16fa13880f8386858e848cdbc769b9221883c707cac6da784ab64effee1d597d503b2a7d0c63081f434616010194ff942e9a7b17cf36bbbeec5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb31960063ed1778a3be53d3ff49665e7ecd959c4c6d5f7ff46f36ae53b31543dc98746762dc2f7e618f13e5485089f1f1807a48ce148b3a2af34ca1970e7ec8c603f32c04fbd2006;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8eba681e02a6db2919d903a01f3a00b648517a4af96450e488dd3dc72866995508b1b3d7a0f9a35581566198c8ce6f32bad60cef88fe57affd7ec13aa31022d3c2c87e4e757e1024;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7253c4ec7e12fd164ea566c9813e1e44b45b4937eecbaccfc69695899ca053b2efacc7e56fc93bf4f29255ea9cc5d0f651f70a7a8bd39592e7bd58c574af004fcc11c5ccddef3cf4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde63218f428be7bbc698c41e685be12044e7d892f9281c1bc2fc716fc503a4755cbdd90d4671037f7da52efeb6047b1603e51824180c4fbb74d718a29fa04854d863ed7d2dbfb6cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcaa5ca9e33e1574c1f0c0370804e7856540bbf8d85f40bb870b291683c19128ce8ad8053c4fa3a29dc1583776bf054d0adf8d16db44ef51d2092e6a1f33450987aec54a861c4f73a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0a40b513099654781b3074d84ff70611baf331cd414edbc057c276eb246330a4936d3adf96ef4c07bb6783560a7a6de3b42b6614a6a4be6e9e28884055a81e4833a95fd3f89c6fd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc41a32ca366e9520e60da2179c51393f7502b54e1c95953d881e4caa62e8fc749221453a581adda50cd1afce6380740d753c5ae65cd5d4c66cf72a1c5007dc6d1f0c2e5df3ef49c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc22d5a34f766f030a3a9cc9d1b36df4fb78e557b793878f199e3819ee06a62a04d54456eb07c7bf821029c48f692e5c88a417d3f622e78fc1b72c648472ab79725b6ed01b021458c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h543ae0119cc53bbd0889aaa896b48215db483f7a539d4447341af11ab85b6916e6b1730c9ec645e810fbee5e51be6b744cd3abafbb1d93e1e7e29c7f32e0d939edb65703f5485406;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6f02d21a7aa5a217cbd63bb5bb2e1a27695cc1bf7e54218fc8309a48406299d13478ab9a3eacf592b7eb19d454f4fa5c42498d6ff6961bf49d4c18b762071557c15aea6bac7536a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6207bd02c8b58fc1702da5e2a30ce6d50a05dd8bac7dab796b137933bb10a28f54dc86a9d0d8f006d3410aff607035bfaf3c9bbff50f00968737e9843752c685e77d9a831513bf23;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15686a22062935bcd2777b4cbf8ac219c7663744baf3fe4975e4967eb6d2def98b915438f629295135a725c7b40b9bcc64a67c5f3ac24a3b2a3dbd61d4eace4ac8c2ab1e3df7dd32;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c621f27a8d43daa32df5a47a3a3f18541bab2f9e9a172c40c1071637b5e75b59f527540314a980be69d9b4f18afa6ced024c1c809ebf7c0548ba315e1277aaf222639139b820c65;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1fc0bfce8a113d34426f651dbff1b366769cc16fd89dfd8a751f5657a1d8c205458ffcfb0cda17f1b93a7f478c74a3ff1a2a1fd016be8ee2a66ca36a3a32df82e14d0de66cecd652;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14ad4175ed5b6f291e8b70056454862beac933f4dc29d29d5be8aabfa636a346067a6bd4bbc702b6daf1debb874ef88a2b8f6f5ee5a2cc11523db2702eeb634951eeb06fdc12f7ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3052683976bf846da4f45a8c0f48b4a76688cbbdecfc2f65b1d7baf48b0dd91135f596c016cd3d8d7bb8eda699afa9bdee80408a1be77e50b42ce4e758915d308a86eef6a7ee0bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8165dfa36692567bc623f82b3c4cd65bf87d873be0d78924544a8dec5ba35a5485d19bfd0730f72180cda8df0d2c585eb22b535818b4f4a58cc2ac8b21d539431f2e75def11f0ee9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0398edb662139ef90d6bd0b8ae486bd0d21c7fb9e2962dda0986f8d71b99b744bc563b6d317ad546b20ce404936f3b96153137acc2d25b5fdd2e67c30ee36763a98a58c07f59c1d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hafb402227db634277430f089e65fd8af5aa651c5b327859d2f65cb89fb258fa9b102776815195262db8d3fbbf78758023e96fdb9e851953a97593bc878c83c427d012a346585e7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda13b3074c92cbe638f396f014a013a39b7982fda0bf23729e6a0004d1f5e0c650a546cbee147747a0e61a53a5a2cc29871f1334f23731c7fc4fdf779447097621d223e0b319eb20;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec55f8a22bcdda4c83c3e543b54880fc9c4750b725c4e1631d7e8c6655c2d70ceaf7fdca1d4da5e6e910faf5d836e6761c149d3885e390418e540b248efcbb03adfaf0b64d0e6a05;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbe9ebf42466f6b78f34c14731dcc4cf65e3ba1d11c522d9c58c8c83e19364729ca507a078cb4523f9faded43b5390b1cc09bc58cf3607c4fb0e7b173c649a918dca47ef6ebd7f36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf6b6e8a699d419d5a0ac24a8d2e548d0fe51541590ee8239b1bc5f3e7dc349a514800bd1de8842b505b51a10726dd656250f913dd0466e2a773e18009893c2a92d4a2bb584c3dcc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7cbcba1ce991a0c96e09ace93c2d4193d4670edef53233f5e2bd1d5b61b371f5747ea09d57ef9e1b27a72b38b8db991a4937a6a10a99b53a62c28cde0197b981922cffb8a7951b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e7945c6b37bb2215281e9502c298d92c0564b481b509c439991378bf53b1691819cec90674c75ae4034f6bcfeaad9544144f2cd5acf833aa51e6e09a12a68516514d3353d97fc43;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fdbb319a2686a1595ef95246c92c2ccf1a622b42bf773d16e8963c4a6172d8a96d5e3d4a7612f3982c45db3fa010f17968b2d3c731c284059b5b14d6e6ee2357683cf4614193482;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8dae490b637e5edadce7a0f58546c4396669e3ef28881329c9da17dbfea841f84ed85fb973723b35bf3bf05238e19183c08cb0f68551f872fecb5a57651a6d09fa16b6c973380a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h333a864625b19a04f304ccea70dfa84c76998b2af16a32ad5eae28dcd8f22c42f9b01d8010300e19cae1b82971df584f2474b58092013d058ee8c96da44e3fc0d3ef46e25d6362ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60a8f091f26217f579b9e9eb63c4e0b9611e239dd55b045460b83c070b6f2a910e98c972125983eb872ec22ccb608d88f033d3a2686f37e6542668c8c20e4e3f4273cced014d7f9e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a1968432f824d7338e4f66bbccf39972184141bc0bcb10cce8b3e6a9c973b643c55d13f283b3e926df66926ac936675395c89dc02207fa2dc24db7d9630d27eca0f63f0a0d259f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ffe23e11414cdd4115146b22cab32e0d6b22f90a95905aab80cd882abfc29ea55895fc557ae63ca2625001e57f149c049dbded9392de55afac49fa124f715b8113698b7a9580227;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedc0f46670b3477ba06cc0fabc419647a9034732f315cc7bacc408da5ea2057084f03b09f91e45a6f97e64ce00bcdaae6b7997a4b9e895931df3b46ec0e7eca0375ed1f08ff2b9f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52b09168e75688a491fa8ec289bfe2c8a088cb361e18ca88f303fe865209ffae062763fcc65aab135270c4ab22f04d766dc439ff806e1c065b86f8c1701dfef3edfb5aec74520cff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4a05bf58969533a9c03bdd92bad2ad9b8ce5e62b94fc465caee3d533c62b6245e3ee368f47e1cd1e10459415359194a337c8184c7e6d0a51a06800931693e3ee62ce34f1b13074b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7895647098c31963bf33bb7811a391aba42cd1313449cf21b5dc3b90d138266d4cf40b3e4a2f26c1b39fed00bbe60b38a0ef83b2cbcc33663da228077ac633e91720073376e579d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27f32fa7e1617560fd305b1b97857a97f31440c357c36339e346b4bf55732df5d2faf8069221091f0d3e44394bb75e48c8033440fc6883c40333917205c5441ffff29a905b4f695b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cf0d1630d3b13f333ba53dab2ef2f0b21069ce4cc0f739828c1a33c17bb03a38d53c5c441953ea14afb506d69c75bfe733e1526463480e7380ca5d540ca2bef8053525fe0496a0d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2266c9c262027af8cf2f864dbf1e0f325c711be7701ae6c9f46fbcd41274b041a490412d2f608055f88617a92c0e4e543a0858b3a13118fb7bbad13f85b7fa17e19bf123e9857007;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb093dff2476de9fb188b7987dbdd88db9e1b05b3cf459c9d5b6c5605120d76fcfd4ffb18d4c8aa7dfc0afa6f8a9ee893ea91b6c117b66ba2a7f60d9fdc1790a943d300aeb5904ecb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h677df5f9c68e84681baa8f16f81d7f9764390662c7df7be9574442f31845a2bbc0461c5449fd8f54b0a79ac02097482690135e5cf7d0dc7ee8153c6a661bdb7bd751798ec5f70bdd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d5d800beab530a96c7f5f5b39379eac75d35544028f5cf0b2db533bb874739bf6e5685a8bf583dd00d1fd4fee06e6d4565eeddee550280f2d1d33e66d4a6da2043a6ca5e9ca845e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a0bfcf92f458cd4f3b6d3ed315d2a3d9ac19eeeaaeea39ed206a03cf84d02f89bb71b65a9bd287e6852820bb01b6025cf5eccdc1231975b25551c88f1fafe3ebc0b4d703d04a930;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e158bb8b3d0a6dec253cdbf83a079a0e284aa3e6c2a9b59abdc5e0505a0387b0ae8bd84a9b172611a4628a0ba0235b36f0d09c38becba2d1d416891500cc1cd6855a75c1b901074;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cf37e3b55e7d69c01993c503114fc540e50724130744a078649e3f111569f5cac80b0ca85b48f76b03cd3fcba1679309dc1c80d7d08c89cef3ad5bcba0b1ee2fe6d5008f72b104c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc7d79f53ed4dcd8bc04cffb3c3334780830ef4ee0a3c11d68100d242ea49e92499f69dc5cf08aa3b1e8d70d11c35b766c4c8534dd072f09ca097c343adf1c6d5e056d340574d39b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80d97f4ce7ef29f7402e2c1e7faa1a4372336d95cb779f2ee6ee36cb3a0be3f63b80c9881615ded3ee6a4a8d46e99a510466174fab843eacd4105e9d8c5993db3e68ae20e406eb67;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cf8166db36b1111815e32188f11db956b2e405cf0cfd1ad7c4c73b299d11ba23e71d955b37c02b6c8e0f0f51494b63a2aafed5c4f47e36d0438c9fabd9be192a3f1aa673bb6bf1a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15d627e4593d1431781837955849a3be6f114cc13e754b538a72ae0422e1142898050b89c7742558088bc9eb9559163f68be14c17c88d23174235e63985a7756b97da415db3bbcfb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a5a7adf7723079123cc062b50175dd83383ca3babbd1bdf962f7dd3a8bc9ebf2146bb3861dc2ff036bb0a0fd10e9790a362ea7fb3c9faab78398bece6e3a7d5867018b05527526;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52fdd018f9d04695fa1ff584cc96b47d58f0e090644a042d7c270edf34a975f2ef0cd27f13bb06d13ca376394cb9effbe5330cb5819e1975c9dbb5e3ccb285ef45cc3ca498b3d596;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a5068921de47790eac137ccaa1d47bf96375ecee71273302806e662be1c27579a6820f983b89f46672cddba963ce39bd5f2db5c0bafa01261eda9a5e792ee6c5fde580456a3ad55;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6531ee253daf18bd818f47c7c7404c8ad44cc9e4027f82682ad108566dcf321bfe50d4b7c10bff650c05a764d9fd2fc0d5835d366f51c970579d1a53781780fec25b58ac0fc24b52;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f0a676104413a7356deff3a41bfeab599f03eb77f428a15a07b2e4e4c36da42af0686720f7852febb388467a4a8ab02d85b7e3fc2940eabec2054a157d28d0d2572ea82693c08a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24262db50ac089838ab9b7de925ac9b2f820d060e9c37b9ab12fbad83f9ffd6be646444ac08d12c3e343c3b9da85b2bab3d7b8477ae97589e4726170cf2c2c1edf04f4e23b34ca83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6318a84428e21c36ba7843147b9545a0cf36c92f3975a1483a52877d429a6271a8153679913ae31604db4b6740b2c23c9de50bcc0998f76412ac636828809b4300eef386ce4d2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3152b9ca553281c075dc00ed1a12c865a537d985cf92d53a906df3be237fbea2f834eae293703f852134f21da719fca172331843bb42ce1b1a8b5f8bf896b8614fbf512f99577ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7fe368f7ec49d6189713551baf864f8fdf0b9b3d7106050236c6646fc39c0f20d86acf201cda632f3a9ca6356980ce9ac980af30c0534edc9312ea73c27899ace83f76ab20ee04a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h407b478c810a077ed5173ac1fbc4d9f6c55f60e62b211be537d98f4b46384295e03485ba5adf7589454e8d1066e3f776eed7fe50492f8e9012862e3326aa1faff2aea6b542f779a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2503968deaaf51d569d27945ff7271ddf349afe73865d589c09b4313b00d30ef96f7c7d82d455b03f9d27825f5842b1e06fbe92fd68804dd04674ccfdc8632963f2d6b19cf318b80;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6af9e06ce783876dcc165cc4b3f526894a3b0ada6616297790d3daaebef3d613dbe79cb3a12a4be1065c269c0df7dde9a33d8ad5da68592b0a0243befe8d944f8a8fbf2c09cb427b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had6a389d7cebe042844684795046da4a2600870fb413cc982e951d22e8c248439bc41b76f871da61512c8cb64c67f0054a055446810577ed8512901b97a5b240eb0ee83e8c4f3fc9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8ec8c42205d897671e1eecadb6b3267534b4942aa05cb650bcc799f370f23bdfbbec3a1afb6830f7e71dc547078a257b7e767dd4825e066b36fedea6c22ffec7ca2cc58fc32c15b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c473353901397e8ae668e99a2f1dd84efb654257748090d9873618daf8f7aebdbc2b03d93908d37cdfca1a0947e01002d67526011869d5180d248f55b0ef62c4e28f57ec1a0de1e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h801072f0c6b4faf146309fc14e0734fa59bd4d6695951f221fc05bf6281d2f4d19406d2fb00af3a54ce9e40982dde11826ec879553666d4c63256df1fe0cbdfb6f93c6ad1f078b80;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5f481cb99cd40e4d0305e094d86e245566be1b17be97d732314d764d757f4144a2b8e34db7040439fab0da06fd8958593aac6ca2891789c7c18633e029ca7b8d95ee8f0db9a7ddb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34d44545956b86ca81553b98caaeef051924d3bd840aa2c1d8b47409479a7720fbf8d17a9d0154ffb9453d933663b8dd862a13a10ccce0add18cd02eeb5d99020244b6bc24bb2491;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f942f8d393963ff67b37396123e91c52ddd776af76cebaa3e68078f427d266df70439ace4d8d57a03365d76955c3c7ef340cc29110e5c649d96edbb56a2bd908c0726d637a9453b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60bb8e77df84370180f7c75308ec6c5346ba1dd7a511b881dad40b624974cf832c0dd3df3e1099514f7e5dca7e6730029315d0a73b72c26d923366804fd44ab092cd4114c7e2650c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2df3aa61c7ccb6a268963923535dc562de44eae7852e83342ed6be6a1503cbfe68c79cbe3fda2cf5f47f3c199c1db10f696b0b8fde5306da4a536a66daf592f8243ad595b5cbf773;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee9c83c7877fec2c28ae143c1967e77078b73971e64dea0457be0f50c98dea0b333dc1b8c3778b77b32dabd0b5bab43d2e81e596386341f33d4569031ca92e9d5f576ec2f37458b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd71e023d6abd6f9cd1a88e551de945af4e1d1b021ec091c065e7da10114ca357c05e2696b48eadbc3d9b5b8c7f47ec0f07d5d605fb9ebfec35a50afebc6d74f01dacce3a42f2927a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10bbbb8d9d754be9c67a57075bc5d5e84ca83d041023d124de81b3ca586cc74b90b3d6cc5e59e8897d38064559717328d7d63d7f2c4d7105c4c39b3bd55fb5e09a568bf448096f0e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d5592676e0e1af6fb76e842f50a0cf0203a1b046b7c429d13484cc5d5d505f39ec7817248d9d760078781e9446172b64b65c4c567478706b8f23c173b1d724de44391454cca3459;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h234ffc26fe07537859eac51000f43923e154504b09f86a5fa8e1b27c12338ca3766555d4474e65c7c91b9a38e5fddea81b477ee41539338e31418b629044ef52fddaee7f7346cf7b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heda6af00a282f40d5d981086b13c695d05bd130b4d9c69c8d561add7387a94e6fcafde234df791cf59cd7fef4f506cf31e99715861c2d3bda63cda341eadce1ea9071d81945ca41f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b55b174f1123a9b34475dbbdfed5df2b0c646c0ce117014363e0c8f65e39afb3e520592a318a206684b62dafa11e6faddea44c56faf345a7e87f9de47b79b72f3bc79f35c9a10de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8360f1cdea0d2455e18fb76bb7439afedc9ed45bf10d3a8dd2d7a4772af4ab6819c08475400bd06688e46a985201b90403e2eee7ae6e8ff91585ae88c16b1230e26e9c49ee9b2b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba697c05b19dbdc95291a6a1eb994f8db2da61f5e774950bf1f0519c6dedef5370e7e5d637465e1bd476aed5e3ca428b20df2b6cf86801643fba10d8bbde7d77287b62b493178ca0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h269a9e7e882e96932bbd24307d2d5240c473f4c5f362c506b867424b5fe6cbca54f46641ae6833544ebbec4eff89779ff800fd8b37e58726ebb90ebb2c4badd72ca5ca1ffdf175f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb690faf802db1eb7a53697cadcb7a8a3ca6214e2b0e2507aa71e99d9c8287ef82dfc16ba6c05166815622befe7812790a8208edf585d3b1418cb46a5229b0c8104ae7cc5e3d1bedf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcfcc6799cca05dd433d4a09f9caf3cc25c9a7960c826943bc2750fbdd74fd4933ab490e045784aea246aef1ea294847296b944351363bab83ae5f03c2f7b1890a718f2cd6c09e59;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb115d2f72d3e288d3a2a9c14d05eae994447c09b38214925f0ea0de6c5f33ff69d7515afcc87e9536a7136d73810a74d24f0cb8d520cf13962eb1c9ae5e70eb2e4e352abbf397058;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9fa62ec0d211a1bab0e2e110b2bb1fe9f8bed599618660e2fe0a26e20f2c98fbe9056d79701e79a73c75508139c7afbcc1a5fe9455c3f92f8d790cfc4dc01262ca05dd6522b77bcd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dda533417daf70c3dc09b03748066e2e24cea9cb3ebd417796c3266fd3ef29fb3d99266756073f3b611513422da3eaaf8c2cbe53e15ae061360f5d23c2a4c859c8a38f6002fbe9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1ef3d2bb4e951ffc8c1b4e472bc626633c6aae7bfef4d693aecde99100f73c68e9b99890675af0ac3fa9737f43c013eacc6bf771088405fa092a00efc91918faffdc90a763f70f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee08d3b431c2cce206dccb0a4cc05a3cfc5b5838ce1e1b67ab77ac7d790b5d24f625dbc6bc7dc5c1236d5b3eadd11ab2228899b17f0d8262aa42774c7f64f88174b15958e082930e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcee055402014452c92edbaa0b943e8a86451468c484ac8514e8b1801f0e2a93c9f7d15c9fa303a8837147feadb19b76000ec6cc0b9dc0ed18b26551efe8d4807b46cabeca2ac3397;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70db7c69b716b3806c3577cb80b6afafeae884f4ab876f39e3401d55da23e598fc2c444c3ed497dc179738ed6f081f7b3fd7c725904718a8fad285d324ff0abfe50817e452a1db24;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h675b4948c7e5dfa3c4966204026a42349ba52d1efd2654faeea1564e16f9acb61b25ceed23914354c8203dacaf1226f29fe915c8920e862e9171b3e293c018b9914f3c4ac620a52e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42952228e995615c7a13ccd8681338179352bbbc061d73c58d07c5012ebfde9677eebc509ea864ee4e4e21c058d213f1f8bc5432d3f405c8f67df1d7427dbeaa308cb156166f7b09;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bab2efee26e57873d69bec46cf02c3c8212c79b520c5ad31735cb1c2d42921c57152244ca767ab54009bafbf5cbd295b85f47f5eb123139f17139d700c3a9870c0064f847157b51;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h969f9d2fb220467d179ee50786867065258593b3a9edaa7e56515a3fbc214dee85b747c29080204e792df8aeba1005c6f154da1a2de687b41eaec7c903a3387cfcdccd732e52b506;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43ecd05a989ee1eb8d1989273afcc986bce43da9042cbe9c5c0303f41b0e32e95c5a8ad1f64a44ce10304b703ab9dde183e79c0ddf83dc42f10da526e4c6fd7947a626485b7bc3ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79ca7fda5a0cc13ae25b44719f21f16d47e6e572207b28f375d82349b7be7f430b17a64e281cf1087563c47efcf6a0c513b7c5649641a3286529251a321a0833873e1278d05fccc9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b864344efae0e5bb396306cce2fb3031261521275e22ff34233a8b71a095de42a1fb4f2bd6e98df655fb1a65263ff46e60a39a4fce7983a5143727eddb3d932cdf73bbd61e908ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb5064a5036468a208d58a5ce493bfee869ec43474e8a492914de159476b1a359f2e1ef1480f3bf9cb62b4efe21493146ff5a64f38ced1d8f950987ea5053de5a37e4720993d0af0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56e6a5c9b88cbb2cc8ecf8a21afcfa55dc2679cfd612a6858fea40a1af2ef226257213381c6f8638bb33fd5d02588d32f86374c8d91c06c09024c7597e85ce1fa07064c6007325db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd0dc0597bca2ec4e882f53309bec724eb1ebca418b0cd7068bee94540b012a8d88d6c695c38633de09d5f020efb23dfc967a2fe5b3daff1ea5e8c3e37f169e41aed56f1805ab82f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc41d075330ab036058b14a7d004f3e8c6110e54f9361c53cfc6f5a704d118a7217bf5fc06761967578fe2ac416853c928bee5b88351e951ce1f6de176624c8814d904c304dae9586;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd38c96895b3e2cf4b9e5445116a44d78fa023b685aede91395e87cb355b8a70bf6e69b0968ae3758247d58c68e397d7a3b43680bf906b152c49c1a3d1da8e53432caacaeede87132;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b73249aadcfe7b76c302aca0a1645424f7e89c03b81b9a3361b5b9b77c6f6d0fd129b72463477fbabc181ce1f67fdc11126180eb97da1b0a3a3af76ff97b2c6a05cddbe7704a7f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a58463c3bd52cf050c012fbb6dd4c35cda6354efc0ad1e5d4a02fc5a96e44d01bab15eb9ae021c7132169ad3ffea4d3ada944f98d46d8b65f4047400f4c6e5ef65a6f6d1780788b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5dfa98a133457869fc975fe902ebffce8d428afda55b348fdda4934ef65f50bd99d40d8e38e688a78714018409d26cff565dd4dae493b594172508c14c6503113d987c520f32e2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4f6f6f307067ac4420dcd2a6d7dbac01e65f5d0d1949039a18b5d25c58b3a77ceddc39122a8008c7613b19503711ac06d6d8d03980a6c91626d107adc89913016e385ce3cb47d8a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c3ace883631e304bfc636ee410675702ceed3a8b646a67b80ecbea49c7e6f478c724994016d9caf4536db07ded57bc971316eccb90cd76058e7c4740af23e274b17ea3b3c67d86b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33e10db3a47025b68f2998d424d8ba77b6e082e20b94f0c4e9f3964ca5e20fb22d9b4393fcf42823ed7e7ede83871b23420e4a7247975598682f152cba0e447fdbb11322fef6509f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5c3d0944bd7adc605a846bb65197213ec029439820da8d1fc0039c788dc6d39d090799cc044a27c83e208058ce50cd885d8d3355c7748bcf2ff9b3e4aacc6f69d2c9fa721c47a69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h448364b869f6ec0cde49110f33984a3167f8a583b7ece4ea8cec6db0d1b6155ee54223bcbbf6014e2f4723116015fb59d26fab591d8e633ad6eb93075be12f5816e887d1d3c507b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19d54082000787797fe9f8c9ce9e04cecf532cc74264ad1a195f16a7f9928a6b747259f11611fdcdde10b66488285c2bc62c1916bc432f10a23702710cd9621dd6dc1810ea60206d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc099b9633d8676a6656cf07321d9473f6698a1c85bd982af3acf6c2ab5ab1c95b63436a9406d429d6ba73255c8b0c3757ffb508d5eb56add1807f09458b6536ff8159a8f8eecdac4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he82a12ed4810249196b3497f7b22d15776af1dbbf95a9be0c8f407975bb8390eb736c883502dcbc6b10fdbe19be96ae52a4643c75a8743f07d6f2c843e210a3ebc804b3ef5d9dccc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3b32041010ba3cfc1836a1602aa4c0d649d1e23e7bf8f6688aeedc7e044ca872a63ad2d87684a845fe6160cc1fc982f1a4481a09f305c4034929026332543a3625614c357817ab1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f7c36e6e397623510c3054c685566178ab9da6711b52892fe4b5512fb0a9398f4e55da5eec537e4b18145d019de633db3c9ca32ac253ddc5bfbf5647101a7d2b0aec5db732135db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h137b63dfa04469d7d7de533e7c133200fab4009726efdb2765ddd9960badd65a2b9a91a761d623744f1d7f031e0c5805840d59643b8329bd8edda310882335c8a4192d7502b7ee60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8cb11691c03f3c6559417b3fe682eb6a213ddc32d7811c9e7a4882c01992745d9b81bd9cddab92132420a655fec7ebccc7250189db0f13aa8c11ae339d49bc7fe5fc31694d810ee8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76ecfd7e46ed0cb5dbfa848ae9504d538746d591ee4e1d0e8326ca2f644f14307e86411a7f5489d42754d04c03a52a5cd1ef6c35cefee96e840175ab0647294757fa6d44faf8dfc3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc97e351e5e688fe0096559aeca0c526c07a26f447739c5e245e8ebcb4462a535442bc779b932ab92f15e4d31fbe3c60e52491a5856a7125c197355cb3462128c59793cb8d342db67;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbad098cc62e73816ea5e6ce0cd8580747e6b1aaca6a485d50f36ffe7d139ac57230c034442d57eb78fef8e041ab02ee52efaca7a7053f4239abde7956f798c3a7201f5227caf2ee7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he173f6352cc201dd8e40d7434361ac820b571985b048a802eda56b05c39a1c0829ee58aa5200a24c3aafd8dad23bc5c41228b522020808af10bc59079cb2ce38838a68472c7bcdee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc263eac669f180227a6948c6e80b78e97670705b3e821b0fd42e1f3cbae075c65f7acb5fd3794a455f0c938f2ed651e3714ca0c28be2d12868df30c59bfc03b842ac9f5c1b9a4aa6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7dcdea44cbb73ac7e0337aa7669e8c8cc5bca3b4b46e4fd1f18bb330ce67350eaa529cf4537c60465ab451e582c9bc0dbb1988e4054c6cd48fa1b1b211dacb5dde18a9ec68331f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha90c8f1c62664c81f9112df33d4775b08dd4fea3c02f7fbdabbba01fe860d6d8b92752dba943c48cb30ebd4dbf75dd22a7eb64b152fbd8134d94e142552413e58266b7782834308b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b6fb23d3944ac3752abc0d1f03d56339afc17b15afa9dbeae55793f822fd46fdf912a14e98987945b7b151ee48f9de7ef0568e6b4af9f11289babc0abbbc38b0308ecfb6a72731f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h576ad4865da5b3198200a9daca712202bd434852dbc02fe54fc7d041300cd9064a1148a0e819b380cb16d2a0471f56436bce34cb062d8a39fd5ea1a0cb4dd562b42534df37f38948;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae12cca126a717bbba5221f619456fcb626971cbe37bcfc691fc44fa77e0c90338071901c18ce91847d9b9f214d567cad43c258bf71ef4b1d79f916371739e157a074f51bfb0e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87bbfd8df61eeecd2ad949589bfa67ffe0e574f98158ec389726ea7f6f90a68115d05874e7500db3d33223bb0442a098b0d7de58954e49eb5de1c095d2028a05cdde5a166bdcfc68;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3c08f9ec6ff28b45b83ba18efea86fda5096c0342ee470301edfcd38754829b4998c959e1888171396c81c4572d8185cf0544654600c834845b93b00d8f13922cbd038e95a77613;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd89c4e94248c92cad6045f5dc2807879942f2f345a617bf6d93f314977694dcf376cbfb891c7726babad2ce8132b349765bc493bb470f5ab466274571546823cba14eac307e81377;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4b42233a131d887d84a0e97cde62e50c3a989663b2b9210e7a77f2498b4fd6f57c571c7f487bc7e2f7dfbef2cdb04b29853af2162227a7f324666a05f90adcc13f9c143b02e5c86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4790f20aa6df918476c0e0cba9593ffe139baa46c45d9601b4d9896cbda30a520db15753fc016fd21e21efe012055090515b983060e34733e0c4bab647ec7f65326203ecf497868a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he266ef738807278f4db66b81b6a6b89283395ce5da71d109a23f6de9d2a10e0460bf5d9f61d3d0df4124a9b846d5095f46fb81378ec66b7b4a0d46ccfd553e6e285a5ed407c46c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8b5e377e63d2a9edade0694691514485b765de1b8277eff6cbb6ca0e6f83ca556b57160674fd7920d938635a20c1003719e558eb0516156eb2a5443010c7f8bde916cbcccc17707;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9f84e8a728040b224c3fecc2bc11f09949952bb2150ab07ef5e6977caeac8c5567a21b097de983b89f357ac1c8e611ccbbbecd3620fabcc9a6102982fe108a3038a97eb1aedca47;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bbe62383ef18e643fe87b49c98b6ba90173723fe57bae9b50477acbc0a95a7bbcc9f3696dbbac8d5685c26e57ac05d347ddd3522427fa26f37d15881d2354acad1ab93128a71bf2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd3dc8aca7065daa1f1f5970fde7815e9250290e82425e7ad89a5012e4060eb1cdbf8db96d6c637ffcc5209e1af10ca6912a7de51ebd4c96a514192fa90e4c03865b6dbf330fa273;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fbee043a4af6c5965d91236c6a2e44fceeb5578875114992e4cc7114f33b275ebbe3fecdbdcbed2f74b61f38f8fb8a4f531095d8365bf10a7a52a43c2f0363ca78b5db171427fd5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3caa06749fd110844a4e596420e96796d813105cdf8c895e7edbc57129a04c44040c84d189420b8bf6c4cdc98f9f1bde29b070f85c1dab3a462be167f95a100c75955a3b7c05b420;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb07065ffe15aceeb386f62b2665b68a52edbc85546c071b923436307ea4158ac13dab3f22e537d6faa3d1b7db61d884f19a21925974751d62812df04f01af9a01a687834540b73ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77a4113bd8cce133430ec9c28f4113a1e0fea558f6b683676635dc066a70e78ec65d65e20dffc96b6f9ef917ee0cb78a03a6d1e26b7b7a95fa6f9b3d6074a2c321dddef5a4b14bb6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h878e96fcfc7ea50ecc1e9e982359bb113555e5b44ab15d6d7ebf3d754478cdf4950b909366901834af6acb09cfb209a8b01ebc989d104903ee288a12fb0811b1da374ed42432b386;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71c591a1b6d926c7c7d970d4150a23227c30803efb4e601f29c70b831b0c210ef506efa729b9e612bca14b6946ff45d5c9d5b88b1635e2d4054d596d654d23c49ddc9bd3c7c5980d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfde68660426b88bea85a37d43e8b91c6b78ceccbe22b4896ae6eda73d94dbe8bee8930c90ef864760dfe7c792ddd43c5f41a0cf7fbc79df75c5d79906b6bc688a2ba66ffe7a01a17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h991cf4ee034c76c6b78bcb5662f19a62d7e602df78070738dc6579ce049137c076326bf19a3f9701e1e7f5fd8c3f2cdde941e2874c7755f751c44d1a24b3b1dcb295e04ce4dd4c78;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h598e1386a9994e6f76b2cb9ce57bc0ee9b7d2618202922a66950d75df88ff729fa135db39673d0d0a5bb997e191f111df4e5a2c35256d4b3bb60cef4f9c41f182ea9487bdf8f65f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf8dc418e9b1bcf0b9980b0670a7cd4a783ee72036ddc9bc32da6a76924a831909488e6e02ce18b9614e6f0b184ff93983fb189ce2bb0b4e1e4c194e2254a0808bac323aa9dfed03c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5db067a7d4d6953bb5cfd74fd1e4bcbebab9f61d5eb7bc6e9c8b9ac2ebb62c819e5fa18af2ff3335ddd5ebb74a01a75768fe7788e916999f8a47eb884aaf917c72c52acf935e6e75;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he74628faf8d5d0596561e096795c02c2aeaa1702e127f00ac8163232ca81eb576f5292519577ea5c4fdb5fd32e1d601f80413c66fea892f19b8b1e07eb9bbacad2b3db91ed573fb3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32266674c2596565e8715fb8dd37e6a11842d47aec1790d30627446195338300e334447e1e9ad040c741df0203530ed4098c21bbc1f64ee41d56ae13887e322b107082bb58cf37a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fd6d180ab49721853a9fd6d6ec08f15b4004a67a919bba8761ce5eaeb12c5d10c8b185e8c53bb4f2727c828a13b23bac6cc89d6ea4f038278f29196b8ec3363d60d280f086411fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d09c8864f6a0da09cb4c140ea1aabeffa15bd1c2d8e97374232492f29b75076979bebebdafa586076cc6c7a017fe83c454d9a79859c000b0345f0ada63a29140f260bed3480ff9c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c1f76bc2a32b6b8b4cba06f42adab5265d7daa4a551db810158fabf1f419c241bab2ad2bc35b903580b2c8c389a4315e7f60d60d07ae6965b98a048dc66ed9e95fa19fcf42f25b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbd7d7b362d149fb59bf5e01d716dbcf63ede8329d0fd47e9772524a77a86cb3028826e136ebbe2aa0985900ead22b93d7ddd7a76b3f7f4b453e27e1663bd71535903f29c051aa28;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7767494b95610a843a0d29a026484ff07385d0e69c384ad3fddbbc13347a7bc7f8cd2e57c258406e657f6ce2e4c9f7a3d910d678a00dc9cba5f0957006f1d2c9f5995c5075e05fce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1a821e7ca03878c33fd80a41751dc3835bbc9454de087960e9f636cbcb066f9873cd859a4128325a780f98856017e87d6d2ad0f09df7823ad82704eeb625faff541ba385427ed28;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54c06c675feebe98972a2f87599d3b24c600aac4af96dc00f8435074c3406ad42097393ea6d3b6a91578a45000a32f49e08a5aa443f773d400bac3669e7fe8ff3635f0cd59f3c239;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43770c9b64d682da240fa2dc0a97271b45698296d1eaf84b27a6edcc5c08a89bd206b184b987917524f19fe5b43a8df8f0684b9027635005a65f64958e3f261b879aa3ab7d5b1631;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf6df11ee783a2a08e21a762efb9585157b1f1b98f32670a5330fdb3907b0f1740aa73a503a158ceaa819de5d1f532180df8d06b27ccfff334773764a0aef487b7871a2981302a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc12dda1b51579fac4af3b6327d4f2bfbe940d8b0e65be4f50fe1a7dca575feabee4d0d12771da42843bf8ff15fdd2abd460445945d90ceffbac2e10e2ed907b0d937297137e79d34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c34abd914ef0ebf55c1f631d00ae008d4b089f3dd005d3a2084492d987bd697f381a02fe53d7ceb2845cad0cc35c6a0ea61610308e892c4fdd096b3ce09160320437fc4855a0ea2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82c34823f66095fb0c0a3a3618f01e76cd63c43fd26ed0473ef7a35c7f64677d8dfc7b42358f86ef215fed68d9921e032c211169649a9a09ae295fbdb1979a3af0e011dcd42c993;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78d7163e5f0a7e29ea8ccd453e31399a06779d887c6865981dbb3bff0e860961df047d19ca450466563e42697a6d8171943a3018909163e81a918fb7249745865b871df127a4924e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffd9bdd7706a955a11cb4c0478512f74c1167844bb1317841b00d51fa4a4751284d452d75180de6c10b211384664c1437e2671f99621e7fc43dc48ae12573373622fc6d1eb4413e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ce8fdd9eee8edde5335f7b10a247c17eba3d74f00f26a962cddb4f15ea6836b2454a2d9c5f1e61eb0d4aefee4822a89838ca0ad15f6419bc287c905c0664a6453b222b7e093291e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h879d2573c8caa3cfe6a3319b35c0d2c01c896d58e2db60202c6a146478c3841e2dc0cf79d9ae2ba7b8e76fde7c78675ffc36a16bd15dced251bd152d35f807f486288bc3f38c3bf6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h817e8e22f8c29763057a069cdc0b8df162f4616c538fdda3c742bbb34d667e9d4e19525874a6384bbc11272e0695a7845bb311e8a24467be0ab0d48520ca6abdc47eedc1f02434ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26e4ff5f51ebac0a95830b607c36433a3eb86a6cd330ad2ba6917d3e483e52fa397d55bb339d92d65959c6bcade6e5da676c89a30930d7dfff36ec8f46cbc7ed7f2e0892406a4b33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2b67da84e716b43ae60c73ba6cab50972fa9b829dc4cf719434dd47d4a1e1528af708daa5ab2b7d4c186a44094eceb3839c71561182b24b1c5c7a51db3a596dfeaf17dbee9accb8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8c7cbf201a444086df8ea7a292dc477d743d6d72bbd998d4b92fea2529b1b0375249eefae851f3dc167ac00c50fea01c6b7085fe06d5a7312d24b3ef9220f77525a63c8488ff04b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b5d9cfcc49182ed1202162f364e07259530a3ff9900c3d64be922cfce57808138ab527479a9d68606a5c9bfbd22bbcdf068b0566571e284463077a7d2ba1d60e81c839a1890db0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h520c8570a50a7c26908afc15b5aaade1e132ef202412ed683b299799d0b4fc14428d816aa615ed54cfa49b676642dae14f37a2c0c9b6d9d488e074093db7fb0961773041103abda7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b2653e6826018940e66045a8c1ceb015481906fa9d51bc972e68cbd21d3fe062726cdcb77c6bdd956a32210084e15946902f27f7dc71532f115fa6b8c9ee156901704b6a104ffc4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb10c7f047bae0a30ff05453058ce80114b1f3d3e6eed10e86e61c5a4c6a30cf5094689303883865681739c1c3aa0c97c88eab1a9f32b48d44e8e58d03ad8124308acc5bb1d17e3cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56d26675384c6c8325c905a72663e9b9bbe5c2e523759723c7e4401353883e489d8ba25b3a18e57d0a89d9594405644508d5afd4e4c677740cce4fa007b162c36cdea1cb0a224d19;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa0f0f2050c67ddbfb0a2bbcd9cf5b957a4f3d6d7514d1a45411b81015206dac3b394ffa593d274cb0907230d128ee3e5cd2a6725daf7a3cb1924fb44ed4317b65ae14614fe5531a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9195e9cfb5e56cfd6894f3a526f856ac9edd2df3566041305d80851b0695699e66be20a3f650a59a860a3713b219709fc31b1879498b3be0f0d52351d222458b87a4dd9aa24e8c27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9d759f650a434b7f495acfc4b3ed873693fc1befeb7978adae40ca5a4f6b346651ad1415ab20a2daca5150d703099fd8fb1201ab72664903bcf4fc2a78b460864d5b6dd0fef16ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41082a90c8e540ea7d9fb6da0a3c9ba4dad9567f98c17610c0d40f682bb2c2d52b321ec581aacee71bd9096643e95347c293cb5e369b3f8ca09e23e0421ba8232839dc57ed56258;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fca64d56002f7aeeeb471524c208d7f6c66dadaf296f0734e05a23dfc10d41c00b2ca8e89999a3a063f2e32c721ba5d7bb6c36df047df60f6f10e730b3112f6be2bd586c46360f3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6680a47d0d583986f486e78c3b2069ec7ff86e4a217b55bae0ece541b2883cd06d72c079f9e9980d97bcd46e6031a0ee8a5a59623e7b6032ff7cdb2ea924b0555a188964acf9fd63;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1b6ff039b840a98369e314e70edccc7eddeadcd18fc6b2eedb793854dd627673ef8c294b3d5e9ed24c7601049eb0f8ce1311cb203da1538b070312cbcb9c9df12812e736143f71f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ca719bf651383f603b4d50a6948aeae4571eab8ae5497af11ef6d0bcbb7da8b757c0a5e45fbe56fa0001ef338ac729667fe9af108b499d626d10d5cba358a26114d1b138abf643f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habfcc3f630223a2b59e2b120cfc469188aa517874938dfef4546b68ca2884baad39b434885c1de4be80a32c0981e82f89c94e6e89c16bea0b70cd73ce379bda8a1a962cec17feac2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h522fc9954a979c4586ce80d787659fa452d7c8f47ad26aba1c00f1102b88cc5a263273d8f58cfbfa732397f1d3850778e91bff3ac081f2ed05f6558cfd3a6829b37e69885a0e4437;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90042859ee8b1f916182a5a13176f90df85b02cd13b7d4213732f54b9041460f953650863755122bc7dff81831d1fa3bf6d23bb313a955cc5771f07b7955ee9808e896edb30930a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ae6d0745273cc291744e56f2959c5520dd4c3c84435ce9d994306a412452a9d62108970ff62ed9b959077993bb74329ed9cbdbdec027d1f240349511be5414891601131bb73862d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdfdc5e1f80fbbbaa98baaaa4b9edb5da8e13ff00d13d35b44b429c4fe6d98bd17bbb62deeef631652522ea902d9519e29f23ade62246364983ab136eb2d870e81a3497c21eefd3be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcbecd2a0de6aaa250b0a9ecc676a96c3ec7b91fabb27967f38888fd5457a565753e42e9b17112e3a043a0fb17040bdf116ccfa76e403af1e04869fc580484d4bbfa7eac3ff2b7c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc199df24ec2b55629d9d28b023f924b55e665782070ec599e67b5405fda89e45ead1608527d9971e3f002435ca9111dc89dcdca87cc40338fbb85812b8760ab444d8ebce5f9b67e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3a81b5555da4ab51e7b1ef670d443e9e14a2a8aeb1e2e507b05af8ed9b135dad5dd36bd4c1c4b11c53b6b13c196c7e78637c3fc2d4e1555d75ca8ed201cecf28877c10f7681bd87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he774d926eb78204e581f158d4d92f4237e41d0275e8e68f988e767a411567df036153949753eb012e6ba24cd03b8762c456030504c9127ca2cc7ce2aed6a478570475bc90c4a586e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dc965d3d01aa9f4f72796e7d1f4baac4688fd5bbf48e2537b3b7b7e52ebe716dcba036108d21f0ae402dad579200c3dc8abb558cd859db086928b134b7d1a952e85d3a7b1456889;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7629fb0696d0fd32b645cf23ab888cdb536c05f158c268dfe524dbd4ffbd79aa5e49b13f26b935de7e897efe361efe11ac748006d64d5728252993eb023008482f3d41f3c903a87c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f2df413d3d1aa4a83bf6e82fc1f5e0fb5f291c576774bb5e9fcf5585190e82572c9c833c0969250c50c17f293590889766a5647550805f7ca8e5099205c47419d3e9ca8dbef3645;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h374ee9d413d83badd1147cd4c173d8e8282506303295e96e28f4a61a6c948bc6236d16a36cf2a871947f6436270adf617cbe47f8c42163c54eef2ecc1b52e5fd32100aed185b3aa9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a0bc8af7e4d2c9ef3396fa9bb79852dcea19a9cdaea019539a3fcd9b0c0ccdd4c847ccf133b821a2f056a97b30c82aa4206aa69c3af9ea5c293306ea3cad2e8a37b515e1b35c738;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54ab81191728df0805c6027c67ef910d91b76b31e8de30561e8218c481eb70fefbf01e47a7abe67c766bd3434e5e81c6c193250fdab2f7ca267a93ae1858e31ea92e13a7ee923379;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf04f3803ed0ae5aa295f1874f26b4a574a46c05ff1082cc2d83b5f344ccfe42011b62f4f5bb302ead5a36f10517cc4873a2873e3ba3006ef4c4342384f15d34ec09b1bda0e98053c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1265987b7632f22ae1d23cf94d06544698ce6f4bc29c29ffef08123b3a4d70cadb77d28493328107d97b0a65aa93bd535aa4aa8c28e122bb03da114138f290fa9e17c47b1cbc93c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13d62ec04de9e736084d628f1cd4f51798ff31114f544e76619813919e634e3d3df84b68f4dd627ec88a3d2d5525a5fe66dbd55a433b02f2d0f510b6fbfe8b277459f0e4c66d59fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5833a5488c2ae07d3c31755848e069816921296fdffbc3ad50adb9ba85e3ebf499fac659a40285c17a33e6af26c6f6d95c2b29b5efde183ae1b1f01b07b38f4f2afe9f84abcd462;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8d737ba5e85d599d5210354ea158db6477d644f4501bf68447cf229aaf9edd37f1d80ed5c4963344f0fe7d2d0426a1fc4f11ab1c4f3972830d207a50746570f14df043dbce9735;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h343c22630a7032d416868f8ba722b427f07ec33affee4b94cab5f4f5f30d86411172d4dfacbaae9b788e860423c625cc814273c9777a558c384379c258f5e5b98a7bef2fe6091227;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hceeb36b958989a0877354e2da5a3bcd5d8245eed055be77401dc16f99c0caff77df879beebb2bce83d65ae6ecbbbc04d11cc5950edc38a6e313415257594ec47487d25dd876d67b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha93dcd1ea5c3a6e686438d27d960da5c21cff3efe54c2f00fc03cd466fa00fd6776d53ecce2177751406e0ec2f2e9256024076ca5ec6a94075af6dd1d4272e2ec16b240c118a24f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48a5c2a06278b21b92530673ad180786700876e2f807361a06a369306cff908d6f5ca2195d1f0c42cabe8d4dec9c7ea10b6e2f46dfef21de9e6816368ed8eb72f6e53108e7ac9e36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf06fdc591151f98d63539c26167819c57465bb248fe84bf53eeb86ad9e42a3c025725d955f9a5c7b15b1260beab80cb351b355be281d3a293b21849a2561e3db53deb91ef23ddffe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7b2f156da61b69fa379c72b3f8a78d250832aab834ca7d1b30d0350944ccf3647e2eb2579904dadbe0807bb170524289f34b70b8ac0e69566206422c5a39adf0c28dda4e8e1859e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h19d412a0cc8a811d73cd6fcf3a16ed209bdb86dbd869f90a5add40692d414073e5788d602bb2597012cd4e9d51540293afb57ac06a785cabcba08b189fc326e66301135be0d027e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha544139408ac6a441fbd2fd44fbeb9ed507cd53d1d13f7566a0ddc464a648ec7bad1c4a76791d3a385ff6b5be79fa7cb6dff37187375612c1761953cd6cef99d9da762943f8b0ff1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1189e40da2486dca1243ecd68dadd8704f1db63c6609ceb63aa1a04e246e99c03f7831275f7323e607ed284abe2bfd8a9e9cd847b1b12bf951a69d207427bc37db15a442a66c0505;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7201048b8a2270b3d2c911ad153990de46bd1d9124f1828f3410bd13a6a2fc7666cc02e301e6670bb5a23c2af9287f88d6e278180079c4ec13bf519536aea9af32a9882588470599;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56c26704685daa082177793299b77ba4849b6143d73ccde0e6005a938b57ed75328d47fc6242a22e66e0e6edaaa21e965119f296ff4d99851c4e5be4643698a09ac823ae16bf89f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73ce585158e0184791934a2284450558cc5f68175e3ba295135b26a6374649ce00237d4cbfcb900749aafb132e73cd1cf40eec612e89368839d1238f9a933284a06ba09c767796b1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6254054d053acc7dbee61204d9e2b8842bcc2e0095a6a5c6136f769870ac3fab0548412b7ef04744890edb10d10a4cca1bb5b438daf48e9d247f05eef77d23e40f9c44b2a1014ec8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b155b13ebea73ea816e752a57841730c543f49b418ed729313b49c390afc2823a2d949d65f95a9abd743424e7b2b5f3cb545055916d0b48c0c717e936f2a2421187f6e96d6aa9ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f12439ab6f191a6092f1c4ae3f461e0dc82ce63687b8c489a64775abc1696aff18ef8da28fa1d240bc5e5e28874f770bb1138b046efb65f39a517ed21d3c4fcb9d8a4ac03ed69f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a0d1cdc79318767521cc4c70b9c8fb8d10e06e6ad7dd9fadf1deeea5f0c268f844fa2a71593857e983c21d735cae9c7234931581073b84f4baf6afb44ae5f6424d77b5435d8cb68;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21e889026581dc3851839920eb822b57b13ff687c3cd7c7dbb127b750446884518b789c816ef26e77dacfbcdb0f14a95ebd390e5058bb8128b76884f140c084414af18b77645fb29;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf78c201c83dff2cfc400550b3eed172bb65c9d4d19c978784f3f7eae5b85d12acf7eeb216155351b17763211966a275d0e94c55978eaf2473dd3cf65a991a308b54fa6c17ad89fb4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1a1bc4b9ebf4459200b8ed98f675f59ffbe1c56a89579725f9148257e0ed9e3ef0c691d89c0ed2deae4ea7f919e9dc859c42ba9504a4a619fac1177b78b39596763422aee1594ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6de9fb962e7808916f4b01d3c000843b9af8698720340bc44db7e7c21f53716b34750a1c1044c6216d9414bb0a46f1c4f9ae75377cba37157b813e2846a2b0bb249c5c8677d7d31;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heebd5b4c484e1ee720ad5007d5c130b579c347da756cc4723ecb03b2bf877939acb25b4456ddcfd6b4713415b35dde0f8c9f27a8b8210ad1aaac6c1398a77e2072dd397b9b785bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haec510389eccd8638b04ce9184e9315d0ca59841fac06ee58e4caa8b6e0914ccef6b908931a694a2aaf483b499765e9a51445839bb5192156beb89094d7bd5ebb36bce3a51cc0642;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5065fc3637e4adc704066115219e0bc3c63713f3f0422e3a6d512aefb352d9e4725888b21f1247d478ed91aced081c24297708db168a0837defbfdcea17f76b1812be954d700507;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95de887bbdb6cc235b52561f3874b7a93cba955f867edae498feea1589ec755c107e1df5453ee070f7758d72c1a0d24042389f637269940974e19760a6bb9e2c1e7fd44fb8c6341f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d03ee6e985b5ad512c89a2765deda0be5620303864feaf1704a5bed0a7ee11085eb9e6cdff59ec1cc576530fbd7b919b37a6cb31941c83df79908007809a38b47aa938eae0a939;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6bb9d9deac8d02932502a80f0a00be220c16f367f9e24411c93af424893a5563881e1affac3fca6cd88fba48b23e27a76aec8471bb0b0e4baae06f1b6aae5a6ad99fcd4bcd96b643;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb178c2d389b63ec634712224d2faf58b3123e4ccbac4f373f3d6f474db6d948deeffa6d1c0140fddabfae80c25e24865914a9518487d31e35cb0436d324a4535875bebc876e763a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fdefa905fcb7979d12d24c1b336c9979ceb0034c14baa08b70082ffc497420b16be4545f83958c863d75d560c976102847cd92f667f7f4d026d7a9fea4b9edd08f0e861b07f6e19;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d29f5c1a0c780a9f44c256eb8fafb0127fed5cf8e3431fb6014cb649c52521f512fd920e723cae0a05a47dad79f1ff723794ba4333ade1babd86b39d0307313c90a1ec8f02996be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b67f9dfc508ebe43ab0739129da857da0a906ebfb299c20a0e1129fbe4e223764aa6015977ebf919602f48fa2c6a4a0480d6c9c99ca19e0fc21fac6e618bae50c5741a84cfb3861;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha891da6ac19457f1c268ecac6eb284cd05ed6cb2587586f7d0d918a779dccd3568d40a7496212e5557131721d848416d17d0131ee0397e3660389c32dfc6119dd2246508d7e0e8d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdb5fd0e269b665b2cb8a44304612ccf28622c88e0f7fe3443cd57d0c321452d99590a9373148c28357a98a344b9609e1557aa4d6d6e8a8c206411ff1a8c7b0e9fd89d4d5a100c19;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h628d8ffa11c5fe3207ef669b926873e53cfa8bc2c401b25b7175fe275fb18bbcb3b94fd225866cd0a094cb35285006112925c4b449592eeb68cade457c8acf75ed02b603eba8ef17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6048c4a6c2d5d91c140c10b30ae1bd444976b4a2424ed4fefc2fd7f4ec669031fa3847bca104b882c8fe09b9080f69e6d1d508e9d13f318b6147714f3b3cbfd5f1bf3e5c435d705;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9859f4c518b87d06e3b7be80a95e495a9bfeae182fc7461fd6b340aa9863ee1aae3f89b5b49ae9539fac42a330ac4c9dc112e607f33dea332d5549b35bd8ebdef846d3822e5e9a9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda4216046d29b806784291a18143305c65781c171416a5d72050b43dbf5444612b3d8048a66f82008c51143d0ef2dac6b3fd74de5a68e513d7defffc8bc24a7ab49f26af4318063;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he099d9177746cc916e967e22163f7326712964151fbaa3b89cffaae636a5765e0c180ccd787ef4cb8dd9b0ea6676f446239872269c84209b2fe57c008ad28dbbe9e3f364e5f6d501;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdaecdcee1cc6a305c972bed3471d0176429cb43ac87f17d1984c965509998cfb883592d7b54cbb3523efc394fe05461e80ec349cb0b5ab66af862b2c2301347dd8d9bf44a795008c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1a747dce302bc6db191324b8438e5c229bd5032489bfecf0f2358046cc679cf0179580dbd8a5e90cb06a8c28610f0516c65f5f00684193edb5bf2c83c64dc32b245e7a90130dd45;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e28d37927ce57470084c4621e7ecd9bedd602c8119bce4b9c742303fd69a56920f0d453cf67cbcaa94106bd6b34f3156cce7fb4781c06ceaed423d291db9174af71603341d0bf37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc26706158f02cee707f1f133b943d66d14282bd90513378df97a8bc9ab2776c868a7335a5a2cf17faa1f773a2bfa21dc8f8370f463b7ef674f167a9be51b3abe35095c3f560e7e28;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h522f04e57c040444504513ee4d16637ff74e87b468e7988eedc32b18b3909cbad93d2c4c594f45fdb7752f646d0477664539e38c307d1aeebca60580341ecf4b350850ff5d3e6368;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd16adbbda693b041ba3d5e81fa66b97d4515bf603e6466710de5c622160d5d213d145f9ab216c540ca4a1c623046c37f0078582df4039e32e99372c0b3925ec87a5fcd7999847abe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae2862aaa22ecc9dbbbbad9cd82f52889550452a2ae935d8e9b60a0f3dd45c5ed348fb9e50746f8a476deff1813eb510cd8cbe6905f88097cfb9da4ace483cee15d888465a957cdf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h308b97d0a1ad7335eee784ab7e08f02b5b0ad8e47440bd2d0e6f053ce242977ca9da0acfdfdc3b8170546fc51a6bdb8d4663382df8d0b29f7174f1362e19ecb3de4cf2fb03d62f65;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1615b3bbd2d43ffd2c2766f90e2a9f8e39064c8bc6544d8e42fa3a140d1309ae73880192201cd38e9078b8b6fdce8c7385ddac72f02d8398445272a61b43883495132f9f5b4b2f2e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde5fb1b808455c1d04c9cb83f3394de45b1f2bec9bd756378e5e43b55cceb1fa27b41fef2136c68f65145278aa383a484dc43087eb4865cbefd076ec4663559dd2fa4c2572cdd00c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5c2c7386bad9d91c128512835c9d0013215a6685924a9d3d97729eddb1cb3b529ff2ac9975f66ba9b3054bc18311ffc6eb429b68133a74ee8002ad259b880532588e5eb26c38be4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca4cc6c2096582f098278860920c34c9de8b942bc1c09d88d6b5b251ec7b81104d01c022585e408abc76a2105980f73d37dbb15c22352e9d6614b83d286fe83aee4ba3b0cc47164d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2dd906db9caa930c915da796210711b9cf79215cfd8871ab229921fedc6913e96d88edb13db287cd3953e363c3927c57acc9b3c215f3bff2f2ca2dedeb91517e7b378b2756a9c796;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95178131a5c297435573a5291f41bdf2325de483d746d61e7ffd142af3be8e60e314d737a704423f03523d101597737499f5555a71d0e096570a4a9eee6badd6a0fb3ef12dfb9161;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48afef09a2c05ac19b754d53ad256ea0f351883f67cce5e24ba96bfffe6aedb071d26c1035be423a85cda6ab8e13e5fc4b13b58c16bcb8f1d5b7b7c9000468df74f3d65fa5b7b252;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4d3f58ed983e9f590d6a029147eaa30cf990b9cf790bef30b169f0b7588938a6f0d85a9e4fb7421f4c2a137e3be5ffdcdf243655bbbe09d4d1f9e606cfcb8feca83e65e8e195c37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdf07514a78f218566606b195cf12d4c3af73b24bc83c7bf99532d7b213f099c23a22a889749cdcdf56cb7209af0a74ea8e586c4776d304105444a804d098f508d4f2e4642f9545a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha64c55e61625245ec41a121baf23f5f5699fbfa5a7d89460a49cd6edb4f44a3ba8befb6740229ff866abddbee0bddd03f65c256717b2dcb4e6ead7cc00506df1d0bcc84bb76973b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9efb48335d971e3ce49e0d6de6f46f26e9f3285200183a49cdb857d620ce5a63918b7b16af8b6c79a59214fc92395d485d73d516efbd0688db21188f730ad6ba1a9bd8bbf8773ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h361e925f326e167737d77034e88e6bf6ee15d1752ec5337bb8bc6aa72ba3bd7cc7645b2ee66a1bfb4ac0d1717bffbfba2dc6ca0c0aecc27575a7e4e35c5b675cb88f69f0fb1afc30;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6e00154941b2233de21ff5a1a2a534eb86119d39b2c74b2bcc7d87f303b1fa4b0d8f6973b0761af952c3b87f03f55e911657545abce42e809ff46c041123f2c107cba15e9d23287;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d4e22bde49a9f8dc53b16afa2b80ef60411554346fd4eb97f8594e786575e2729e8ac3ec3be53a2c7689bac1807400dda7fbd8a77990d4b206a6ca2340f5a747daa6e3e74039ce1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64df55c0baaf40db46a94e562d298755fd66693c302d4363acb9cc77149bcce9d310511987db9e1a1abf42f3ded1d5c8a07d0b1d58d1ef85756e52492dce794637a5e5da539f0d5f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefc53abe97003b4cd40a09d3a66977bbcb7399eb62799eb05f5c9a377a8bc7b54fda23b925fc9cb5bf2f746d55d687e961c7e8c038dd843d48f32d15f78e1176556775f435f4f675;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40a5d1d195cf618bbc1ce54f575fa1ae6e4c1331f9f7ce1bd565423718b563ac9e00842a784500dd933243a0fad847574ae8706779d7fe48630372859f320573ca122deae87b883a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h837644848f45f6d3b007c524e95c6fa383f1cf8137f7965718e837d7455eefc386129022364273547bde7e2abc4fcce46c37037ef9c019d392130e7e0182f8202a2160de6dc67a2b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf03b6ff86380dc43a384e013ea42002d3cce819bba73cb484d40e289ca7423c6680bbbe08ebcffaaf293a94b226eadc7d065847877281c5c292b9d86379a5c2adfcebcb7a45ffb6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57e5d604e64eebd22a087ca86bed000882cf49b0190c8794b6bf11bd6a349169e6ff2e906ae40051f552ed9b7c7bc87d32bcf04560379495175b83b6f63511eec317acac105aaddc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h526760ae5d904e94c64c1338c9040ed2487ecf8b75923e1932e4c016ca1b877d6b06b0087b330b725a4a6f85cdbaf955e0704bd63a3947f2b903693f17b4f120e2eba3bdda7f2ecb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40abb538c654251de8a8e2c69e7f97dc9a770806c325499d602c7470a2b63919bc9f4e69ddc915f26fdad560c75335a0a689ae07629ee4da169ad20a178760c234458a9f0eb5309f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2190581b29a47271b52b5b1bcdd02d468bf4a8c460ece73a2bb1e64ef0ae91d281efd239fae33c9c22b1e9009960f5842e9182fd30c506b6792cfbee11d71b35d0941e6662b5af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cfc1b891559a958da9447b3b19c9bea441367cacc9e5871d1d170ffb258e0f6f9f5d29572e7c2c1a8ccc347df6b595f6be4f244058cf5004498186326d75b2b5eb929f61bb8cbc9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a3d995a05ac3087b30c116c61094e04a3d6502099d442f68e9c6c73015cdb95eacc1ebb0a8a318534aed8946f2c79e5da7e9ca23a176e89901dca0f95f41d45393469917651c772;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3b9aaac90b0838812f136e501c9793d3a45dd8a491339a709637a02d88ea0ec60c11e783bc0e0bfc312cb8ee988402801bcf06004d1d47b886c698acc271b9997aec36c66eb4052;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1bce20698ae0674c0d44a38080c0c4b428742aa07ad167d26ff6b9a87620e84a196813213125fd677b30ce2594b3313c68ba49ad885785e5b563e7c9be64c37e6ae7d8844f77937;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h843986828ecbd0bba16acff1516165d8c86da8263489c420b16b69f6eea8e48635e150cad1e56b9f6bf9728a6be1c575bb12c13feb305039e3b597a2ad6f9b0ffc9b06af15447c2f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25a2e7f974b169f5158cbb19c6b9d38da715f66cd949294e31354c371ed4d93b21af3fbc99fa507ce7e1f3a28ed5506266757a498109124085ebd5baae58e7b928bd94f06d91943;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f520fd54bc7433d1d800c8d15a46899db2e506afa54eed3e31e0c6a823d3d51628d7d7a4520210bf0caeb0f7ca44de9ad140def3bc5cd8eb4b72d7c0056cb2d96b7641cd2c8410;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc281f8713a2036beb80f0cf152482ffb8b571fe4cc531054cbe99dc99ecc6f4be38aad8a2de9c171abbc488273f4cf52d766c09cb3b7137f0ecc2b0408874e2ff6eb700115d9e3bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd20a2ef1720927b0611ac4953ea9cb361ee17b5938bd2cbcaf3a791806fbcb736796ca1f0fb0476553778972c35d20e5d96abe676261d32d954fbf32c83926a77050dda1482aa83a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31e8a7844f2a6533b23b950c0e9a735df8db0ff834190088be7525fa807ad61a3f3674634bb192420231b5a9f8ef0b81ecd4a8b1e653267ceb069c4b32f1e51687da590d80b15978;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h961750ed3fb63b6e1ee2091a774375a56c9f6a5b9aac8810e601e4146b7a5bd3a10948117e795045d965b488dd0803f3d702bfd30316a530fd40ce3089fffec4679275c2193d0254;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc3c731d94bdd66028253819d345dff081f72b001bd470cd07fe1c84941d4c175261d19a6c520e9fe74fe9538560a45bb0ca6c13938d17a8023bf341ac775eb92f3fc39f1612d925;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h768c369161f4f52bf44c1c4cea00534072a522adc68ca76d5f80d5fa1faf63437892325e972bc71ad37a0fdc0ee7590ce79d55313b779dd753e9ada3972d71fd15f8c271e0b6b930;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1abac07613fa3ec19961ec1bb6a131cabf5c4b5a6012a369ea3ca042c39b5dd19e7b67bbc5441ce25531aa68aaa014423dce691e98a84d41567ef73babf99d5209c06168c478c35;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e1f1159975fb25d6a9307ecdf8c2328093c949d235d1778189e2a8569f1b060b1cec5eed70c0f9e31f301b4d49096285cb1b7cb3991e933b11f7ccf9c27742e45eff7d7ec01a7dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfedf7a7498fddc0b88559fd64cb9656f6744e8a2edcd8ea1190b50da61ecd5d4e742afddbc11b93f8fb5ccfd0330511a09e3636be45c721286d48a32224e779826feeff39eb56eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5173152b4954c78abe7b0e8de59b32dc720d33c900da88c57f763493e32d75eb5c66c84d96764b45d6f92a807a307f12a57b587d45c9368e153407163db1d4016730a88e510083e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h172e27a183cd15fa94b77b866a812ac3d39e4d7b93197c61ac620daf7eae50bfd258d32117ad53e5df7cbe785d1a53dade3647e42ea48f3d7efeec36eb80678be22f1d274210f84c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9388f9ce719aea00ce0968578bf752b41ef487ba8c2bcbabb67a0b7fe5cad1e3b2f5a4fbb7d77161d7a67e3d11a79105ca7ff3cc6abea1cef012860971673c2e0c7f39152edf2e87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6710d18d1a8c6f84634746adc8515a23d78a1472830d44967f408969f9258d4aa002f084fa2d2e6a2bfafa2db056c13a820d0a5ac85ae7a579a4f1661593e36adb8ad9435d159508;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4c3c577f57566c1e90deb52df67a0e507ab122911350f0024cc4c714bca3aae99b8ac88070a73ea79555846f38447bfb0825badfc4834b757e13abeb108231b08d88cce4e495ed4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89b4d8f66c4f43dc1f4da4dccf8cfe716787dd57dea64b223d9b89cb219ddef1dc46cfc0357111528f61f8361384054a3ffe781dce80ed6b4a84e3c5ceb97aff3483ea881dfb36d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde89bef57267178a3aa2f81d57be258490610883ec3b7a3e75f0287375564e7fab42e1bc0bcf5acdf28e450c7177222ee91c5768dc23157828945c2b29a818ef0045d9d9ad6bf9fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf85f3dbcb04fcffbf382662d6a99933df4be1612d37002bac2797c402e2cd0befe8edbd71e756c9cdb96f6379a70ae0160a528e918bcd17c05033b76202a3dc2714f1929fcb7b114;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bacb452ea4a10a43cc4e6af259430486aeddabbf8ff231e4cf5d59c462bf59499bd779bd94964471d3f33691deda30e7c3a5fd37c731e721d3e3c339e19945b6914e58285108b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf42de73932d79777aa7e3d494098e905bde9d787914145783fa9a42862882af19f3c39ae20875cfb52de8651bb953e966010d67213824ecbfc8969f6abd751dc9f860dff25b2012;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21a3fc71be578932fdb8f0431cb7308383e5ad5730b0333d0911301f68b5db495b90afd95c9a5182bb0a1fa4e2f9fc99c96e78908ee9bcd1853969c5ff76603b02ae282ee8bf7125;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c76c731e0b30b3e83e0f8c61a50d61cb9a4766ccb7c6a4e9bae51077b5c2ea74e38c1c5c3e6ccb262227705dbf205cff01238be1ddada624db5b672164c7c285c07ffb947bd786;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1aaeb1fc5618322fbd1b0f1870813eab40c3e9c4a51e6f031acec8a07a889ac34e158dd1ffa2f2e586ee5199fe0549a6ef94bf0720bd9110c838132bf5abad323634369dd10c0c15;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50cca54fecaf2bb0c75c21ca7d11a8a3381d24d731582ce0ade33658c334aa4072278aa968222d4a052a3ac0edec81aecb48fbd9b7e2d86bed093b4114d4a25aa00f09200ce5737d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e57d1cde1692f654998b2e6e43298d86c9c8ab516a6bed9c84c8db90fe99fdf6f839889cb74bc03b1082f9926ca47e65af471c418b4038d530485c05bfe6991bbb1fcaa5bfc242;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he34e8ecec935cf4171df93616efaa76aac25f9d61452330e9a2f9d233141656c338cba7703c5454999c8f58624b23145cb205d1bae56b597450233519a3c669945d76239304bda60;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cb5f644743c67e04c33f6783c46de8728113a607501b7c884276a7411f97837c4d82b93db7503ff36b7f291ad882de93119da03a4bde0c37b2bba58404f5120507afdcc576319f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc2dff24fefcc77da321c62d4ab3bbeaa4d14f36c1909d93a4091aaacbcfce1b9ed654651083d275775de903d94fe22a769e8e3d5767292b2fe40151b6a2524687be2b00664efe73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5c881bb3623bac1329087b847a25fa76a60d2f68745f1516daeb972300e76c1eb4ed600a6f172d41c24e69973850846152eb6242638dc09ecce6c1837f9673463934f5215a711c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb56cbb19ccf6af32ee90829fcbac37081f16a91e5246ce4e6b6d39f0cee4b94a3746c2fb0f9d321d071ea947fb0601fe7815b7d65e12834730cac80c19fc8740060a1231a7f84ea2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa05c62999c169ef9487c24e58158c784765a70c3bf6ea08fdbde2424108f022ef7d620a12d45d5cf0a1e7617eea3193a1b1eea04b7b3af9b5d89472e53483c7fcc983b338d15f0b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h695f9f58bc64a38e6d92c94c8377ff5143a8963406087e0388acb27606ba43b9614627f2e143c95b385a154c559bd5cdb51cd11ba031547a5e72943ebbc9f4b58668ffba922dd261;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4bc186d745b6f16dfbc46032f4f4de54a119d564d5dc0e26ffa42020f3f943c4222955e3b0ca0dc1d6b071ac9a28be56cec5aa8a94a82680ead9bfa426b3c91a9c150c8e2dd8f2c9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf701832852d33b7fa547eff53ec37d1a3c62ff8d1443a7e21f31d05cb89d5bd4fe51878a033a8e60aa4de3b448c758109e21b9d58b819810371341b39329bc5253e07916744c4b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd3c0fa06ad1b75f0806ae4516ae4b681cd6ece760ba01dc22d0bce74e1a35c79862c483de87b088d5bea215167047f223a09f8ff58f44fbf351076c8f8e234e1d9b267dc2f6a5a6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29375e5cf4b1d82f212a2b92147a41bfeb3a2594ab236b0ab436766d1063f3b990ee2616c2b96c2a4092c8ec95253eb83e9edb6efe9a515e6f816b528080440a28b2e07d671db956;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc860f2b7e71d3d624b58f4c8599832c4d4b88e45218fb510e3b836a44e125b9183db4fd126defb915f6de3d58c64483bb5afbce3312c5e3a338dd58307d40d00e489f6a9011bea34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58b87bcb8f24556d22f1a51c9db7000e34e627a5d964e1a05f18d3b08c02dc4ad39e703c62df46f8cbfb2025305d4b55c01f4926901516c751d229851e5508b9d5d1764406d2f786;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habb9e2af4642097651e828981cba16f9ff96950aceab270c7cecda1821a6f1313875d74525eba37b06ddb776bd5e2c1c0f20a09491f4e230221dfd5cde3455ec03ebae084e001061;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e37bec4c709efef8667e3f904e3768648386ec169dd6bd73e133de067ca5ef7ad93ee1d10fd50528b08d6c1d3ec9a1f9fbf821c68d8a76ae6931d6381e913dcc5bbeabbc4088bf2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22815693d7d25c0a1ef7c04e77c55846c7bbd27d9f5ac3bcbfda74795a8af18c05beb34b05a4715f69b54d9496a00648c68bf08109e9accc67251c6fd129c8832e90fd75d7ab6316;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h667f6cf8bf3ca921c50cb8010c1872e97115e540bb186f1f7e171f5be647155df06ae8242a2cb2a21d7907c7e3c2e3c0a809ee14b436f14ed16047f1f19b906bd95b4f822d30a110;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7da5347be6f5f517cb3895e00f93026efa14aa062672c4a5f963b168a2c3367b87df38529ec7072bfb32fbead593926d8ee45aa135c1f9a9adf2ea14b516513a1bc1b13836394cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6796e45bc71097b04bc6cc47b4744b96351719336d059851c9c05192002da91f741bf2d433c9c54262bf7c0171e1afdd52410a23b7d824a0f94f0a6b979903c88a4d83b269c6194;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3890f09fb2bb09f23834f1381ef22a74932d7ffb4fec996b131367adbcb28abe82e95e4b301bdad9a9dca42d37260cda6e1a3be9ba9a8fe2055c3cba648dea32e41bb779aa11c86c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7be4fea2ced0086ba883061e7826865885d29cc30ccf09dbb26105b1fb1e32f87f3f4349339c534c44a0bfad7da13cd70e9e1fe4106485f754cfb4da8cec016cc69b42353e1f4832;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7b80015e1853b5487e9df54ddb483ea3ac82e075472c531c5d921724e608c613625e3fea12b238eb2f96a80bd1fc5537cf88c5adfe84eb5d72383d669295460f8a6958a410b70bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6b6c6556fa070413b4424de6e528f6e86ff464f656bd9d7d03624290fb94b4cf12bef2dbfb3d3a7ffbea60b74a385c6be0a2d75ed5d6ca53da897113558de310ef6437d0cb6d6af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd433a111c89ac1566deac664235437a9e9f9b403dd9e5fa44c848140008106305e500d2b5217ac1a797689ceb969c374e66949cd0566f8077d40316f516a08d7a457eeee2fed1b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h796ca1b82cb2437265b65e94aec28eb4f560ee9310ca057a41ff1b0d07cc24f4db4d44671e1a66bdd783c504ae19d8c9c647f515dcf8dddf2c1c324a8ddc520f65d21ba7600f9763;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4bf75618eb61e16e0a4b94c003e59b196a6036d2ec1b296c31b00a5408026fca1393b60f904be05327468c59bdfa500116012d07d580b282499d58f2b7f4b0dca6ab9854bf9adcb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h554a4ea5de4210336cf45f1f8605c3b317ae900bff3665e8a0547c6134465b6e2b11210af23f8cfec8581a3574a26b80885724af4ae455dacc0b8c4cc7cc19a642ed401d9c70eb49;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf79f0bfa76ddd29e58aadf53b1296342b39cfdf1b54d8c590c15f326b713676fbdb298fae5c95498db41de91223d984223a1fefbfb6b3f8a0a8e71fe4eae28ac450a5392676eb2ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd513767055d029823c6dcbe187358f92e0f07c884a0139b81098c49fe230ec77c1d293364a8937872d0ca5c68d166f29921de3991c9230aa53ba3bc5a93ed98f6a5dc25e006184f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a7135f281f71b8c81a1d2ef7a3dd96240216311a8e85aa84219e75f17504c5a08a4085390d493305f6eb292b11a54137bea6e2ea142d14fc3305d271e95b78ac0432ea9c45ff1fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd896195b06650f22c6ac3b3ce577ce5364346869e12d0b3a45dbe386314f5a0a5553a9ad547e1131850c4a29cc713e1ddf1d7c24f19fd8ea6009ec8acc6b7b32ad695e8c210158f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he84bfc0e84c423bb2974f32e812030d659e1325d03236a07ff6b04b1a5fdaf789067467f2b37909681337cefa7a5acf03c7c8285d85538bec1a8ab887ea1fda82e978797d239f88f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44d8dd33f01a559ea8ad866066dd4e2b35ee0e815485503f65ddd64c0e3dae98c6a50aef8a7e01f48c392ec34b9f07481fad3b13928c31c24bece8300b7427795bfacbc717d11f47;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4106f50797980bf06ec90180ce5d23614db17de0ad3fde26037b5ed6aee1b09636575726de59af2fe6ee0c642d7bccf886d37af1166b21c8cba93b5db7f93e3059196cda99e736f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9e0354f014c2fcbbdad1cb6234301c2d6fb14ff6af620e34d4d881e4121250bf2eff706dba1698aed5eeb80005f5a1b33fdc881127b7670fbeb28dc9e54b94387b5ee33061c0fc0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd03d474b92fa116369c80ffbe28e49c4f3565610de81979a123eb493597ff7c825558f4f49261b096b377d16632ae44d28c028ac5c551f087a1f533bb5ccbd028d33d1655f493760;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hacd6a30315249f94fbdde90786e94bb0fb7240ccbc4376e385f057cfe9f2831a77d3bffbb3fac088a07b9a041ef14b4233d2c33dc0ca0e2cae76be64fab90d8267f28a3a8f28c8b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h456f7cf8b1b43d4d70b606de48e6b28c182ca29d923e4747480514b0df2dff3bc45968cc3e76358cd601a15a63df5d94b23f10bf3c537ac1ccb71ece8162d0f88825a753b2e741b8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65348e1982a7eb07a0397f47d2ef47d0c3816c666c9ff68584b48ba24b7049a967779535b0a98bd1bea479728f93e59bec4d2eb720b9f511c1e24b3b069b7b68488ea88404cd067a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3a248131fddf2d10c94f23ba87ec75fd170b9de26f15ea3ce17c57276e81831473742b019cf1d96962be178afd80d95e60e34deedf594da36d55231730e30378d3bf57bac39c9bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3321bb3c8c0468521a2317060b3798dc5c0bcca5f58eb4ffd098eff6f1b8d1deb5f2d7c72954f5a7f23362fc2fe057feb8bc3119fece3528d73f72d39961c5891fb4858008771aba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22ab93e3a190cb38000d7ed44fea6bb2e7a7c43bbd51a213a95edc4e0d4e2e25882b7c3f3bc38768ea60b23ec5e01f7442941b1d4d05f41a2bbf052189c6a9ed6a9456b011c82ef2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heed4c7d3466d22a211890fb53d4dcf7f53d0482c5da4de560f465300e3b744fe2db9472cd1f068952eb8f65b4da5302b09146c224ef192d615ae040b9a547108245a24fde4b5647a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd843c511c02441012e9d1aef3886c8f3e0162d66280e71a39b1faa75be1244d7ead902ab6c1aa1949a7d5760642cda491e36edddc28403094abe9006f4c091b63dab00b81fb3ce0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b322435931c9c1d6c0203347f5200681824f701f52fdd74e2d721e7cb6a3df03eba15a38451634453e6a5b7ec31d41410599a4e793a1d7b13d5708361dba4a09bb58cb3b62e60bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda9a1c2b027a54bc37254b8f3bbe91de6699a5d941f22c1637d878327c5953b9eecd1e40823b627279d338406b3402657263fe6075cf2c09d00af1bd64b51f8922968e53ac4dab00;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h484b3dd481d2361cf7b45f8e71664b73242fffb15ca786fd1e728762034a05ad15ef3165244293d260865572f3714fbf8d0608c557982d4b105def39ed755509fa387718f1281ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f03984e1616ea153dffe4af6bf7b10a7a2178f25b533fc1a4951aa3d8f575fefd03599e11a3281b1ecfd7d23a43e9068e2a04b8b8a8e43c441e8090dba10196170017f9d81228b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88b8f77b4cac0463706aef1140048f45c83000d37576fd5e5d4c613f19ad7fc105d4a4cdaa7a3b2c090cbbcf11d9fd75b04cf4dfb0990875dc05738dbccea62951477ad2e808c6f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5348e7d17fbce23de7617f9c3ad3c6b2064a03a88d00287807f9aa3ae59715ad93b896da24c6534e8e24aa1737867c56a8323f6c9f203b4c1093225a2bced5bb81aac8552b4b06e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18d1b0e8ecf5cc62a811c5106b379a230c3e76fedf8470fbc3a39ccae530f7170aece3e3ad43e370db05e4b89bbdd37f7c7eb9a2971d6e3f5e331b6815b75527f5bb64890e8d7e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa0ec26512088ce75d93b6cf2e3de0940d91ff622b250555874a6c570294ea300298a910e612824283674724f33a114317c8aef4dfff8c41ce0184f424225d812d58fb6c7ebaf320;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36488a91e01ffe41ee6324407b482b1e0da140ed604cae7d3abb21812f2936dcec6a4e0daccf3095154a878bcac0452e1af7b9a450bb6a6c344db1f8f949274a5d516beb57009685;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cedfe14314e0ee78ea425bf91412419a0c0e16a6ec3bf3b2cab220462fdc3c2b9b70a4813f680167d463d1d43a11c277c288873ff784524259d869f0a86575b73d9e5d2cb83ca90;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cb8f7b5008bb0030a1b7ae72af17d153bae462cce08a107ff1022b94be39c7bdb543bbe5d01f087919a0bdb2b869e6ca10cf9b9e454b74ad395a9bd824068300d4f79c2b0088416;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55911ab35c7f6ab02faf6ff82ddd2b8d77bb7c44452b4980ac1341272de92e6108ec39c05bc92370e27ddaa23fbf8867461f2e0601242445c140363cb0e9b02675666215696a7f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b04ae44b5fa9dceaddcb6eb637cfb136790098badd93c6989ac970daef1e66c81ead02db0dc7d0dec1188dabc6817aa49b20f52969dbf4b279e128f953ad5dbd7eba742a726dd69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81232b42186fd220e2457b625ba4db3b8f8486c2566fc52da08ffbf411090607fcf4ea686980a49d78f2a3e0adf543befe56c015425974a08b9d2a8307fc576feb8e0d9a34da9fc2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75e9452a5873f8189743c650f11e7289adf205f9c0c5a1a8b1753677d5669f72c4d895ae47c1b0a226a3a0ed13ede0f295a7eefae65a235b6d4a2ad8840d7dbe50b7e69758bb19a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf82b73faaec68263214eaf8f87858bfb81b2bdd57539bf102bbbc4668b9264fa9db77b92ee7f1a48a8ab18a2bfac0649f771b82a10be232b68a5c5a149fdd5cbc3ba4b82ae57683;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc1e055d4b05da845b32aa10474ccd8f2788bf0446dcaea848c3321642712e39bcd04248ef673007f6c49194fbc5bedbc113bfb9d123ac85baa7eba5333db5c3aefdae637df37499;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48e437ff0be6487264758f878058dcd0df4230a105dafff1c7b2f81f10311c30a07426f70baf877fbba0676a5f467e58070b57ddcf9fa83effc46601148c444f784ec0ac89016699;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce945de111e64d27806117b4b4a79bfd3e5ad0e0a3c6215e6915f9e0aaea5418b8b970c786ff156418c7cebdcdfc9884e3229a9f068a32ee4c569c75c8d5a8b81fffb3816481e60f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cada0c27e2be6c769893c0e171f9dcd437d420144e00824db7f80f51db05541185ec87f56962d323eb1bc84b7815662d89d99aacc98c675972526919a564abf59b5059fb724f47c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b3e1b7c4a4fb78eeb58071a15577fa4f1f7094cdbec6ddcf976375bd5f5987913d6466c1628e0a581725238d44edd0af251aa9f9a5e06153cc996b96a17130f14bb6221460e4d8c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hced8cb10c72bff11702b159b3fc87f0eaf481bdeb9366a49dfef7a47f7896ed7558ec063a81d9e2847fe662c1804e0ad658d3f3a0fe4f487dac2c5d8801813f619e8f53bb4d907c3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb91d608f06edcc960fc4b792e2810c745e17d3cc6d770ea2802efc0180cee5279e4ca366c31ba5fe2f4b25cb9f4cdfbc977d8be839b07a4189f770f18d0aa4e44eef087022aaa319;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h151b6596f72df350b8b1280617941db6623549179e59f0cfe76bc43bb49d2ac6fb92cde9bdc82b3b811155cdcb0ee0c4adb29d81bcdef53a1107c7d8f61970a04b24ea8396926bc6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he680255b7132f5afe02a41d1f6ac572ca7715567a39fbbcc9ac1a458107e053d022a9638322bed64ff50036cf5f38be1ab6b97f96dd880a867cacd6cf6fec850d689dddc5567faf5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haec427c678935894c8faef1ac99bc78b3b659e158dfc0cbd53e3ed5181c00f4065fb234f1a56afc89addca7d146c21e95866698b24ee0c05e8b07c37d91f6ccc79964c6734f9c48a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50ed3026ba9654ee0805e2c2166a9ca4e90ce5c430b4f9ff24cad9105b2fb4def6d0c50a78ac873f3e21744bf9ec79bb83be162dc9085547f229273623c90f4d5ede385ebf5e8b80;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h133881a17629d5f102e099ff73606d36d735578bde27c2386e1771c461c1fb004b401881343addd244a81366511d97c5317182456630da6d35f3fbf727e8f579a211f3163788e327;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69777f001e7201e7f2c3f08c28b130e2d2854556bb4e4899ef7531f019f06222da8236e60d3eda018ba8619af2adf7ad39f1667b3afc4976d571eba528f713c3ddf0224a1e8de99c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72cc9c494201eb16fe6b962ccfa9d7ae4197b4fa8876920ce619d2fe8791fd0804c82098bbf54447e4acaf20bda246d0d95c83d351d80b15447a1c15246abe87f58b2c925ebaf813;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd33cb7d028f65641aa3faa18beb67a78330ad2f6d3b279debb0359560fc63fb581b73538e2a34fc04e6670b4303d45760114f4d39fce1113e788f98854808d7bc749b3475dde158;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1e8a96426c1e25eaa1404c34d6c440d0282c96676bf89ebed0e5f329d7b5bf8fa9bcbd4f5b16ef879c24b394b7eb80ffe65ca575a62c9e190d24237322528463572859f199fc1d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b2e053a74fffa92f8472866c9e9e58e491399fd8023c71152363f4908fb1446f5b9bcad165d1f876b0708875e86502ad99867473c31b12b94c73311a94fa26134b534320291c5ca;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb514810640bb92cba41d98f13ed75922909e0127f160b5022220c57a081fea110b7d067ab500aad7aad67793fec59f03328a595ca4c45826f64a9f5c2fbbf64e602ed12522e264f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf76b1d4f42c8aeb2e668c1827ed31ee11b3afd7fa1db6cc801ba1ec07d7111df984d5d7cb98f9c9c80e95de91e49cb1efbf0fd4927aa185a20b89aa1cb1f0f881ee7e4ed7ac00d74;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2928da1c1faac5bd3ec1083e238f7534399b1c6124fb71c14cccf3dbbe7df858d2fe4c58f7c6e29dcd9f210addcf59adc383bac99539056108b5b8b30e3dc98d3e6ed84a4592761b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3190b77780ae0b4944d64e52277c13cce5fddc556925d2ec16611db60c5d0adbe29a1bab50a3fd91591465e9eef3c659706a289d13746e332b7627a62872f4055ae784668290bb77;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6eaf6e2b67914f48c3255da45b833b0233bae6737bddbb45b29839c42d2f78b3783e57b6ee3b633ce73221613b530eae9060e81e647795f876f0325abc46d8bad64ad46b82d68037;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h257ea7b501b3cab8e0fb13c3e1f121ab4b5145ba58cfbb6eb707df191cf72987fcc9e5053cbbadeff09a38a1de59344301f96d753d7878e156ad11ec2c53922be502c3572badc082;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9570b6db34c711526d6feec41689a26e4e6d43efdb65fbac3ac3c19bc22616ce12981321f84dda9039a81a252787af8262b619ae3a0cff528c1ac8322a4905974c476c68ffbc45b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h631264e9a83b432934253216a50db96a52fc1b69a9b6708d0a9ea9633a2a4b09fed2054ecea8aea10fcf32ae01c9434055f792b6c688909124a2eb168d32e82d4a28b2395f47707;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf42221439eafb67e85f644e9d9eb5f4c2607f626d68d1d97daed47b30278cf8e040a930d03a394b04f305e5b7c68e1804cbf775be0a9745dba0ab325c42d95b81682f11829ef6437;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h515019e18a90cac2f5115b8cbdcd76b675bef7d97c36dd127ea2fd2802a0cc6d60008381a2b4fdc4386e5e1385be99d0a0a6e45a847a67b44ba38baff3899b5e418aa8e8943c4a47;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3075ba1921704684549c1a4c0ae392c8b016dc960d50f8407158f74ddedd2db51175f7d37acf0f74105a51d276d0fef880208286c365631492eac2893a36013da5f634b0b543e1f7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffe19c4f3651e3c7ded050ea0a63d8a35f96f7af57b0c61a38ec88d89b9f91a3b28a14bcff3132ccd0beed84b27b664448676226dae7596f995c53c61a4baabed24007e261714a36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91b3c0fd3f3b3f150797322b4c4ef60bb9a9098979133b755450b93ec817ee4635bf5318b8da245c5a743dd722e4084a504c5ce65e39cc966cd4ffcd4ce36fc1dd42c9cdad3df651;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7397332c5990993fbee60aba208c67f99c8e9a18877b84cd03fe79c321654110ebefd98d6f2affe99b415aa3e2960a5f64dd321397b0df4d8b107e4daa22efff895506bac5120be9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h762a99fce9138e2d8b4af1c99d57a18014a1bee804b85786657bb12b169ec4a5a334044adb1ac2663a98fe79c2870bf0452c65e387f5ac4736bcf1534e6fbca87673853e5c60eb61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed4f8c7cc4235116485306729513766780cba1b1ae02980857e0040d89de6b95ee2ae22c52fe541c3d28011257af07790c0f1d8580c4f5c1d713298ad01519633afa22657882601f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha318a4fe409a4bcfa3b2e09b1db561829658a81523ef876ef446581c6415091cb507c6d073a866712691604637d0962af6efe740d547cc6620adff5e16ef132fba181733852be4eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h546abae083eab588286a42235f29f759d6beb656817ddf8e64df4c34e459eefeebd0b43737694380c0842032b813218c18e458913c8141de6b89a6e99eea3f9b86d4df7a666dba4d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd63d5eb9ba5764e03800a3ed07d01cd8e2eca5aea749f280bd31d2f9bc1ddd5603c1b4f883b6893ce1d4fc57e20d7dbcfdf55f8d25319ab19b48f96adfdd56d6423124faceea6fb4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd31006fc68b63c021f0944f9cccfa7edae6d39eab12110d17d62580cca5975c8c3ee0438a96568905d44bb06c7b122f51d12100d7685003301799fc0ce87388ec9591a75f40f7572;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ae633dd74a5b75fe95f5796dc3d1b1ca0af1e3ba6b7ab9cd10beec0d95ed95a36066a54cbda6af387df371301935aedb5f263dea0d79250c44ed2d9bcf8e562295c8b53a5e1f974;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55332ee8460f57c0eec5dbe2ff145010f245c4a07f12088b234d9952b52e7ecc2455d0b6b15bfef6fd1f7cbb5263a8ff1b02e3249705403cc3701363795602e08bcfe8de21dbd567;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c106ba8e4c44b58bd43784bf05e781a3f19e23d52c049aa447e974b2f28f7a974aac2e3e0ea147cf1bf2262538385281449c7da485bfd6e154485e4c9ff3069a33b8e933b726e98;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73c5a4305e81ab48c6afd4d3e2938354b447f1429d067aa871355b662dd9b750167332fbd648a8a4963047329f8b2094764c93df7a3a05557be3e44c9933d0da46c6042963468232;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34780842ab50939b2b729643e8326c586dbd210c917db1f82fa96575f42e231b94af9bb3f08dc8ef5e4664de0676cb6fc46ca5ced1527d555bfda7a51c50e0e4dbf0abfd857d6ea1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9a24a8db3bb6113d28ff278d2e4080b00c418cb427ab0e0639a47268dc0421a78b02ca376b174598bfec63bb1a01d672fb0fed8d9573ba106d20b2acc26d304d7231409afd44d1d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6029b2a91400b5a2dbe9695a6d548bdfdd130e3d3bd61ee57f71ecaa2ab535c5f30b374a2cb66fd6dacb324c76b8dbcee16728487a4249c2e6319adf4c33953814278bfb0ee81b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8096518aa90ace4aa8a44f460e36e1af534cac9fcc12209901c17b6b511559d370984fdfb8161442033984be1b3e949984dd1b71c2babae8056d4b5327976dee0eef272509981c6e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd347722436393c92141153aea45cec39b84c4157d8cc715448cd639eab3fb7bca76a8aaea317d681b0b810649e70059edf560dc17fd16b11399226bf89060fcd2a00bfe1824cbbf8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9393b3284db0b2916ac69a56cd991d9f3421b5bb7566a69bd1706b2d09004a34c2323cce7196a677312531d03bbb36306d2d471e6558f085bbd94f6f02d1cd805c42197687fc64c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd1bca76782eaa19f1a0bd9e99013967e7145acc8f620c1f643bb43d58234aabb082e0aa0753e546a92c7f8df341f81586c6d27432227ea5c34e50880307e3b7de0f10930f185d13;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h418ed73ed2154a734baa47543c7b90fd502ea902ba82362caed53a8d021f3268e03fe509864fa0f22a89c68d54a8376d9abff968f55ad48eb779380c3daa06ca5f963698a49d2321;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95f2e05f50a70b21ff697fb9644efec0e70b44b523241078402c5a6d0d6ad2f6397b45c941e8c1096abc732ecfb0ce9911bcf2f88de8f5f876985b91cc4d943d053e94f9f4345d81;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52aa841b98b140fc9d0ed4ae7830d65171da9790b0ff9663b511d95633e05e9d456453b564bbf3f00bda569823f28be0d652deefbec31302080a8c1acc7e2d938f029e83986fa24a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4cd86391237a33e4cab25e7b0e57ade7369c8e9dd070729f30a6fb03d71fe5804e37a2b33441cc2ec389122f08c6cdff4b97ae1e01031a29a5e49e0ff610496a794dbafe586ad657;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9dc8eadc08b81fc730762be35b76d94904395adbbcee5d8d9ed98671ae8de8c7f0e43e424b1a89a30a503111892bdd8fa2c66c1985afc374338fca74057e51c93e82f8b4d047b04b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb225dbc27a4c3fe5b99569f0371fbcc8e23c87de54c1cf27b6cf5f507191b1651b84ddc5a4d75374d6aaa01d24a0957d539559a4ce321add8974dbf011352a5d290096931b0c4c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb700fac4435f1a769dca8cb1abc5d03ea1263cc5308d7f9e16cccac716e2c1683af7b81445cdd39cc55ac2cc30c0a290f02e7a0ca76e69f040f1ae63a57d1094f45a03655a743479;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e8b428326c1336e17965e3c8de4913b8b8fafee140f34e2c353e1a341c83d41290aa1eabe7e4add761bae05766d769350b775f74a85c5ef45159e1384fce099d1848868f67216b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2c5b86973a38c1283e0572c0862593934e2f28612638e4c142f773457ecdddb93d7018f2b09991dbe7769ebca2508d61e90918ce1f89b35c1d5cc38450e25a1b84258f359565b83;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26ca477a41c25d298a7b294be9a0b334028d674544b5ba2bb665fda82557d5a75c7b42971e330c3cdf8936a7ca9bead73dd429bd2ec8ee57b97d4cc4c5f881f0bd53890b21e9177f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4eb114f06a218c9c74ae489245f10c95a27b61bb69831775ebac54ed352bf7269c3c5442783956a826b4d71ca69898aff7fcb4eb67bad1537d4dd4ecf220441bfd458b07c68bef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he52b43596218d1fc174b19f8dcfde96acc3d87152ee1edeba8297e69736af33c60ddb7f230bccfb44a6c793ab86e65f70dfa7cc338017a2ddd092521d77727cd5548fd45d528f38f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1603d13509e7ac1890e6b7db5f5c9405a416ac97280a7c22da2611ec003b7472f687bb9c8edd2ffca15ad545c0915675286e2c815ab2e92ed5aa4175fec9aadff9dd49076d6677;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h866ef77420eeea096af4a78bceb17764f3f36015042477241d4a94f836dfdd2cbf059b9935439cef1d87da549cd6891e9fa552d43fd901a8f57519e6df206688abb4e8dc1588d566;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf42ce4d84bc22ccf0f205e8decf1efe8eb7efaa6958fb257d961130c2d4904df23a8a4704243bd77f0c40c58bcee105a96537648cf9c70dc720332381aceb6ae1e441d334e9cf133;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9715bc35a449b05273eebec1335b250199a4a3c2e6a83bca6a2f534348421e960f81595e3375178a8ec8347029a012ae44acb571ac60ec40036043d84521eb5502975ec0fceb9222;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f030b0fbe970d4e90dfabefe8cc03bdf3e98cb6e2593816817b65a15c384073d820a23f04ce72e31f9b94773f52e2d2402dc97f36920c242c0f05214c5b6c76e697df3621f28e17;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0ffb68794e2e79c088a9a92effac2d923ed27ef1776515bcc22f5915b33440ce615078642a476028b707affda8e9f00ee3ed76953d475ee174dcfcfcc74aac3ca8773e759a6edb9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd70c0b672f96d9982e2d5783ebbeb946f83c6fcb7a196d80418de73924a33d268f871ecc3f22a53e50ec66a904dc223e7ed8ce98533c5bfeb2bdba106ef23ca5e4da38f1c357f0a5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he0731ff451a367620d90d7312d53001a13182409f21ff451690c19cdbf0b73d6211eabd898d62cab872c089fc9b12bc690d3ad0aaccf27dc5fd8d801781a83f81746cde7e67b0ab9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4767e9047c3e2b63da5218864d893b8671505b9bdf2cb97269b75e37e5222f46cdc436f90cc145fb073744204458c7cb1035b77c24aed45a1f76013c32cede84e138104e731d91c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17191fbb6215e00b356d190109b2a034a2a8663306b54789f3d8d22aa42e48c130951fc5c22e5182339974a36cb3c7cfb19c6247973d448b1a22a91f25822e219ca308e3390887b2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd5cc3b227a69d908e1d8cfe6441de48a9865e81004d439e6149c90fa2df199f2588f0e16bb6633c36985aa0e8cc2127d710fc1783204838b3c1bac7f9da5680304004f0660cdfb0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae0eed736142d00c4345448e3030fa64380539377549798612d3be9154c5dc5d9aac6db8f344b77f39c965c89dc8a1966b966e7dd03434b2572461018a60e16ee553825325eef53d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb53ab070a1d5ec6742d1a3853067b378382dfb298f82229b43c296cc72208f9fe12aa3481d2f81f77493562c2ce04e7cca01305eba1a3b9704be66327f9d78ff3272d27610caed61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb36ebf0215fdab3f4a874cc78b2d2e6cbe98ff3d55882c0e77bf39fb37e21148ad01d9ce198618283ea47cad5cf78673640887ae758cddbaa15bd433adeee437d18eebdbd2f8d78d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf42d0b513a4a9cad20a9acd32cd10823fc08a6cf765607a2c6e0dcdc06c8455e902eb528313cdf663fbf74d162ac14e35d812bed89e519b5d63feab1fc9ee15ce9507e428818d13;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b65798347713e5b3574f942744b0b21b347db6109f3ef937a74dc19ed97679bee2abe0e8d1208d838e236ff9eebfc1082049aeb3fa9e46624458c1971708f7173dd9f75cdb40646;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0212ad94065635a03abcd1766fa2940cf36cd440cfb961728abce7d7f96a9508c8837971aecc06e3ed0e521fd366747a4d39ac08afcef90306bbb4bd68a52d2c836be6b82019dd0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5698f343acd163c55d20f8ccf911ef62e8fe3500bdfadc7e8c7905255a6ebe505ad41666c9acbd36473cf1ef33e5e21325cdf243dbfa0bc6b72399f81a0762410bac5d4043ab09c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2646b8e5f31a6b9f313a3539f43c9f062d58efb62a2d800e6edb3ff09eea67b01f5c3d238f570676be9b5ebffb39e4892ba569bf6cb788e66de3a019bb442d0e53c11c13c406d0b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37ea4a6167750363a6416e0eacdb4d33856f1848fa985d269a8c66cf8d33aa455147a1dc45a901884b709cb7298c95541d0f676b453fbc244728b3cd40ebf2cdb2630aa03fe1a875;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51d02cfbb3dd081b18a5d0ff0585a1dec3599c1f10ce1d0f2ae1dfcfd42cf2f67afea0e45656ddb7dda60ebf38be1316578d51f8aaa21842f78a213fd2c0e0a0bdf380368d06f5e5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cca73fe039767bf91d73824b2bcbd8d67549a6352a39941d30bf7362763fa0d8762f41752c3261d3ec3741273e51e10b7c1ba22e7ab49c8229200373f8af3d9b5b2d8391cb39d62;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b25c25659a35b1b3d4c5d2b3081d09b8990707038eb14a44e0cd3127101405714ba31c14890e6a79e97c1a0907a982824eee89ef51f509dedae9ed70083995463ad49ea4958b3ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h743f4dc53b2f24130f6661bb578f1396317bd7541c3f0083a889352842c900c26573ae4e3948cb0c228c7b78885db6c1d574795811d0420617f25c3064c94a36aa04c4ee57ba063f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8edb30224b2433e2fb54f9c69fe7d08332fc4d3a900a611677ccddd79292ca929c1013d61cdcd39695c017c10513bc351006287676ed49ea4aa8086ad4c8bceca691697b9a70eaa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81a9b9af16c2ad69d1b078fd5e49e1e95ce924c484940eef61b18507b2670ba704a1f4518ad930f1344f7e83b4ed5ab065a23f342f7b230dd06149c2303158edaba30907ad0935ed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h556865bd44414f330ab79afe514f47e61695532ff3861fdb910ca132832c836e424e9a9f7a3bad0b62d5cd2d5bc64d422d6af6258080389b6d0a7a8cef5be418437342ad9bda7a68;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1c7ba4c797e4d49bc3f188e2c5c7409536ac4f9187aeed48763938c7a977316e1a79a08b5f93358f39b62efc57ebb86a3b56473b3e15bea659c6fd8d30ccbe4e42b0ba8af027e2e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2729c24b2147ed4b686915d55acc142a4178577495d886bf107615b2e4f7ca9e1ec9fc8a6a2c64c89f300fe9edb2cc42aac981ac0dc4ead325765e902511c1bd54baadf734061eff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4628a67e1b6ce0375c69c5d39b15f0feb8002f1d7e500263ac8692c4f69a237d6b92fa5146590aa814be0499b77b76f6c6b344526e0a86d37adb03b46702f4287d401bd4e2fe66a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12d23d964e83b2b3a837d81b26854ad42b05814abf9d090f6f9c434807e8d74395fb494d4284e7b384f44b6e39554fbd9cdade9477f796fb6ebd62cd57c5a173f83c1c7587e35387;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72ebc099e85f1b5d283f632e83d517e657a8d42224fa87200de58561276a7f846eb651d2bdb5a283c1a05df956f69abb0b7613d66e62754b2eb1f7c5ced0ca52407a5b88990e82c9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hacdfa1c5b77202e98677b580d5fcb19dfd1364ba052d058fac79a39c18c2449e271b3ed15d9053f6118de42732d0d6856048d910e4128b03b53a2ca554f055cdd4df0228bc6d7d64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he12d8eed2b37252154aaf552dc34ff8987ab2cb7f88e032d5e071018a6d805bdb2c26563aee947fd2d53a64c157c7765790c4993fa281807784895d553ac871cb9e8d976bbcb5c6d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h423cd61a4e888876efc8050ba12674c7aa51c9813e83df0f37a6eb0cd40064e85035f2a11a965e15d90f92346606a3156da92a820c4730336c3af1a8145cd408975d66840247b2d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha540f8e6d5f8ac9dfcd2976f060b637bf231348da425852ae6784e2931a94f3a9c3b73e656d31ddaea5cd55ceb92081d094b296875cd433e57f75cef437c77a960003652a35fa4c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90fe1d62ab1f8004e5c1e50b06e5936b50cbb4b795b66cb72b29ee204baaa06d899c2550d4ab7a9cc80c673258a13a29899afb6f6b71d782d217c2159c37b0d8eb4a7145c05764a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51278ab3a374ba7677db848c8b513521608f3375cb9589de4a31fad531d1b0c3003b3c90c942a8b44abbe3eb61103f499cac60407c1130f887f83159e83a1388a39d3b495a4ff7ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4cab315683b2adf26f97849efd9590bcb8b569d325a781dda1ded3f746a36bdf0640fc2026164a4570e37cbf29599d78bc6371644800166ef5f0c3a0a6a3dc3f51d68bb7a25b478;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba05dd3c4cc24811ec1be8d148ee6b9e84067ff3b2da0c4b441d3c4df113b9746046088ca81b07abfd995f0f84ff75d22d4bf41eb50bb8712dd3e919537c0f6196d8c2b0020ad644;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bd144fce90a653ebe44c162a305fd9e8aae6621109d72d187f1c855e4a372c942c7e6379dad7f9316146f884108b243d82e3fb7f106be1549d6624fa055d229f6750e7b64c9cb86;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc7c9040f83c6e5e4957348eb122ddb1fae5622ffbc5433a1e79fce40397b987965a5437219081f5e3b6aa8bdf469110572a0570d3232583db44fa8f4bff2adb757771bc87f540ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcdce6da9b648df668871931d273d8b4066d193074bcf75f126c56b4a0392f86b42f2d5b9b8624cfd376112934e0d9c3d38ba8b6275b1b5926342f187505dafb2018249890ed63a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a468f1c906c83d1b51ceb84c47bf98289e98e9be61e863cbbbb1f01ebb40738802181c0a38a3a714882ddfdf07074f0d73a938944a1f512e011104a301b8782c3b9c5d72f03c83b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31fbe8555f6575295ccb0e70cfc4545f03ef8e5ff77f4fda8c041766ab514b44d3135da0978efd61b22b8c18f3a280f04038ade0799ed64383a5537b96374e9e77ec752767c9d1c7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42fe87d83c9fd6204d9aacee60c8186ef611f6691383bc2f7dacf68e37378116772c5d0501571cd3f9c4bdc6250b8418b20a3378ec01b13af3a1e3c4ae02e5e490470e8acad2eefc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf575042fe45cbe65e3e05a6474129b68a02ce90a439175abbba076c58bbe97b6067b58a66729588675ee8c66474109ec334b1635e64d0539e3bc3604340a91410dd8e1f5ef4405cc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h816b33a3b3e1686d7af96b17d38a9dd82ddd8cbb0a803e215c44b01431924392205ca152a057e5bfa34e6b1c46bb3c25d5bd1a07f9408f8f7dea7692668cab925ff23b9eb4670ccf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b44ed5515060ba844a21f745774db43b3a408d6fa810e70f6ebfc3f31230d41a492a69955d2358ba9055ada801b042c024c6b297a2e3f2a86dfe412bf277af9f12d53406d94f375;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9191c28f3c0213e80a0d047f0f18a7d1822d0c4968140fa681a9445186ca6a5280e95d3ee44909768e01287023a8e867b98c5ab6da851675a9e641074b286ba8e2a630e2088add5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb728c8b7c6fab3e4b3fe143ce369f818f37a727f14bc0ecec25993bcbc94a2e0643eb295fcd5f9c0f0c1b973156db5c2ed577ece8a321ca9e210acf6b264e19810acd2a23a21c87;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h204be2eb23acbc6270ccf7dc4bf8ead330765abb33c7a0e77ec2797e865f530f7e4e1ac95b648f361301fc0d20d89848960b92d4556d6e12b90821b718dd68d7b3acb976ba51dae9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf281a2429d15043d124f267beed29cf9e292fd1e61a49c7d934d325d4e90ed1cd146f73f93e3c49ea2f8e542888214f9601e50aae67ba6b7670fbc85a05b2c6f3d06c329e80bd9f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc50e88dfd1b7795a3cf8e0f08854d29dd419d560f877c7f674537b6728d05ddeb0b30dbfd8e38e973f6b24a4cc5927b69fc530d278a60496b3a02af04c2865abcf799a2048a4f4f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43aa25a0cd95dd2e028ecf003c1066333baf04edabae6d7f3f05d7c5c8462d4c95ada3a5037d6b089e431b76a43c2391c39b4f723dddc732963b9a9afae0043e285a780d79d20ae7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6b0c6bb3a00040a85cd51a0131d629038e7428a090ac47d6b170af820061b5dcaba53cf5e19caab60bf92ac4f2c659eeec9738bc4328c85c4361779df595e5ceacbfaf47742fb5d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ad1490204a128e76ad8c80d9f3476f8b368389a0d784d71345184f123d0ff0a5ded5732cc0afb47f7bfaae46e7d6d96345165c9cabd61bca6bb32b9cac7f6b50f70f6fc8b567227;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21c6188fefa92935fc9074d024f8414b091ad063f17035ebd7cf9af6c4029221d12a77e9bd60bbe3ca94e713d4693d5078892e2fd47a23d5e49d80837b33ec360adedc6c5d8d032;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4042e09c9fd1af75d172ce301ce6fd8e1b09d7c18df10265ffc4702dc10be330a30e19e13bae7d1f01f8a1503e05b5b1e30bb65ef2941ad2db41a58ff0dc258809c849d14e04c0f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fc1f6ea24935afb6a2aff07d8b940c105f2559afdd93095325172bc60b0505368e6ab48785e61abcca899278a68ad805060afeda135f0f65b234a61d8071480eeb2235d6cd8f466;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64d76fda2055e5d590ae3809d46b55a3d7c8a4fec0b5ee1d63ad428ac1f9e3adbe710deb33fb5a9985d9ec65aa43463e4dde85e23cd4964e82ff5e62931cbece18895695c9b3a4d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65d697ba50a5e978157f97599719e52b927be47545184ca01714fdd17a26f27d0abea43986bfdc27248bad459f731e8998c29c4b1e90e0dcf6593fe7683dce45a02da33c6a583690;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4806be6ccaea39cb794e706cdcb3bb5e72f720f90aeced00f51302a9b1ad7fddb8b80f2f6617a657c75a18b39af3a84a9e9783734b3582d5f4455d41aa91be574500ba74c1030324;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf299d7b5e11958994db66db9600753d7bc4036c31098d26682d36a21d6f26a0f2f341439377e79cf467068ee7bf495bb3eecd1f366ba57484adb6f64ee03e8fe3498d892b89824;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a32ef92be01bf1eee02b4a39a0a4609d9bd717f3ff58ce19c69983d5bc32f1a3170bd096007314a5e83894c7c19d8bed70afb9812f757f50054e76bfcc4148411096614fdde0385;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h815895502c5bf59e363185819e6ccb6836b4f8484648b43721185541d4e4696159e7c27f26952e9b999a91b0e3026cc07ad4e869fe1fd4cfa481fd84a25fa4cf757a9ee16c9c3394;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd87515fa1312209600e8cff46754366f5cac683e6eb139f7f544f8149dd8f4713637eaf001dafcedb3c83a79dd46d227da4243ae36c90f60a1ba8375f275aca8270ff5a96554b4fe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h481f47cf44615933ffba2fc4992f06f6897b7b290fdc59a0561d18993d8f0d467f8c258337908ba60d1edad96cd185524cfeab98696c5959d1a6652d62e3c435ada652318daaa60b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6f56ee99d3a1aedc7c419f76073e821c3cd75005d387fedc9183bfa6f2b3645e4ad5237960ef708d37468ea4b4cb15e6cdd6d0865de114bc1fdc19e411cb0f1a5b83bba62e8e8ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he090bc93af63caf746343e242026985137c04abf15a7fcf74f877101cf07f2d32cefcfe54b6c6bab93851754ccb763d2771825888f369be606a5fabe5249562f974abb6fb0f2da7f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b0ca802cebfee75be16634b88a61cded5fee5dd8f3a07f3a3d4dcc2822f0f0eadb802e8f4fde8721b4ffb5ae96f2d93dbe376e10f64b6ca4af7844e74df707b53ba27997f0d679a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab409f4babb6e4c2f465b464fe42d7ea22fab1c57584b5e9e0a1a8e432ad90ee3e2c5a265754d1d1e80bdbb423473776ad9b0b1e6c5e1acf123492eda3ad0aac9e49d75c052e26db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde021284ba7cda3bf23f29e7d231564cea164466431965cf16dff3599c88360a481c1907df6744a277bd06ca9418a653c7ca9d6af5f4fc0c2769cc5f0281a53cd527056ced01c1ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8be28a5371f7d2b37421ee36de4b597eb480347c760fd820056da67e4398d6c3359e09db6ad6d251e0fb07674b7fa9651b7590408eeff353167e22c1aead4aedda2236166279817;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1eaf6e974d9b32bb57fc11e0ba956ad66531c73acfd210a43a66536949537a05c5819c4500ff86594855d417dde779dd8176c6ccd568765a35e09be8362e4adab63a3cb743f80e69;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14aaa89677fc022ae2fe1d6f7d9b5786774f35c0c41466a30a4353c3bbdd76bc202df77dc0c87c704dbd8eb8c59971c5a1c2cecaac4cf685e24a05587baf5e6685671dbe1a6a45ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf474eba47a7435333ac2dbd56ff2b3e068d37d473de36362c21fb15ad9c02645191739956cf7c2a8d9c57f04a2badcea7fb1372b2824301213dfe1389804426799d71442358985e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd353e58689f06444fab08e462d9d7a8519f28170c286256b7c7378023d89905e195d1530000c6eb323e9df01ab2fda6fab94b0cb6a46918040f7a95ea80593d301ac108e7bf7223f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe1058305e47426e6af5c53473268a27100a2357d6710c26654d7c8ccca264cad1624bdc9864a9dbe4e41fa7d426a3aae56a742084cc38b118747fb948298583cfebf2e9e84d68f1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdf62eee2edb977db9d75f10658894da7dd16ed4338123ea545ebfcad8209d45c4144913b07cf0e657e2a6deeb92dd1774d21fa163fa560db18873ba71643e5442469ad8693b7aa5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c8ec5a3a4cf284f806d8c795694d6e24d3c28a381fd6f811b035c6f4d21be0bb516c74bea934eed85848b17f794c46076d05fdd86df8c733ac601dfacdbdd1e2fbe4815b846b4e4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63977bd2afa0f087aef75e84404ae372f888a4a22af8da176ede47371fd8eccb1f437c19e99bb1f86b343e915d39aba15da085018e4b1201d6bcc266e366853f62a534f0cf321eea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde2bc364e145d05cb39fff5c914fa7a787e8a51da583cb4a764487fb20df46dbff0577aa8223aeb5b27e123b9d03577733d8aa07c8581d6b1ddd73afc68fd1f194aa1a68f69278cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h325c1f5adb7625178f3da10c03e39e2593da0e39d4827fa864172c361afa5c3bae104dfe54cd6dc172d000dad4844b9d5c8e9a6061db6712d1ab632aa886264fac634befbec7e193;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2857dd69256726656665525ad9bc0266083cbad901fb093cd4584ff652943e2159ea3c40d8b614a482f1080714ef04e4dbdc85479c0cbdba57a51002d542cf89a448c5fb5533a47a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3199541e56d0f0efdc4596cc44815cc84a7b0489daf19a9cdce09872f6853ffef495fa5e4d2797088c09bd559c91b8cca3b4ba9e3ba4ae48ea8ea253bd13977c463fe128ed79d340;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe04b85892fcd7c83ae68b1e594b56d6ecdcf5a46308587ab59f0c3f1cad8a1886a347045f20e2f2e9dc7ee081b56485c3c656f56e55017f3a72d9af78387391d6b1060e87a93881;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30ada424654642c5daa859a24cfe06d443cab0103eb7c67fbd672d44397906f754b60ce8b9505a10f035756402706454e5a2154e10d75321978ef0a2ca1224eeb282364331733cfd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b502e9ccc3ee36725b426b2cf98d7b6515b92168dd600564492f1b709433a34589aab09f91f784cf67c4a936d8b781fad51c864822274c24c267a7da61b104cbfce71dab0eb4ab4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fee43d9331f0fbbc27e3f95105be106de46a25083e5fd1796e0a8b83a2d371aa1fdb056b2d15e94e9f71ea7735497676a9d0187baf3f12ff3ff47c1b3c4545be4a7bf318386fff3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h354e3901c03550a9b27cf7021c5a905d297e05889dedc507d5305ae66737ff5d8f7a6cdaa41e9427f15bc2b6e8ca5b25ce11452930ea892b7e02cb5b3511a03ed86f931f7ebe2d44;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h135bf91c539cda00be4907de829576e44bb55955777c83d81f9b0275164abbca6421e789b9ee4df76e8ae69fd5480584cc409946d517a3cd67ee3c9a805bacce19e102e89ad5bfce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11cd02e10abcc783a5d1dfd200d37ad729ca118ef9cc9b15d9bd7e133563aa4271bec1bb311db9ffdbd82637f39107fa71e8ca08493a06ff0ebaa6c4609f04fadb863cdc090beb1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f25433a0debbca944b05b02c0c6e8c8434c86abe883b8b478df786122baad0d6b7ea1d52b6f360a451c57654413de556bf5f5befb5df0d968d87bede85dacc7967149cb2e01a86b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd128872b20e962cf95badeb6cf56fbe3974cabeceaf0b69414b0435ab518d55707c0dce89e205172685f42c256535d779f9c6ef68dbb328d4bc2bbb6f9d0b3553c11ced6fa1552ea;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5fc6eb70c36813c5cef00147fbc102f738446cc498e301ce560fada45234686dc7a5aed4d3ff86f02b645a02e00d0cba23b507475bc6c4276cad362c521c3e7d3293b591c443f60c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc22289625d8f4985feda33f2d7da9673c625489c7ccff9a1bc61f7ffc410a2b7c011b7157e5ab62298d7faad9f4ffdc67e6d2fc2a3af088059d58ff1f5e4c7d5f60daec141a33a1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37bca3538dfaf54ac98432846cb73839e813fdf6b017c1dafb49682b0d205052b29d4eb3863cf4e62823d80b0a0911c8ec04f3f8d1fc88370fa24b057555521ec071e54cc3427921;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f9d9eaf651f46e1e1517ce9a359e79d75c5cd39d9c0753fa320787eb72fed72c7efeb55a52fd8fc8a0330d2ed68600668af8b33d01ec17ce9253133c8a8ff80303b99a2c28a4699;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce5d2d5c73080b7431750c03ba82bc7050675635fec42eb1afaa452a0f9b98f7b640bef4ce115fb9d544b51e11725364c0962c72ed7ba95714dbc913c43688c340aa670f871371d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb22c097f5e0b9d2664743b5ca3fbd767d6fa73dfa41fe898c2af8d93332384c57ac8e363c0cf8c371826d445e3ab8b4f72b045d279b8f1bed8877082bdf8d067556cfaa046a39ce8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9cf7a03aaebe16b10acb15bd6e5c2ce69af7d7cacf4f4925315a7085daafed62aa6f949c3dd33fa8237e8fe8dda2f2dbb15f11624b8eb12aa63646504cbcf7387bb52fa13cb4814;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4fe604dcdee23cf7a401a3e44c236846c6eae17b26496251e924c317abc69cd3b13eb39be4b8166414a697f9305d1c82adc23ece3f972d611f0e4a7b91e77d097643a22c7af5c46;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9180663dfed6c3573ea1d3482d6e7538cd730cce50a1064eb782feaf473cbe1f7a9ff1235cc7ddc0c6a0e5bffd982140712c2850a41da8fe20ec57677387047813bc7599aedffbfc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91ea7d82081ee005fa45cf71ebd9f28fdcc0be90ea642972fd51af91647ef0adb0062900f22910f6b8683a5352e6748e7e3b1d95940ccbfe42fe1c28ca782d9e1e9198d3be271663;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83fc6c137ce89c861688ea320cc7fedbbfa4b69dd4d30dc8c8cd05aa5684afffde38d7b6df81f22a66a5f961b523a51b5f73cb3eb7d76c48a06b3dbba582181644696960f4c7b867;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb6d1d1e4317c4dc7c68621f8d09f6a40360aab5efaa5770532cf3a586cab3b6182990a53cad82e6ae55914236fa43020f1606617bbddf21defe5c8664956fbca4ecd038e849a9e6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h323f762e2314099544a2550e159ce9adf396a6620c94ef1be6681febece0f8c9dab75d64b6edef5884f051d36fa2c98ac18f213d68044ffad76efc76b3ccf1e6efcca79a7d6e8ac8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27cad238149a80a7ac0819d836641ab4f9d9cb0d2713fecebd16a6f7c415aa3c4beee9cce0d577df3c96c0207c78d0d3bb5dc51ae32d1bef8a65bbef6f0c272cd2ff5a18426fd0bc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he60f3949d2e70eca3afe4f979c10af7b044c053c7c917cee2df06980638a7770b112364992a86f7408930c056501c62373df6188d81ef2ce1a6e81df3d89c8eec64dbba1a025d684;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82d65b27f6c1ef90b066a572573e690db47d078452c0a3b1b8da42f41f102060862bd42c8d6554a59e7e732f8357faf2ab60a84383127c30e24958982df7780aa77d680eb020b410;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3b0e732c061ee022778eb60eb6f871bd6c09155df94b35fffb553f40927e4afd2c05d819d7ccdb4b675697505f63c503dee14bbc8d9ee4fa9026026ca8bea9e6be200ae86af0383;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11ca6dc9b4553a9569392a79751e7bdf1083ba7f233f03f65b0dce7d03dd7fbf619ccb9bcfa2ffd1169c4a2849ae2307449c349eaf400015ef402fbf37d4ca5e7b67649e96f3db5f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f81319d6cc3cb98c942ed53ff2034c604254a035731fda3928e89024429a1d249a10eddd7b4750249bacc591be24b3aff1eac754507646fe02fb38b1327092a75303f432fdebdf3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea829e61d23efc3956a97791024251c266a92e4438580cbbd05480c008638ee752fdaccb32c09f581c58fec52339cdee09e73d9afddbdb9186cc565a400b7802790af3dc0a8c84bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a93cbe4cd4d4c21de3309c5f9dfdc5a73c3861f8ad68c77283a89f6d72a2a2eb59fe734bc6655627b5180f6cbaf21f3a7ba4056858734f385e595caa3274f1f2161e7b190cca171;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a488154532d3fb6a1a6c8e3bae65c30570e7d9b019322719286fc7dbbaa39a7e87d56a4b300f9c70d17b8918737fa1336f64c8b8fa87366a99393e92f5d342b73a01232d5cd8afb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76bb72926ac57a63c30a0d833ec107491454573a96e21fa4716ca82434db1195ce2677b5e87bcf5e2089ae0f6e9e6507e2f6caaca97fe8d287e5a2c6ee371e2efa94511abf953e53;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc66265109764ad3a309af8e363dca059182ae8b4c24467f4274f310fda98258d21565f0e1780f4c3faccde213d0f220a5e27e04d42a8f590c080c4c83308316f0d9b46f742cc935b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f73eb6837f69075291f8e1485390fb5d303aaf9f9ff077a7d7235c070d8d3685a6f24f20c1c8633c848e7e7836660d8b3c4bc102b739bafdcd1dd4d7edb62315dc9d2f060703f1e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8af58816bf4f08db3001775c261ace845d363a7fa8862ab29edc18f90cf2307d2c77ff278286ee51706b19d880c3f4970804e5170f65c9a8c92b9e864b6f793c760e01d414fcc3c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c8e2d87a9ece6eb6f3f5c6654571e239594480dd1726a3d952a0b49e7f7b6be6f2a12da1dbc1cb856196b4b9abb5bfd0cf99875aba72692ddaf1a1ce9df5fdc3087c196d90a0826;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfea18b31fdbd0ebff719ea6806e94a2827d6e49c5c50a2951a3cdc86b704af9949c7c73b6afc7ab85c3d73f33b4a17b183124f538af1430d04d27afa8728d6b8d7f758a23d5c7328;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14d4cf013fa2cff5404f5379806596d8d772578940e9eb114ed5e3e9236a59976343de752f363aed252ff7b3fc12c05dbb5b3f8c204170f7c439180a4cf7dc871aa0f7e34277a141;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8204263fc9c1779cdf1f321095b73d0fc9959beee43c8a10b3bc15ea37ce58262579bb1996ab6115b0a88dadae481163050933fe754d46d780cf1129b7e7b8b3a2db61624af837d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63ff18d026c3bbb0b498933a7f175ceca108634058f90f55f1d0d5db71a12dc71fa2a5243b27c133379e10bf3b45a4885780875d7c933ecc95fee956b6fc90e92704f2e278201125;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0837d394fef18776bcb2504ef8c514f5345b38a9002608134bf95748352df8e762ca1baedda2f5349b54567daea87d30a61ead5e8f627304a10949f51dad407b7dc0d67b7df223b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b7f430f7566a0105fd35a74c735574096e009f141b9a2c612be361dc97b9f00e84921671100190a80be65604f6f9b77bc100d77384f535c42b7ae5ded49b147e59e5e8172f57b72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2011c615c224696f090edd4a2f454d0e703f0ed273562321ab85034727f66c89e47ccd3c8b185fab1a672741d8558df96d22545f6bc509f3a4d544146586fa7f04df973a7018e1dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcec4e19e8ae93c35fe962042f90ffcc52a6ff48683c29523b7244b09956e65d099b17f1d9e77442b07636815fa697e475a965b41259038ca672c3f80264d1b3071f9edeefb752f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h529f97d4586f7c6afbda01b6e160ae8804a4cec0706ce2a98e651b2269e7834ffca0e8a8c5c99d517ecadfe2e19904f48c39777bd92c230db71382b6813c17d8a23c296dbb5f881;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf050431de676f89b6551300af055279fc151f793d23ca6dc3b8435d987ac50e517e195952806c047500de7e590da1809bc3aead4879ba8d5c91dceb1fec75c7ef4549835dd85f38a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd96ad9e8a65c72380a2f4cd6cda892fd6319c768dd488bee1c2408a6d6df2a2f3d45c4badcd31108d4510dbb20aeb24ea7cce3ea61f9db16ff2afe26d30670510329bf64558a1067;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5711583752dada527058ece9045b72d1deedbc6527497fc5044c0c8a43322d6a61a9c69b65e8f579f182eec5ad147c3e511079ccf94f5b4e1aac79007067a6dd8ce41cb01c4e5ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b269782b4a6021137a76343755a7ec1d06debac240c943de54d44338af43a8d2f4ff8512faff130e8b89a1814e9fd771083279c606831df5b1ca65f4aa8e11981ce8d6dc98a0874;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0318fde46c79f56661e46b3b31771a4f1d270d19aa8d155f7ae0e5c102e3defd2b0b9a3c18962048cc40af4cf0bd290ea430b4a30ae9fd9f6bd74ed881cb2fd78f69e74cb50914b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b5d7660628b950b4e8dddd44613f03549eb4352e9acacc9612881e8e7104ecbee36d3ad52ba9666dac400b6f95040d903b51d0f0b4a5ac80b0cae8adaaa851683cec5963f8530d7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h818eb8a04520eb3220cfeb7fe77e5f5480df5b80c69bdcd8c0227f1d5ecdf37597a474196afb8a510641a34730c8926ae8f88c512ad5c9674d27f4d1548bc46d3fc965d2332beccb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58517665c744bdfd8a2f7e98c8da79e8a871022d658c59f5b2d37f58daf336229c265daeedd5315b307f3f0499528436695265892f2cd90ec3170c5cf67ba3e15f571cd67272ce10;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c966ae8fb5b7e3b7de6262e1f188c8162a12d70bb367e0b011379836568ea79c4ebfbc9cc4d61476d41e6d7619b89a83c56a6ebb614653dd23bc6d233863a7e7e5e1474685905cb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35a0ebe3f2ad583e14ccf66997d078523e665d5be67a4e734901bdcb780785a97d2799491077afa4a55ad29f80730a9c213532f3e535b5009e18fdff29bd625e9bb10d52fc2738c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a962291b7da2f0fd453534c4e8443beb1fed0eaf13754802bf347fcba991a08ae26e7cd2c4fc2e542b4042e12da0952a47424f30838adcbeb9aad17a5bbed8b873a23d0a48dbc5f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7db592eb3c8af33435a80f1eff02b9f291d2a5894d58800d4e54808a8e4e12e020f8a417d30807a83f610e4ac8497dd4c3c71b7048cb521ba26db7ed4eaca546f0613f15cb8e313;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h140ba4270d19af94fca88de17f49ffdb7ee794630638277ac50862b43833f888dd64ba56e712116edc4e96cae4ab18f5b74bf51e5f2c7ef105a031ea304669d2e4944a1b4544cd2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf89d8f9143c7fedbdbf607f108e363e7ad2b801e503d6f47569a01451cf2109613bd1309e7eb21a87688ed8ed8101d34da774a099095146b2066c5dc5f2d346f2d72ddade0652ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecedb0d4d8754921edd9514c076da3d60c924785cdeb152bda4e60dbaee8a42e1fb7e9b000e03bf2e6ef00b90445ad161b5209f4e8656393de8618facf110ba0b2985f78652ac122;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb95798c9d211a0d5e4b817fddf35fa0d73d00b29f7a1869be92f95992628117c151bae917853a1a429db648e887d0735aa8726aa78c28bddaf3cd09e8ad0c9155d6cb7042af5069;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44377994e1fb6b54b638b1982a1e9ac88daab03df88797c7c01a570f18b328cad8239e884fa5681e03fe345aca459ce1ef8c64d613fb4ee667b752c4dc3cd14164e59f97bb073097;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53da9dd8869317721b63051d25bb93f18a411a219428062bd4635ea9f79c2616f73c60b604a404c500b2a8553f7f8caf30f4cb908b717e8cee08b46db300d7b5f1103c684990a68d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13a0443243eadbee3f9c5de85e87485c3adf050125a462226e607115fc135d1320de3015aa346ddad2791d3bdf28ad9b5fcd245207328c6ef7a6ac4ce699913a87e68d75fab9507f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfee77d157f1a704f841c5fb8c2c0bcd9b96ad2575a87d403fd9b42bceff893bbc20883afb91f412e599818bdf52eaccccc71b49a00d42cab3f4aed41e4ea1d94e9a54c56558468f3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b48a9c86be805642bd182b37023c4c5d9fdca36aa746ec123577716fb44caeddeb7b914b251de7d600c8ebcb301139e2dfb9a5f48b932efd69deed41c13b4bc6c2f3298df98eb4f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd65c132e4f421c01189960e99240e838c08caca360e18a996f3f152c7eb69a6acd26b5ec43a74cd1e01ef3fe43e292df699ce59295c020485da1bd86ab95db915935fe5af1606ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46747afc62cb0cdc22064215a9efd3282e24a4076c88aeee8f028172a167ddd1df5add20afcc4afae68ccc85cf05ba734c76dd149438d43505781fcc6072258e7c075a771ccce80d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52b82f39049755ca2084fb17ca886f8d3d03ae913db2b003776ae610789500ff29c9266e8742ae3a0c3f22154a3ad31261e08ab1f9a853b3a8cdd704370e5c4348e42434b000776d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2556cf1067bb7f1bdecab26910acf3357889dc6767a728162cdfd9c31070cfd721ca81dcdef377fb1bec451376d64dd9f770bc3cd56a7a7f94f198b7e2fa00498b4d20cb91d5238c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h430cee21cf408923072f49ed000cdf09e3620d07d8de8f7290a644621d6d9850a1b5de7de8da283cc045029de465d52a7b4508222d267607895913b72221101e6088f9c3eba9e88d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h639447953cca3178a45793ca4c7056e173577152ce48338f75a5a2647ffbb0532ad6b86f75bab45424e6ec7ad758dfec760bfc570ec12122ef210ff79f847a0798e19e742c456f4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf60bacfb2c3f0db96abe99366b20c77357011c2332338f4795e286eeecf9cf63d2c807d1900f896063a15e71caef70a02369db8bf84f2f27a8334e00cd472fddfcd2e75a5afd313;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd18e66a931b7128a1d740ad7f1f0b05a982e160507b84a2ba06f37a138b3c4732cdadfdf6922ee0630c56f8a0db01605609d49bbfc51e2fcb0ffd3b6e911dee5cc35d2032191b303;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ca33e2345b054a80cb01431c7e5324c97f7c826583f4df3e375e4eb9c9e1bbc4ca0acfbe936c291c6a68ffa12dedf1ce3ad8dffe22666677a72227ae1533c062496359dce82ad62;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc00bdfe97eac3871e511f60e92835e5341461ef5601494acba1415cc60aea754a0ae9060355c9b61176242c37da5634db2d099f207f921178bb421e1267386dcbf686c84bf03b10;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bd7c61d738941acf39b1fbbdc0302531ef6f2ab080d768d6d374b93a24528f2b59d331414efccfa1bc299cba3d4d40e3ace0a5ad3585f5be0e8e98fb38b5de26b414ab7c8e638f6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd492f1d93ea86c010995cc5e3a5b19eabd51fee38ee9f98702e5be83166f31f76871b7a087ef85f0bc0e4b375e2ae34840ca341fb97e2ed8dc2980f39173215db7c2e24f1b0bb20c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf99de8cb5f89ea319f236a54e5b06f5c89db6ff45c64079df2a8aae11e0c3fce3dbcf8220f42925c0221c0c0ea96189cc315313d7055ceabf8463e6b545d93f6d340d4a8787ed140;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c00fbbc518bd2aabc2a2304e0411b4c16370afcfa0e3f58692df59a876381f8dff6cf78f69976772150e5ce0d3f16562268fe7d960d7dcb3dde8b2c9aab2acb4ae720b8ce5a20df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h478c6a8e953bd7457fcd1a12a8a9c0651dd5b8b1548a638dc09173d228a128bbe5a6a1ab23f281edaae4561217cdb5151a21d179d3c256eebbf4a41bce2840513d9514c180ef7499;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32b04861ec6eb4a540a345081468d3cc3f05f4521ce5291afb3bbdb0fb716dcfe59f1dd524e18d3ffb8d86b9e17dc3015ae4d1847d3d6f5eaf5ccda21c8e4d9486554eb23262ef57;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a7802301d5ad6a98643e0c5d0d8dfa6fb28fba783cd86f6ea6e68deba92a0e53933486413eab453dbfb7d3a7cb0143347d8ad4361f8b14a048576ce1b4d7f192af3bdd1f2876bcd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9eda3379dd1df3a63fd6fafaa8823effeed84a5588d54395df27cf3d0c2f8d103a3190ff81bf2c1d210cf9f11570c429febe68c9e5c04f3044cc95a2ba9a357f159e40203d7ad9ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98a14cea3e4326073a98c96ae3fc0c2a2919678ef7be1df9136b63fddd4c8a4ec7c9d937fe3c405ceb5d8d6d14ead00c2967ac55a890b1471bff0d13c7eae07d7dc9bccb06b8b17d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b30e898ce0381a566ab2ce5c6753c860afa4367e6eb8d9f033cc6014ffd1a213ae287090eb8e2eeba6ba0658e5fb20f31393d7c4edecbf05e97f4cebf84b295d7be511e6147e4ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85f0e4f876e1959545089f388ce97212d1cc4ca9b18d1444d9cfe2af723183c10bfcdc6033f67a3f824c3e8d8daa75ee4a0916930848d8aba220d1d73128245f809434ada753dcaf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9883efdbd32f1258218eb3634a421819ba183ae95b4415fee819a7e5b7a25e438c96e55f611df8a7b3264565d84a72d7419da4d7d652a2188c3255e608c9ba4bde882e3aadd98a01;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddd86f9e5c7092fa28053b7e098754e6b47ad385084c6d9fd70d2a05bb29ccedbb0560ed5defb9d6be45ada18cfadb286a64b7d7b241070cb0ac99afc09648c5fa83b2a5b41dcaf1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc162532d49c9658c58a580ddcb710a21151c213f2c1f5bba314d03747d13bc46af7dae6135ef51ba0cae2d63c30cd7b9cac7a795567fe3bb0dbf7506dc3bc0126985ff865c438310;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72c93e3e1402c0f3ca81c4719fa4607370d36ff63fe0bba6a949afaa9e0f00b2ff597a02772ef25054c536ce38501f9f703b797907afdcdfb36b11a58e9dd2a831c39093d26bf72c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a3ad41b9854d29fea6b983e13a75fa1c49681cc2f1eccb289abf5679380b58a5f82d56f76766a0230bdbdc9b759fb5c1e8c481b34fc1a2a4492b18c6aedb4df9d62e06a7ce597d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hced3d5256d09b0ac0c327ed4bb46d25feb7934d00869350e0ebd450132dbdfe8585c9dae3ccfbea35735dd88577a279c299aff99539254c3f54062dd1a544a35947278c9c232c618;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddeb2eb3e333d96402cdfcb146985a4d01b16bc966523614f6ae169c64ee60b6a23305cc976b3fe3a7ae33df49ca3af7017763007799d82860e3c6cfc64a1773b4ab4fb851f852a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h676b77bec32289849c4cc3de2d41ee35ed7658feccc611644a5690e648ff0cff9e967f5fee96ea361bf82cdeaf2008d9326496e1a62a984f420e21a3932b6926a5c1699645069dcb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69cac59ea4d3841c67af64355564c71cd19d9c4ab68bb1bb92aa78170257dcc4942b109fc2fe87a89d44b1871c6099c9481b8b992df299b534c682e985cf9b3b0865198d988a70ff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h893823dd253720db467521000517837ecb6931b65939690093b19f4b6f765ac248614e825eed60f84594f7cc5ef1a1ca9459487ce8ebaacc4fa7f848fbdce27ba9916cd36960677d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17a7d55ad0662ba66084c401508544b0ea2d40bab2ca34dc3ab045f6deb5ef3ff822535bf24768961015370692a7ff9cc1ed1ffad380ffde8e106d0c10226f13a5013f3c947d7f3d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5db69db5a38f825bcf337a4e0b203e09ad9bd9ac1619dd0a3eb97970846c14317d44d854e809e1a238800742af56c992ed43472d671d03932b5e54f41748fbb92223f7249b7f5678;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30696022336c468e8282bb4226ba9f8eabbcbf496708531b5a1ccab5440fd9a1e80b1e1060c8026ddf6a813f73544efee5371c3eea0a3acaf3a9eaefe20f85d12e6bd7cdd7050c9a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d2bfe7dd7ae1a529026a944059928d56395c962424980a0e4fe2bd20d596a36c748302706be81e9749c755e0e6f2babcac9c6ec8208b2fcff93a7a20c2553da5e48dedb1c5f7d9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h47427bcb687509562d0c24c80ea14f064c737f17b683247622b93f9448cc769a5b0839cb8257be71a5cd3103d2603725dc47c05d15afe0757bafad0349917356d82e34f0af8f858a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bd50c6bc4ccd327431e170494e0a3a0dbb00cc08f560f8356f62405c5cf7caee6ce874eae422a1ebc474b3ce8921d647921c66c96ad2fbe794e4a19ca151cbaa347980be603e925;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf309b11de8dfbec1fed2f03076db3d2c4f52740f347d4786e6e5c24557c490305f8540f8e6e6a656cca48c4068ffe898384d9294cc30c76b2b92147b19b343612682fe424a35e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1ff29a8c2ae503eab5e549dab9584a5bc17919741f8e1f1d0500e2e704adc767ec668bda7a46fa1df057f0186dd2e8e72bb66cb8e1e78ee3b3d141d577840cadd08d713905cba0e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3e1563b66f1ae389fd6071b151a05ea2a7be75a8166844cefdf5bc74bfc6ff5a4820aec0488255d21099b28edc9f2ce386b3e00761a68a536a60691a1efe2ce18b709ec781abb76;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9dcca8cbd7ec17dca4622c11c0d96689c720583f8d2cc1c11090cf976c8a46407c3563c3a50f2cecf4320cc32555ebd25ea1b19629e847256793d8e10d45d1a0aa86a0c514a94d32;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91a76b82921f174272f3ee3615817e12f8020b3111b39ea45e031f375d5a21bc0d00caf86c6f03ce733ba5b3ee1790fdf2ea23f3754ec46efd4e7eb79aa9f5ea2d1f0724b6c6191f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2712eb090155bcc70b279ef991cacc2a158c41b4015c8696550e961f3f5dc6f239a6fec7e5dbfa037f966c54f4c08eac1ace51b76fb7e27d2d4c67ff0a09b618ac8a2911d63900d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca0eba1c822283c7870e494c7de3ace237a160310955aa2a20e3e26a316e70ee4fc40b6031eb0ba9bd892d49f8f8675b39404eb6e286cb8eb08dae081ec7079f13357cf9942bbe02;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21d4a4b25f46b207fac464ee974f735a008f14bc4484d6d21b04b324237d94c6e4aa11b9a9ac49700f9b2d2e61d6a66bb0d01c4c82ba7579d7335ed3ac1df8f19344d51206c0176a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c20fc0de7cc10827f97336b65b5824c9f6dcd92d4737ac5d4788cd6acb02982d260f903989e6a456da01c7a0a7b0f11881472b83c85be2566c439cc38b7070db90e9562a5a83cc0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc04304c3ee64c7642e9519b02f751c5deee03ab0157d7fde0d5322215c5eddc87bf5a7e5ea9f5f458dc58ee6432a2161da3ddb7d33b0ab3f00087ee418f644091726530d9c14932c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee1d663f7d9d34a5861746653987515bff05f73bafdfd2426b6ccf17ca2bfa9eb61f5fe39f4d3f6563d7c2de3f83cad5320f0f1ed5e1ae1e481d9bd4492bcf452d92d0426bbe9857;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ff022f08bf0388c4171092a99ee41875f3b2803cd594771fdb7e8210a348822d11d130fcff2c12bf8fd8cad813dcb967bf022fe50821b8a1c21c623d8ad94202edaf9b017380db5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82993151952784e2178ec7a8ded623f622eca588de5b2a1208c0d14afb2faf416ceb30321b444349e9e17bdb7e999e907602f696627f75dadb66625d536abd0596561e872b4ce3dc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h846e27c6290c75f7df1c1eaff1e37288b9f25f28c1078a7ba6ff9c1b48b858f74598b5078343dae20a986f640697422b2b2c8f17224a370212160344dfe81423396426c28a2c2ab5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb15b4f9b81122515de49b24be2844f02f773741191d8d92b4955ae09f75d991f785180268da3d7e08ed45071230026a3aa2a3430bea0eb4596d7dc05172b1b56c3d7929c4c09e80;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h824e5fec0b7b49024a07ef8b9a5417391395c2f0194c061eab24d46f47b8c3922ac6311fee2f06f57b75b0598ee6b81fb873189cf3b34a01a9e75faef1bb9a61bf57dfe54220d8fc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f16151cd32785b3893368eeb83ec35d83a034732e6991d0e12cc85edc398fbb31e63963eb75039e6be5bc9d2825c87196c8135f386e6fc0affa7655ca82c1a7f493d434df2592b5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd495ffc330d06eb79ce8dc5621a77d52b6457234d107276d8708ec57154b334d3cd44e1732d63045e48ea25c2b69e29549ed68307b3b6d4832652da5d4468cbb0eb275634b241ee7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb23ff1ab1f12763ab980d70cffb4ac6d1e455dcfd61b0b6956cb01de55ee5ca8295536beeed4ee383b19b1ce39f8bd6264c33b18503c712a6c42e9c78d6c58189c5c0d90cbc3f67;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b10f586f824a04b3740b4b4b101b1345d1107b5cd31b7c2a34d755ce5bf5c817b5e2b202d2dd1f8e78bb1151270aae510ea53013e63ce2e4a2a4cbf24341f262ebaf0a3e3d43a3f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h427cac881e5283b106d6ce67834be13af68ecca2d0c5714b6f88d837b96fa840ad9fdbc8dc544016717c7997c4c1bbfce1d8e50abc44617b0cb71ac63b86550ea614dc8827c3dece;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7777b9a1445186e8088bc393e8e4ed7cf61652da949adc5901be1f9b21eb4b07cac378534968a9fe0cd4a7fa693d1966d8d8119a4688fdf17551179b3bfbd70f7fd36ce31e3758ec;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha514f1f2654bad7ac0b5b280717c7b0deb512913b50f010b0dc8fbfc2eaa886964411dd783af917d78fcdb2c98ed2327115c49c830aef1d135962599de964fc42cb726b536b7629b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76c75e214307da3a1c87615e2ee711c39c41de9ce4a647811088fcf41dca7f5cf39e41ff752d8dc607c0ada190347f25d29c5ba331a1c70e55d750845772a98574bca61cbe97e9d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93567a1f3183867ccce3c9e9c7be883150f174beadba76bac6ad26cc1c8dc7df50caa62d896479c051a165b2be5b4bd99df5fee568b19f7a598058894e91ce4a8b58720213a8c116;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c088f8b4036aa1080341d000722c68b873c4fc59b2bb80e07a0d95116975642493a00674d25b695d0240382b76e57f5fbe95d8f811994f5bc9883a3b48ae41b302a26b1df07eecb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fc88cc1a0a37ff6e8cd4d1c209e5678f638091276ab97995c214c4701d1eb083fd7777ae63d82ce8684c978d6fb54cee915d0664982cf49fb01aa1938d6086e28987006318a1258;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36e0f5bc54aa0fe5b6a363a43594f4ebc4dbff5ba6866ae1e283353643e78b6b349e02041dd65adf1e3846eb0cbb7f87819d8ef0edda41f93ff6fc8985d76578a082a0650731820;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a8fcb321c1b12f6f83ebf12226f11e59bed0217d2f3c38f26340c59e0dcfa4d32689bee8d1d1e9087f480e31f33234cf30574cc3db93e5f6f5044e996229245dcc39409a749c130;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97346b636ab9f7220bdc9660d5ad1aa4e45926241f24d9505749cc9a0d0005ccb7f384570a87670cd899f741a5ba1ef9d2c57596af9ae712444180549962dacae29c6b494f6682c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he27b8b0c80870f8195429c1fa886df911093991cca9954e046b00262c3e92584872a72552a2576d2ded33f27147909a2ce98edefa342336a6fa480a1e63cb8586bc2fe0c6c94cf84;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7049746306504dc65d8d7ebad0c8f774eb7db641b12f384eb242adc3fd17b3cf33dcb6815b971507a047a9e030bdd0cb897ed9e973f2c7da4c255181b12c8b4b7ff54fc21945e61;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9da251686f85bb8c16f88691002e4bde63e6339d158eb704fcf33699c0b6e0153ef77061205c5058992d9a83eb191da4060fb8bd6275dfe920d2e85e2144d360976599fe6c57e62f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cf2232c7220edb944dffafdc2ba902e370e2c13c28cbfafa44f894268a06829ac2e2b550ed3dba010991fe32e788682736e3c7e566749d792204ef02ec45b91918f96ab106b0461;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf44d07d01f6c8b6c53ca61b313dba664cc6906b90f3dd249e54a4a69a462c27c9f529baf1b16583351535e492e0a71a59a85a9964a5c0972489b8a2fd23993f29da6e7a2e9347841;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2eeefaeb28639c41cd1145fd17a21bcaaab7e0354e4a40b87a87d300f915f1c822ed3a4f2ef98a005f05fadb3b9f421cf683eedfa81fe19eb407b170f4bee9d23abd19644fad7955;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a9dad6e716f20143b56d28bd3279e0047708f9efc79db78875e026ab946b4ef2400e6995b284a18f74ccf3bffb87bd2ec6ad8dc2a6d7090a4596cdecd58ab5f6f56edfbf1a1699b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61fe3510b77df5bf674f0eebe99edb8427ddd66c759619fb74b99ca917290e8d4f96a69c0d79d683530ee2db779e72e473d6f8c580d91e9c041dc37e5146153cf91d5684b614a040;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h883fa77477ff53f5e78ff379a0fbcca138cbefd1783bd01f34a30e9e815df40c8894dafa95065b4ae5b065a00ee6718419d6dda8bc68507a9eb6c1f415d6e00d70a140c9881762d0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7346f217cb27bb050a59ea1fc80160ae8be52800f21218e53edbe15eb158c0e498dfcc34aed94dfcdc3b047275fabb227a2bbc5fb7c20b488fec67b51e4b788fe6e588f55b0fc46a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f8e1045a842f144713376bbd3687568039f5b00947cc0443edd7bf399e6e104f513f80b92a6babe0ae40c3ad06b7da983bcbe12c90f5f1894b3ac5bf59257c601d6924c0862b824;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4dc1bc4fe990d84fc84cd3d820f607475528c33580ec7951a98aef9d4bb93ea58ee86096c0a3c32b02c7d3f8cd83506d52a3178675fdd2ca45f097666369e65f257e715d5b8a9565;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4b96e596a461ba861a29659306d1c9eb8c7c7109714d58110aed4e474c596df562c65cf686305d40466253c99ccaaf1291910339cf3b630f263a14d6995dbfc83a1368d00008c6c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45c79e9c95fe88d89d5994855473648088c635b139896ff03ab412e54206f0ad293ec724d31579ffbd96de999162d4c61fd82fc5e836532642eaea3816c53e6ef236fbe0a6966b9f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9fc9dbcaad24b31d37cce3b078be0c17e90ee97ef5222ddd9ec3fb0a50e87ec27817675a25ae504f7ffdf944a933dd1a25c5063d484eb292fe56861addf84cd76c8a409ef40557c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3be194337cd4a0aa10e1c4489ed01060ead76ec46f18b0c9070467d46d4e016a7276d2c0ce5e54b0312c57dcb9c96fe35abd084d29fc7586206cd4dc8a5ee5b81126cfb20887b63;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h90ecbc55a5c11bf4be8383dd14917614aa28141f8709bd158fa5e003187f39aec5670b27f9dcbb3f563d15500be12b65b1ee5d74fc9136c38b73d76d63020f9802bd70cf1412077;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba59267fccd1851f0709ca1ceb3aeb2dfb706c0fb4b00eb7889a6bfe6d1733be91a22f83b51cee1ec47cb67497f244b3a929264ba6546975581fda3a86dc6d843a029679e5ae307f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf8a240bf413b62a66e135afb2a1b266bd654bc7f7ccd8ff24bdea7c6ffa37650a6f21252c59409bfab631886c1245fb4e057f5f6dcc93a8796400c793e64770661af8d6a6af30b7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13ca73b405c415d74ca63870a320ac09853d080674f816b89ca6dd89b94498069d9826c1f5c1b447abf39e59e4548ae6e28a5c6257bc7720d261b4ac5cb56b67dced661bcc53b279;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6093db1b92023308c96f0ececd2b9a6b915c7ff62fcde8a36b57bc419f2bd55ce01338618e3ff83d3304a6bdb58292635f86b63f0c9352b084cb8127534826cec4aba79b52253985;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcdb144a8e850b8125c554f5972342859ae7c71d8a883025de0ec600f0a1c5b3211c5732b5570204da689632c619f2a9a917ba3d4cfdb251e4bfa136af4dede1482206cd818e9d64f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cfeb4395be174f9a98d63a66d1f96b98ededd34bfd2d6fbac84096b1310644b109bc16ec1b0c4687556ba66acc1fce41d7f35d0b0e6e918ac6ba346a5e234466ec2eff43fa3006b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53ec89a5e3af984d481840d27086085aac1ece3eb2320314ace99e312127b4948bf967b20d765353e12da8514f2705b89c62a794082af7d0cb54c1b94ac0e0d5407dd40c012365e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h929f6c9a5f62c5cf0745514035e7a17c297fccd19a580af4ee0a3cea28778c314853e4a54d0078723f76064ad610322ed4f01960c575596f592de648645a4f151763c856b770121d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heff0471c89af69acdec823173d9e7aae3910523a131ebd31145c27da6ea33f96dbf38ef957df341c56d11e66b26c5c907f683be6e173dcfa1e1aecdcdfb7ca26d6fb13cb004d69f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h974f16ec89d31ba0ed44fdf4b7f6959dbceea35042fe7fc4cb3461110814d20c7c751d48a88eb34d4ed3109580d0ff0ac4037fbf48ce0898a56079335667d1f6d6396c509f7afedd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2871e1e0035a17ca86bc6dca190038d6a9be112b0bfa731728204f01f90f7b55aeaf31ed273d91e3a6190938fb640d5da7144b384c00b50f6fc3779553fdec7f4f3dd69c70a67ead;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecb089138b856c4e91ce2b20f27b274dababa035d9916c2c3af8668a2936651f28ababb5ef3f470a822c80aa00852ccca8a9d23d070be44dcbf93e2aecbd59895e74de906d2d5542;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he36e1971d5c9074d107bf2ae85904f8ff44bdf1993724f47731e85fe020112dd567eec018297429324bb38339780382bca6f6d3f4ed9bf1cce56fd6f30ac3746824b2ae16d0e3868;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28cd62c96e7be9a0cc06938ca442aaba1284b005edf88248b07aa0111600710204079978c530d2174ac94b15b03b2511fc448db116189e1976993bb4b8471e104a02f4399aa23895;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a0c4b7fe8882ede568e0a9889d1b7f2f08c819920b2fd959179064b7aa1a5baa92b8a2349f71291614c278904448d2591787d56f11a792555a1659b1c656402b2f5c3a507870460;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6c34f8016e8fc2f2160d75cadc4db045d0b7a695ce552581ae5c9deddfc54928b8405c1d936668ca6cd89ff2d1e084105b66a585a43c6770136b38dbec92f3a5fa751ce2114ec91;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a78e32bbe689d12a2ddd1c8e543f1044d6d7c790fcb61e81d42103beb238126f9d8ecafc5efcdf2ba98e6aa190a347154a6daf2470397bb13c0cc2d2da280fbf3984789309d99d9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50c16a9ae42e5ad1f34eb2180fdc752af25aebd64684c9cdf0fb1973529f7d12be623644a7be7c7070298a3f0786530f832f12798b43d87d96ebde0245caf9a5bcd3d3bcc5322690;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf85d2bd2a4ea3233d7973cbfc3a639cebc8377c73b6e92d8ed73a27b381f01bd9f84c502af55efd2d297d0fb9aa1e068000cb7a073f626478d02fbfb01bcd6435874081fc97f1b64;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f01ccb342549e922253b27fd73b3dccb3d366ee06ea559501489bbf2353d68b447e8ef21a09d1447fa9ffe13a62d1167a034d14327a6ca16149f18da1e1704e37b09cec087e6d36;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4931df78d910517941ecda96550a955eae4cef8f1045fe090921d385372c405ae5515ac53b2fe0b87670b4bb487da50d2a75e9f9e0f806ca4657f243f0fd9b89a9e63265e31f13dd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6165780bbff43dabd727d1383a8e2937eeecdbef7c816c202fe3c62af8a0bed9f72a34325ef9709fee50851cca88f33443041bb35e6a3eb53041ffa2a4427bfbc0dcf6ee73138a33;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0b517312cdd91d3920e32b03c17e1b5881f77ac92f49896b7834a62f3488798550798c00b85d4a9ad23d24a93de324be37e8dec91b5b5a99502b4b7894077c5d875fbd62b8c23a0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13cadaef554ff2c1805225cb04460524c3b04acc7c26ae97e2c7fa297b851bd6759bb72107999071ad285d08dfc34aa1010064f11ad02f3e0919089bf2e299586035aa4469bccb34;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ebc14a93bd5a913458fbb98701fa2414e421e8eac9dd5450fa9411b90128810709ed848b24d3644d3e5c9d5ba69d7112eff8b282e47bf48445ca83539ad585c916be207cc4b42ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6958c0b5f19b8405cb07ab8fb83342de6eee01141491ff423f940306bf9c039d804bd9b99dc110862382a5bf7b6789a9a8eb662d76bdfd4391021a1aea30837ecce7335f0a7a87a3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e37f1f731c1bcaa3915cab35ad9eed19a2a7cd9fc9ec51d11661bb1eb87402cded13f33946332603dda8ca5ef0f3833d8af7fa29052a62837a62c2148c2dcd82518a8ea5f0d953a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h563370a5eeecaec63ac6cf166dca6fbcca9fd922d946e5f3b61d31870d12904cbfd541503e663f240a004b9edbca605795b711d72744075a75175cc4f9e1c5cfa0a015f15d1635c7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb436cd8e5d5b9bc55ccd1272ff76f51d8bc22bb2011888913c448c4871f6efbbb152a302bd37426da5a29caf0e75b5e5c857a7568b346df959ac6994a4b874e48c8287b8c30a9047;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8127610f951cb6dbdf37c5c4213806b099db024354ff68af20a2d7ccce5b74591918a0ffb7b74793cb5e9859f05fd86e1ab96f38f5ce0cf0135b8405d21fbc0cb1c64c0f8663843;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92332cff471b3c8837db08d8d0422b048241fce8c288c049a40a3e8128c86ae186c60c5eded5e07747768c263edaa74f25b97e939cbd6e8bc5e636ef7840ac243f81db3dd3a6037e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ff22d757dc29fe580b31c3f83e2bd29050913912c9e8404d9f85d92a5bc0849f568fc1680a222e3eb08fb34c4659bacee0f37b71c2237a133841bec408027cac9a64fc18b530f3b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50d38c610c6677fd4242fb33d2b18e28ba2bdf8e75441dc7183c1718cc4ee30eb43c67f945645a7180f9460607f726ddec15f44edfb5e6c33a2efd88a73e6226213e60c6254268c2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f42266364e8ddcd12f8db43d3cec2e29ae1c8b2c4b2ec05a0f6237b5f55caa37a50fb273cc66d31d1d1aa2de08db136829df660008883dde312ca04c6b37afb5f8afbd89dc5b3f2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfaf999863116213e1f8c46a71b05df9da85b5888def57f3487205e3f7921755f5d504cd5e53195173f3ef7c0ea4be9eb6cecbc8a16845ab86edc81b351a7bbf507a77e2c4b41a929;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb73faf5a569475dc7758a42572e1c5d248ea73f0f49bf7658e36b9d770b74e5e2c98a97ec925702caeac60a29148c1e0fd16892989b0833ebcb43a0e5d9d0ea57c9b10778e15709a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9899fd39695190f7a6282b924de87efc7981da3711317edf88a15e88371459dca5ca4b28b1289fb0eae5c83741c6c188b1f42b9c63641c6b2169316e5fe3aebb6baa2cf8eee2a402;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h184d05e0a51e67d6afb61a391a2f4d83aed800c6ebb8e0a0a6ecfbfae07d0295d94f1b8e2fedf0e186b5b18db5d249ac6fbbe08cd37829ff4f45b97ea56ce87ed5458b72b91fc1ab;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h814cf3a3a92016ffd9e2faf688d31dd55ae86706c8680c5b8a9453b0ceef40a181bd6e137c37492c491ab5150eba12038750f6f1656257f8005c1f4c5455b42bdc0bb6cae6ac2ddc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ac00e90c26e54c071ee2b15fb406181e6f9ef38bec97124619adecaa1f7522f01691a355b6aba872861d375ad32a8da5b76146ec4bcacfbe099d74c22b572885235064dfafbba3a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hceadebdc2535266e11c1c8e56fde11a2a5036f03a0d0ca1eec3f99eba95b698af2446439a36a3d67a3eab605e61cca4ff28ac583eb45268fdc1549a2eb4161b29b73e3923cdbe391;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a1a5f1c4e6435798da77ae9d6d75a9e3086f1e7eeb97a03b38a93ee7cdf1b20d4d31ef54bcff96fef3bce6d09d83fdceb8b2498b75bf056cc562f4d5d3f6fe39e27bac2d49433fd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24291abd1dc234ae05e21b63e0159faf00d055d77648262e1d9acdffc5046b2e02289496eb12c4f1cab19867ad51158d2c905214a1e1c811ac1b6b52a61c68cc2d1c8f7667b452a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d3b2e4319d1dbd20f831bfc3d52440e46f9781c6330b363c4c8802c704012e81de1523d96b52cf2212cca398a8ad44375079c688b73149512f896be35093c1d9c5770aa452c92df;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b92a978391bf88b0cbac69fda6d7cb5f6323c103558289c20d7f39fc9939549d836175aab5007093593a087f7d60a85b7ee0cc5c2999ed50e327fb2b4d17dc2b70243d8086bf998;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd672e0d496c92127b5396509a9c047319a233b8f56ea1364c04fb8601507f9c80f3f03f7869ec71f9136a25ba5dfd39ae680fa722f6227e0c37c3f4ecae019f90430022e60b891ef;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h311107238e98df7bf5202dd2fff44d7164b3772e3d5cb2fbaf46c5461a24057f5f5411f7747e996e158a5e4e067d9bc87b6095f587f5760cb9b53d515aa460e573a0db88cc487df4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha131adc73c634df49224b1021e0d23ec814b51de5395a9c58d3362b13323f53c5f1b05a67a137215ada0b96f79d6b546a324416d7727998ad1777d81db7500a67bc5e6f76765187;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f614a066841f6259120c471fadd392c268c763d8035bbb2073b14ffb18bf9bb23ce9ecdc93b0ed371da62c683e6c5e58f70c4ac5e7efa833588933c525dfe36c9545ac77a027d8f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4db685c4efb849e933a6939275702bf6df3e34c6079bb13df7bc5dd3fbf0ce6b32987c6a645ce8d6ffcceff01243006cebe2a86ff0d8a6fe8c925bb2577cbdf1631419352d77e0b3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he129255576466e4dbb54ede724c0391004866cd2599ba5d7e8a2d3dc15d6cd389a558310f4f19cf806bd9523c751ce5f68858918afe9f32e8e154596bee2dd03196e748ed8ea754;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf16ea2869aadaffa55c47f9a9d32b87b794e7add4df232ba93aae738dd12a418bc20dfe125ec86488557b275aa111c502d9f5978811d66adac22350b637c8df426d6499bb0a8ae62;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfd8f45eca1826c8175ed554c10be4fd1cb21ed27ed34af43030091b13e686b932cdb3c972ceadc12a5e01cec250b7cde3f7bdbebf44c72c0285ff875586435eb582f16a56789886;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7fcb0b4435544ac5bb0283cef455d0d98a2e8734380f8e4646bb8e46087e61e7f302efb7426b76cb539d289ddfcf6988d9b35f6b420dca15c08f01e423a976a2700fc57261aed875;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83abeb1fd5ec16c8f0689588549c78032ea74dc97ed72cb6a710d3f71ed13e42aba15f95e0b7623b6186e1dcc4934c71f40d95732b1a9f5a82d64bc4550958ddf808bdd892d5c4d2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a34ae622cb2ad1aa591dc57bdd76f7042125dca1bd91315f0ead627cd194a90fa437786dd86055b9343af3fb605837ada74be013f960a78dc0287db290101e275b03d1cf7181e98;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16985968ab39d9203cc5a8cdea2de7eb41aca4ebdd608c8254861a3829ee61f0b6a133ac08cdf904c4d24e070319256e162955f427792e3d8d3b1e9539117de15e82513c5ac4b3d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbad891d6da6a1c5cd933fcb6809c7e9b88644ef66faa5e0f06a41478598b416da4b3b9093bf2e790c9fc362d8f3b565ffb55adc71b3e2aa4ef54e93116bf873509efadee52d492d8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f2d09a47902941265aef0c076d04a95687f8d9b534b6ea21928eb27725c5f16c5b4567fecba067121a77bbe703b7d9303dcf98a96850c59cbe7feb0e336e6fda4a11c41de06a69b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he83e2e0fdd3cd80a14942415415dd24e090b2eb882e80570f57b09db66129fac943f4d2f7993726e73c3e7f7263a7fc4b4f4b70f8933a227ff3ab361cde58a280fdb7c6bd52b563;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1501ccb272cbeb50ff88a202506af553b772bb40aa56fb99aa6d96a9d26d766e0510e81b9ccb2986f4e8a0a8a347cfb4b58aa23d2fad949b6570a1896d7edd856951eceecb0e37f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23f8b944bb7507fbc0e61115b37feea2d1594c6f832c55e7db7119a00db80448b53d437405826f5daf19b002fbb59414d2d88e6a70b90cb14ca992b51eaf26772ecbff5da8eb66de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9ed3c0f8ad806768384571bb863411fa305ad8542b087f4aeb6241490dcebdc304f0ffd212cdee984259e06a8dda0c11c65e02796222e4666745b0b01491301a9217e10e6df996c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc22eeaba3fb0128501a8dba5cbd4eb8e670428c8acc511560fb6293925c8a54ba79fce2cf9859268723897511e2486217481ae45559b61b05200c147f409c99939d9da884a90734;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff66538e0498ac4a4d4d59aedd178de7852ca0224453a4a731014a116cb10785ba289d21a53c8bd960414b33342b3e0c194f70852f794ceb8a377ad3483d2cee5104ac5fa42a75c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f713513cb17645acb93dc66c1e3a37f86ad309b56738d2a72de661918e249b94c41230c3806356ab93b85597a0859250ebfac21800f8d5237bcc42ceca5b691da8be30558468eb4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb9453ce12f417722707157edd1f7bd5d1077b0777516182eec0a8bb04de49b9a6c157f97e821596aec79415c1293787c37008cf69a37895efd9f4656f3b95cba90a681b5b4cc783;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedbcd1b26603c21b808d7000d10732d0859d9a3480282c39edcebf8c3f7f8e0eff4966f9e3e280b73f74a749b5c10e629c85576d65357deef0234d7942eb80205913b524d38d0de7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd0f36471629bf6173b7daa69090d812ccd99dd9177fc4d20a0934e7fa4fd0fd7e8a337af6e642f6f0ebfdfebe2510110838e36ad214dc66e7b015d6dc5c7dbe3accee66e4352494;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6495cb134705dab31d5d79ff5af189c4f8311760627b0cfb74ba2af0877e6ff696bf59052a7ce5a0d004c6841d95688122476a605a127ac49e6dbcf0579646326cd546a45a2a39de;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h200d8d54e3313e80d41155eb8c23777decbe39db18080b16ed4d490b0674a4ff181f72dc34fcf790a9c2ad0b12a58f94f09fa466c27eaa6373e1f3e1b5b2a410c7fe3fdd31aea2b4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h431bbc3d7488927d0a6e6086a9e9083054deb89a46daf28aacc2b69c490805060aaa70befb3be84f73548407d82c2c09d0ba45e4e1e11cc345e725ee4f6df85af8abc0a86823a953;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d2badb51c5dd38af19ba62d1d54e4aaf75180c6917d549ce40c554d306048173bf03de2a544e148db42caee47da5ddbd85c310aa60572e16c549fc06716bf137a647838d941a0bb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4b261cb7553bfa80d5126c760844474a7114ac0dcab889412f830594926636f0b6ad050564133dd45528c5cd0fe3c037f337d48c85f2c4f63f38766d03dbaacf0e376a2e7c0429b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee0e26f7bf5187fcd1ca5a7b69a9c57f86fb160f94da28949994ff420206a611aa5286375264ffb3bbdc22c88adcfe8451ec9d1e05d388f847b96c75c97425d44ccd965310fa5800;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36245e952b3b085d27c530d7845249a6de0360b027bb6b275f5c415b2927266b62b6247f35963cde6da321953fb54449edaf0b6ca5013e9bfca1adafdd0b0df7d4a20704deb73848;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff876a33dd2a87e8e8fd9ea6cfd308371040c373a51dc918f9f0d79d3e15b011d594520548d08e4c6de0c02963d559cdeaf93779bee0526c8f6c1e291250c5b5d35e2430cac21a7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e36268f1f239ae88e2d53d7f26ad26be267c9b9efdf2316215aa66fe62ed78a535c3877b54909947b61752b522967930594e3c982261d89c4a3a563f6cde1fceabaa08f49d0720c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c2bbb7e22553c5429c23fdc71589a17b021736632e9af7a9cf29e54a3cf9601376eb72592cf40fed6e5beb5218583aaed9945e871a90603b642a5dea13419f28ef40af05bdbebb1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha83e68cb7fbc67b17fadb3e19b6ca2434b8c3b69a03d56f93d84f7c0fb6fb85c8a8a4b35e0a748052252feb7c84e2e847bd268bfa70d4302c5a7db2a4c876ce1f7f2fe2238e3d4e7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf693cf405e91e9df242a9d16c0961f7759b5c4f3bcc5dff328f49612150e39a68dd3184531562790d6dd9bc66b3301c5a3b157f4769323404546977ec8182de838aab0c53bfec083;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc9cb8d469d3ca8b28d5977910eac7890c40164cb2a8394d426b8cc8b61a9a3b563d3537be03d768c27a399c37a1e511c64ecfc443273ce5bd6d63a115563ead51c71c4bb5c8c070;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf79959cb200c45ae81d98d3e219387445b009d24d4ae2c8f2092ebcf35ed70490c85f8dc7aaa776adb6529b5a13c5150cc9226d952f2d1898e921fd8dc44d1cd707ed66929730004;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c9bb5e121815a9f19723fcf95df2ada7d957948313665a14d1624dbabf06b5e9c4f5c1f87ed720914cb58d45023a8d9626f11e453207c7acb82ff7f161952672adc7dd1f3e78ef6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ab2c44829a8eb4d632e6c0a35e62dfe9b8b27ba1ccb875d496e29face4c56b9e74799ecf52e5dce7bba82b54c0e15ac3e4f28caa5cd7a5db54ee68ec3b0f96c3abd054f5a078837;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7df07cd9989d680b0bc51e189e3aa3d03a025fbf8953ade1f0456755e2ca5b7ba1d2954c9b0f09ccb91da1e09dd39200bc1f9510877046142ebc231e32337ec843bff231ffb3494;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb5fe45a999a9bb6f14c6054b7bbeee4a5880f09af31587694944c5101b87bc73681a75b25d16e8116a8a12ebe897137e86bd9395fef73d61ca106738e9c278edb872adbce1c55e98;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h206c5ba52ef58aeb2c07cb21964271b1cd4a03f40f8ee3123577e9d191dfecb4d6e216cbbf94fd033d33d6169a58d245b4fb0a3d1ebc93b73df09c3897857b06fb32bc0e3fa9fad1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h560dfe33dd1a1be8f83b892780aed12ec005a039f17d5056fe5414cacbddd9ed614f90d6f378d7b8407f871233dd5c5ffbc4f3245fd33fc67306f56bccf87d187dca8e2b31b72045;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ea4cbe82c93f56708bcc0ec089fb86dd76d3f5a4f65de0fa3413dc0ae0b3e9637949279fac49f0c52b939e8b4516fa2d57b59e58c4234b250f6565c296c41e2d3e90f3a5bbc3807;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38cedb95239a836625637a105d656626060ac4d8f43a6b8ca2b956ed130c2c00533cb8cde8ac8eae877ccc941646b90d8f95658ccc9f4edd22cf38b02fc403fe77da8a2267f3e168;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2774f9d63f6041bd995e63b2bdfaf3cd170634dd1fcc7da8838dc0b7da0425848fbae136aa47e0bfe4bad1d38dc83260d5c1ae9aab139b2006ae2101dab622fa964976115f7bdeb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3db9819dfa96d7bc1a74e825af9a58f739719dcfc056d954e060f87c16cdfbada476becac6eb5705db52ef7fdd09b6333e08621489551dcfd00506c77a89f8ab4cb6c1efa15e70a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc82182597847c91c634e6fe10711d7507e27e214e492db0420ad946f521f7e354cac45bd1374b7f369191b6573e319e6e20810c34bb8a2d180bd6a67e9acddb5e557a7738d06f582;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had3a3775e841390e0097bbb2c51a13614e100c94f767ebc0791513408bda270d18fb8a03c2d716a27b02a0379cd9ebc37ea36900e4396b72f3d0c32e87bddd85961d3b9cd1cfd783;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha876fea0a0eaf9ea9ad30c74dcde768dc6f595d93a1c1449b73eff8a687afb2d6b69789f409c233127f6ab3e5f4c2a85df3c2f5d016b618de600e6303960d93f09bab8ba35df55c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h374f91a39d91dc7a1b3e6af44fdc2d209bf27b4a33a342722f80664958dcb7ed200ba16352ada9363dda3c535b02994784def076109dea464e938e777d92e4966c10e74db619ac5a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h770981e831d3149f4f4aa226631c746e27a64de9e695e31eea803bcaf6f83bde521722e6fbb404db18e3822127f32bc564df1885f1527fceca72a6dcc5245e5b8cd8799098f99850;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had18fc02852aefb6d3734524d47842f0274c74a84252da01fbbc6859397d315277484bf53dfa9acbc0ad5a9c29deaab54fff9a52b73524afe1edf505c24fcf378921229de4ddaaaa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b7bbacc04cc1d65d3ebb6bd30d7606dd4713992a068f78aa86fde4f1719a197b76bd0853d6e1bc8e7f8db94ac21af947fd5ec2b92c6f343032a3ea9c29431b8b053282f4dbea2c8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha66b42adfdaabe4ed3f2076feb18b64a88c54ff26e194a177a9b9d97581213ab84a963259b95c7cc02e34aafdeefe89a97d01b234134e9f7009828fd55a6acc6c4630fc486b42e99;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf703ade0bf8d7fe2cca9a9181080df094b650e82a472233109b2722e4ea3b8ef22e48f3ad3443a798d3137bf7e4c5d4d58e046ab45a68fe76e7de79a3fc81893d0cc439e1838c7a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e44ee08391d81fb9f9570d434b66886f33185329e51b5c37cad201010ba716bf540198a4369ff99c99694390c52ffbbf5d7983c6b26035f241df50c80de313f4dd952194ac98daa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28edd03ebf57f25b03e9f4254e691ff6e251dc378fd4ef40dbebb49e2bb3327b739622edf38aa0e1f3821203f28752fcef78a5269f73cfc7e3bf66d2c1cb976f973601a46a4cb36c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7934f3d7a038078102d145ed6ecc23b1a236fd1f9aa91afb885eb8c62859469bc0878a109e2abab5b5dda00bfda9ec8e303a3eed481f88a71933018f80b853d696e70e02284b4af;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha45fbf0ddd9a9d530ada7cf9df2821f8afe18a861a11997f74126c585e8abb510860cc85be4cc1606dcee5d4548625231f401c0d0ff45baa8768bd3442fe9a242422c9cf44a3f595;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbff5b730b9fe9577d69152bd40b9f8f1c02d984883b96c7e9d835dfa03cb380eab04d2b602fe528e698dd2659ab940dffd9c832cc16aefb2728f964a2f2fea04e3836ce00d00fcf5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1ca28537ac0ff88421c4b2d41dd51b8ca2db9745636e9576ddbd5b111e43c53cfff5919ec32ff26be000654e7976d51d23a4ddc08484b2ca72f8b16d264a1d8d1d047febd90dcc3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6887fa920df77ad60511ace25e2ec4409d1f113c2fb9cc14aae2104db0751c0236ba5c536872aac38ad9707081aa518b04d2cba97ab7c4ab0b2f385310c66bc993b4918720bbf40f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e4b2416c11e63590819467b889a4b19af4b5ea2e628ecab06be7d7a8f0b986176fe4f939a4c0dbcf1221d319be241ebb6595f732826869a9ea5e5a78e989db07d58df2d0db7ee85;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77dfcb6fb8999b27ed8ff27444dfb36c4eabe8e793c0aee7d6bdd171fa1f6bb2ca9d298cdff1da4a842af7b7e26f81ba0e13acff614dff5d2af422c1b18393ca341669ffbf0e9822;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4369865c76488ed19fb5d77f2bea2e76decb30bdd1c9917404eea9bfe1b5b9a1dcdfcb65bd6a5fea377a87aa37f1d690624112a7c5168fc69a9e80b9fc4060b7d5e80353e5f70928;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca264a4d11e05e3de246b90e06d2cbc0e082b0f23ff5da686b88c470cf584429ee2c0dab247e91a911f737891f175012c4290350d4eb0d56a015eee0eec12c2e8a3c2d48f728bd90;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3568fb7a2878106263e2d970fd8664cd92f37b891377f70f9e0e35f0b6b328474fcbb32a985f851ab1731c786eb57117415c014281c8e5d5ac3bc64e9fad3acbb0959da4fd069ee;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f522567c4613b336dc147a81be5464d9179738109f38f77f8f92055bf43b84e30256ef5859867b6f395c64cecdb6ca00dbf34b3135d6f2f4a83fb60096ab4435580eabf26d225ad;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd660514a53b689b49808640f0d7b723be22f6b16275126dafc352ed05beb285807742d4ac0480234dc60cfa52e18017066077c41f6be9d993898ef670992a08b08ec31bb721fd584;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc92f4231588a4357ac014987f7a672445b5021de6945036653b810627a82fe2cdce14f53f075824b249ddce5063b02d7b456a75f542a6bf52574408f7992e06d1637be6e850fc26c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h23c15c96bbdf04c74844f77de848c42fc439cb6a2457a6649b46f4ffaa233600c15dc1f64feeb701777ff0e636640b7c033f485a66310a9d2dfb6405ca56f3a3b6d4b3bc3769be41;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc76cfaa16665c893e5d76cfdb8cc89ac90ca9bd8445956728b672b909f5cfe6b4f44b2fa4763c58415308403bf9de5d330dc2c3b343796c210610d9f22c553f8da1dac4b6997461;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24726dc29ad90832519577f974a3edf327c75f640ae487069bd4ca0bb3d10f2725615b1af399889fb9f85c9cc4360df692887115f169377878ebbd3792831b1a4d47f5d1e6c2799b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46e70298e9d29da2dde3fdf95f0dfc574d33183fef68971b49dc2d389b4de1b00ca7eb0100637ca3f8792ab950922c7b3901e001bd0ebae22ed78232c0f4df2adab10ed2bf56e5f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5aa9ffa1ee51974889f5e9839d0a4c7080e94656a9e9e622cf10a4a0fc86ab7209d2580186ad70eaa0d9c07bec9071cad53dc82d66bd979851b1b8caed9543946910e39a8a45ff76;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e0a4803495ef215db35ac8a82d5933288e9bfc708462115dc39b70fe648113c6d01aa120fc8b9fa5547e27ccc064aec48b7908b70c9f67ea634741aa26687839b3c0f3c2a1a38bf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae0439a97e72420b34e86b8b932f763aa461b59bccfeb4554d1642041c60f3d41153025ed2890caca26274948c53197be4f4fdb57619fbba5dba42279e397fc5267bbceda35033b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3d550d98498df402cd7c6d6863c68ae121ce07ea54bab6c9f665306b49ef890362949744c84a4f40072c948356b7f9320436cfb0a4721bd8a054703cc7044e6e9d9a3ee03f65256;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h720b236b1bfe930de0ff513c30da15748f75008228518c6e2e9ebd54362241fa2f91229eb40ec9596651951c3e9663863c1c9e5f73fed7a7eb615fae80c9629b4d98143729093153;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h244d3393bed11d0b0256aff960eb986a64b376b00fb3c16a479487d767347005420da09ef172f09725bad17fe67798ab929a9eaa82703727db3bbcc517c95a62e89b7d886dcd84f3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63fac2f94a197c8fd1d928063ea8578190b5485af1151723af82bfe1f9484aad21ab5d81e22d546db8a975293c4df6411b4cd9789c944793e2cde4d1ce558099b79a0bb6920d912f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63902f4d36395ef6a7fe7af3f4f1b47719a3c7fa6bca8a87f58d3d70ffbb3df903b4ddf8d3959543cd51d0172fab047f76da7e578fb80784cbe848261186fb799e5060662cc422a2;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe3ca99271b0123d16ff8589fe597cea3250432bb64e4fd46e6586ba258b9d9d46cd0304cf9510d6a1ba224895e75b97448756168ff9cb736d3c84765406ac1a3dd78896c6477b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h59ed6bf879ea3f7801e71e453d1e4396197ee8ef0ac5327fea9f84e2a072e41c5a2b4d5a1e8fc499913c5251ad5db099269e423a4ddbb09fdd78933100ecc6e126586b878585e80b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5838795aed1733c81cd981900bd0ec34ff8c35e13618fc01798abbd07ee55716c823e45a9238ec1c2f7a0f7f8eed919eb6621843d204de759c3f5a3c993659ca24706d26a27fe9c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a5baca6782e6efa53e66aff114d8329e24460b1210f0f335c401cc342597dc98760a03cd8d206bd8570747d291bc8cda2ff7e9e627920bee63954d2dc13d6e7bd8993f4232f39c5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58737c37069d46e86f834fabf9fa0546d1ec977d9702bcecf1195bf766c569ca387e6977381d96a97b3d7ee6e37fbb4b2f6e22a9f96389aedb22e6aa9fae2d062fe133dec27e2aed;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0de85fcda43c3959e9711c7bfb91908f1fb6214d27395a4e4617f0ed8ee1af6d12ff02b1bbed3baef9039e5b5644a08221128bc561450e1020bacb8c0615fa406e21d87079e02e1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4da2b3c9ab925107c227201746dd8283aebdce8cfcfc7fd11fec2c6d19b85c5f5c4f3845c4813934b2308fb9b676aca0281efd1e00a072eeb7e297cd4c44b85c29f927fd037bdf7c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42bf684cddf11ec9bed761a15abb9507222df5f913cdd11441e78a5f4798d7ce63582f49fdf4ca7c3347c06b81d4453008e08c2d881d458e2b2522c3382d10ade1aca8a4336da62a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3d2421b883223e2439632762fa2a444af5bad1f15164e910490fe156fccbf20e21ba2e7f5a4feb1f29eb3acb9c26e355f498df0920167fe537fb663ac7e1e7ee647cf59b8b3d842;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44e9dcd51d17f2c1f2946de17c1ad298a445fddff20dbd7c6f0c9ae480f76c87266cec602c7408a584521dc4a50e539acb59e05481c6f5219b370c0d41fe7448012b21438db77686;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91d1fc3cb531d34871be648f5dc09b11e279893708a018c82bcb9185600ea74cbc283d5165e13783a1dfb52a9f849c304532a0f7247af7f1fc159e5db6f9a57d7c58f973e2205dff;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b0b30b14f99ec6f29c82c6ff2d1e36aa087462e779fda28722ca3abc10d0f6234bda2caf6956ddab5ccf6e90288401fa2e6fa3e368374455db67871e5da304588d34f909e42b582;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35cc2ca41ec8be28598f777547283154b21c8aec2af932af5ec9966e7b87721713a0d58ff7c7d82222ee3ea9e47afa95b967ca4cb43309d65d48ee1c9a9c0dec11998f9690a2babc;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8169142d04e720cfa2b99504242227a458661bf5bedfad2f8a00c5e56e66583361150ef99a3dc2b0a86d102575ef2c22c484f4f77eeba9d71a5673c272130e7df669f9d12c9544b9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8fa3bc830ec5ca5cc98e789dfadb626e1c24478af089c63d8ab8816f2ecd47b26c3ac1e3c8901433d236e5ce8e08c4aba5389daa8658e81628a5bcdcd551602ec0fdb40c9654718f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9abc2fe246bfe3105402c5a028a986c1a89619ba98e777bf21710bbdc3aa56ac6859d8bd257f45435d88fab8d1d16ea4a3bd8bdeb6e25227d70dde1cda5d75790999d39678d163c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf4fe86227737a0f790cc7a6d30f3403a19ff3fc03c2c729d370aadba28a105fd3c9dd359c7dbd5fd18d51886578eee8ea99859f0294e719485c8302ee52ac90e39475c9bc9727ba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4548e02c7035556742258b7c8555c82e04eb828e5baccdaa7e02662efd8aeb1918e2fd8cc230a3b4026a554f79e2c81dbf2732d02dd575328f171e4cd11bc55b4955db3350eeebba;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd24d065e1a16cc7d3e63d9991c28f0d2caa0053b7e521bed54ad90224a6fe9f01def60eecbb25eef9b9812766ba02a87a1636525e6c52304f628bd6b51c6ba3fb3f5c47dc09d2db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc17a7cacd7adabc775a86f5bf524fd18600c91fc1ac097622d0a4cb1c14b364d7a413fe352a66d0d4718ae588f574d6798bad7d80031456c7d374eadcfc103c6af8a5fdfd7ae32b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf38ccc55b1952b655a0f5cd2d9189023b19bd1752f49e1d7851bd2ca39ac841e185517232079accf55679dd62f7c8d11b18ffdf57267a568c410510ff2e694847785e90ce3a71a9d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77e12f764d5f208c0c122f18f493e20f3d648f150422237a6e84f2a95ace2dc1f530ba5952f2eb5329ad09473258f5826a415e2d898c4de9e6dfff6017f2242bcd474c80180d1add;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99fbd3cb939cf7cb81d4b5abbefa681856365a0f75263139afaaf88e43d4e5cae89cf7317f15b1a415135b0475940120bc37719fcd1143bb6e5ef20ba78b0030945bfc74ef5ff758;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e39f2ffee56e597f61df0094a3e868febf677067f3c79268c49a1a8d1d07fee0a57fe627d34e6aed5851f07564d37d0077e8721a2ea468876cb227e300c43c762f84444d6532445;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91669b6b54dac1c55e16acda404210313278b28c9166765e45292893c72228fb32cc97ef356266774e84de95f6952cc49dc330d05c9336e5376862ff4575ee0dbb293aacad49e1d5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8448b7fc98988a6ca5fafa5bf4090df2b7291caf1858d5e6763d6372428c4296d3b8c85d5a112e21d9999df5692fa46374c4faf6b3b7fd2a4f5d5601acffeba77ce54d1f830eb45;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h862d06bc8e0db72fc6cc4d73787dc474c20a4a1bc17783e03481e3747d489c1bc9787e2f2a93009f856e7799875ea3e2965deaf2d231bd26d4bf1aca1e49dcaa075baf2a5fb3544e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h77e1c39c43bdf0843c3afe1b817a753eb18f632a66c974fa5138c337aafa2330fd27ba87c1cdda6714834f2150819cf7f97e03715ce920e7b9a88b20d9a504f280ecd6a67e3d13fa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99997e56f1c5e9a71bbfd5065a8c335fd14e1ab4501e23f296f50154436aa9aabbde8bc7d18c86301f37fa84fef613a42e1ef24624904eac0bffae0509310bf52efa9168e8ce017e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7d63da5eacd0dd644c687147e7a90fab3ce495df25d3f4fd53c65565294ef674b77ed5274319db6c067725be8e8c4f1acfa6d5c3a8955e492109d5ea328bfa3516f38e99ed2784cf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffd94243e166f8c1dd1a851c22efc7992e14c3097b63c6aaff76658a63e25aeccd42b4fe39cf737d4f146256896df804319a34ffd477687c26f1298b266121fa36b2fca178095ca6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha83ecf9a7601a6222a63984075e594ba4e739fd94c27edd7f0868ba34cdefb2ebd5a2ac9056f0103d141ca2fb0bfc187cd5a44486989c67139110b7e5d164ab22453c3ee994a3383;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4d8755de92de586e2ea0dd6fe2d1d3e5f09f8a1583d2389d20d338a1fda3f4b94656bedb9295dc6a887f30e8b424a7c764e7abedd19e4b8405ed56a531db7e6224bffba5f9fafc10;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8cf98d54d0571ccfe8c2a57b6d867d30da0630e62e8123cc50dcf8f1aec1281c350ecea76af10ed58a30f972cc4c2ff8c5f7affad67f308d53a085aa224766bae1b2b81e8d7149ce;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d6b8cbafe5b3dddb0b2ba850bddfdd7daeff08cc53b82d4c451896ece9d2f074dae4396228aedba94fbbbc39bc1816747edb8d1499af1d06d82c5ef9159ab8ccc8e2f78bcc5ffbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5a69fcd727125246a767ca9de1ac2c01bff0fd07de31f4c3b7c3dd51153c1a3b498564aa2aa99a92adc8f2bee9c3ca617ca6d7702e7188ebf5c634486efd0a1a0468858c22303bb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6141365f894e694249605dd59afa4ab9b5524bc19bb5d2e0e1ade2581d98b6f6676570167bbc305b2272044ec08b6a497067620405d8894ed081a254a2fdab6101515d3287a80c5b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c788639859030d1325dccfd251a5659a3829216041610a003dc26e5cf9e3ead947eeac086de7fcb5aa355357e8c492adcff711a34b5cff339ebfb4fa50decd138a95b547a3b165c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9eef839b6afad37bcc141857d5dc437c3bad30baa20cd6c61d7cb4406b7c360a02bbcc05d61f4c0a64f444141f8cc103458ac6e6c013a2e25fa55c1a117042c6d0031875b624421b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e9a5d41f92aaf3c5aff65d326896042097cf6b68583c850bd5a5cdd97472eb1c5d958bbe574e175b82b4ac7c66aafcf12a7b7e668fe866255d3bcc9cdcef37259d55583082df5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he95718bd7e16b1b2bce0988dc976dcba1d0fd9d5e0d226375c90f90f1e776c0ed6c5b272b3d3e2a91a1ef3239399be216e7ef4f7dc5d8fa762a0d52c65bbb1a678cd0a4f0e1ed4b0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa4fec2f8f62ac92c17527c53775af3b3fb51738162ec6a17efdc93fcc2a7ad83d32b33b83b3418b9cf42bd51307416beb4cc63ac6a72ecb03963d156f30d2aaa2c7d76ecf0b3c59;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27717ce0d1723905caa835b2b881e4a9de6240894e589b4a17fe43b9c003210e092d83e2af6fcd4e985aff24de4aa4efcc21926521989d448e5f589f8e2dfe462028c5e6511a3c72;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f083cd02f0139e4997e43ef235bf67121f0f34aabdc7197c6d275152e69c92f438ecfe16e1a6a14413368fddf30e829ae05c9d16dde81f241f1ddb624f05751e78e10937f28db66;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d9e66c8c66d3a2ce5e8a06f2902b48ca05afc4bef8bc5c73f3157ce8a35ec5ddf33c7b54b43a8a822b08845c1d17989af4ca1888cbb304e92f4034dc205312708893096a416c818;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f70feab8c1205e65394f41578ccca19cb398382f06d57e6d96b85dcbca0317d5c1949417b20363c2726064a701e92e1c3f6b1194d2cac0a530d851a89a6a0c45fbaf12a300e047a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd220521e25453a469fd4faba4708eacec57dbe34e8de4d4ac384384b4cce6ffebf0ec614107ac4437118ff1fe3e929a7e9449567b3659d5c94aaa6fda18c53fb4278908501842cbe;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h703274d6107461833b5a8a73a2e963c88f618e824d84c1508b74ab3907c96ee9d209d6709e4266c6da8524db28f43b1e1dab3b1de42899e4ca83a6e690421947cb1f6a6949481ef5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6782aee1a7842d24827b75fd391524654f7d1dd90251f9cc7a3a94e6a0a85d66696f0811c5145ee62518e238941864c612d50b7a19e221c4fb993982288a65697c94bdb9a6107295;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83343d828c0380a0be17a597b9e43e85541218835035fe77855eb0133df2613117f98fe192db84d53c55ac1e738a6cc529e1a227b3a259774ce9aa6b9707bea7a1db611c3d8fd7c9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd13cf23a7ea3ca260283543f30bad4b2131b87cfe97f9510381cb283c2afedcea91e5712af3e311db2910e2ad2e5429b4288b4924d89ed7a7626ec4936d1c9150b155f4d4bf31d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2190b81dc68a084d2f1489364e6004e8e99eb816b342ab8f9667c0d1ab46f04b3d4f3bce3bde21a7b4f973760f615564f9204c14854938bd51785b853b91ceaa5fe9bbcf549660f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d9380a8207a73408c3d33f9b3872b46b537b0643f4e6064ff5f02317ef3999754e234ce6aeacbb74ea2a3e3cb74a3edddf90dbc4de4cb730d8e7e46bf7677e26fd30a9ef74c5cbf;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h995438235f1b88d33e2c3348f51feeac6bdcd4c36beb0f48304daab7074972ff5500e60b4226a03fc40cdf6fa70c29dc551e8e597ba4f8635b1bdb24a3716a7d7fafc686d1fb16ae;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha984cab26000f6d5b3197438cedc36dc96da696054b784eac04ae3cbdb7324910823ac23e8998bcde97e42e75422168d7239675ca1b490080657f67bed82379469fb918a22093b90;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb24a594ecaf69693a94853c3d73839e2ba0738bcca8804dae6660c8f5439c7058247abc719f9de5070361ee60d21cf2207584f23dd95b03581a0992b7487649d2b29e7408dff32a9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h202dc0a175de5dc18fc2bd5b18dfea5d54bd1e7f58aeb6b0c3c89fc4a0ed80fbc929c94fb665b3362b32c080fa0f4d79b97c173465bb5765a109599ff044267b4625c86c6a517696;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68502c139fb68d3a352fd33277a546b42f985ac66725e0bc660188ac84661185d0e192583a2cf292ceb269ac0e3b7300b700f2c82ae85ce8f086f411132e308f8b35749c5c4d2084;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71cb3f935a79e81d78e64f24027e6207899330e03a2550c59449fae1dce379096d9dfe5824b4a39384abd7e5a72abc8b0427d6033b901f6eb661727d66855a7229f58a0a46f4be85;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0853b958e8492c0093c16981fb14c8bf4c05bd2428221c611101b6b0c001bf19ac88d388917cbfac79b48f1a9ae999f8bc19646961da25bff8f9c75e1332902619313f2ba38724c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4392117ae454860335f4eea207c10c38e42316779d97db38ffd321b01cf32f1488371c39281dd6fa642e84eb8343d9e17b93b3c02144b318049f3b2b04a59a69fb4a3c069694f102;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habcd301695f86173a9c88d56236e776b344a0eba88a6045009baebaaede8b0ea64cbceb84453c4c7e04a4eebb721cb3465af24afd2597b2504ee7aaa5927acfc909c0be7db34d421;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9046db8c62fc43f5291ff9cb3cb6d5a7f16745cb9a8b6a35869c2abfdf85357a382425b4d4201569e2ef2d8e49969c1a19d2771169946613e89117edfb01cb8179f648167e178c25;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he356b3f31ffc2aff5c4754339da794dd04882136c40a8addfd1c59d954edacc2084fe09cbcaadaf922c5066b5a7493375f9f5f06e23f4342ea56d80040401beaabb130ed2e75ddd7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c6ac30737e2f9620087087b20a3a91f101f83d2cc9f638738259e8ac7bed2ec1be3f81b593462b5a276b0efc7b04bb1022f05c6b98cb8094031ab9449bdb5efaf0cfbe234f41e6b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h641027199d558ea5479668fde3961d403a92c6d60554004d0a06db35fe8de246e95ba43ebda08d2b77870e8fbbcd7c71d4479a804edf4178e24a54ff945c8348563b0a061a2fe979;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he80b610692e78d91707733d9fb04aef504dd76b4b9502d55e8b80fed9c1b48dab722eb8a01efcbc307385dc38acbb274c158d8965247df58e53e91cef447f581e0d68a4af108b38a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha6d3c8bfe8f7b4b0de8d12e5983b1cf45aedd806bc0d83f618f6e12a210d97386750eedc1c8d580148dc6b7268f219778a99d9c809c11858cc605d0a779158c78ffa452bf481e6d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb36395687868a17dbb40225591ad98b24d9eb7d5d089754438a83c7fe210573029b1783e926fc2329e8f7a635e8d111f44d254e69387adbfd716b8bf9ff91a296edd77d0a7b7396;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8ec9c820e3f512c9d21328647105de1db632fc9612a712493612d99a3f0fef236476f3d269a4152bf25f1b7b1dd15b88884d2ba75177de2e287f518e759f83a6b38f571f99cb93;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f2e4984d459a3a377cd9a997b321e55a5ff4fa0e57ade3ae6cb396c3dc17f528373579ae059d0705e48b2a72f3a454605e1e97c089c6e3faf1cc8ba9c48e4a070ea23de1397d781;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h215762ed200e93538fc6ae5dd26f9f1866cc45d2de19186bf00e179c25a42d95574939d80d7b42c1318d0b170351f06f8485178dd018f3353f2bc084f04c90d41c528fae930cb944;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18b751405320fbd3e3b2d1d77b7d133c4454127ab7ff680de1446741c3c885e75b6cea898ad825a0a1adb80951904ba1bbb77265e070a0e1508ae2aa0b73756488d03c2279d5f2d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e8820b1dc27f52104506c3140e8e6fbc478fa32f071e74caaa9f9c3a219b96b4f7848b80c4535d57288369c56ca6d7aed252527e6203c4154bbba977cf1f6f8705d6c6fb37f4d89;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8102b2751e84edb98dae5a8bbf3610c55c5fa2202d31bae5e2200497e771f20f966c3cf34d1f782c476364e67dd96d56bdfbfb798c52600701d668bfca55332c857ce2394f2e84c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfaba07748f7b5e3d86c3a29a63819c1b4ccc3d73080347582e03c19150f37baf3bb1458fab09d6f9f147f6978a9383c30e326f2465735fa4695d9b6b12bad8c45562e6d38d01836c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11a4844c333af779092bb1e479f09070961d0d99aecb23c3dfae4474d89106240975d47978430d75cd9448cc0a32fd1f49b44235610131c39bde42904535b29cb4a31ba0ad992bde;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf36d9e932719ee6afeff761e9032257db8e7ca54a7c1fb4fb58b7a07e106c98184ad76c0330927f4fd1af49bf06e27e3b8954eb54a02c1bb76e3c33e5d56f3e768df8ccad9bc297d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a3cd3cff41528887d48a7221117e6e38192825510f295483372c5ce2ec2e633f36df3503d3e1f7f403fb9bae8dda213391175a9a8902693934994f1b615c7efd1183c3fe2fc6e8b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc2e337f8f707ff298273f928b130083b2a91c6a6a3f37632b74025fcac74209a43c5e18c0ecdd92f1e6cb0c938061971520d7232af156fe76c7ce69f24d8ea01ebd429fc95e2bfe0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd79b46e4f19dabf750cfe63b8000e6538cc26365a95e4693b80338293e9c5df637fc5b7736a209ceee9428eb0649704011c13155a31263d7b96153b920b693da4b29c1c9d37c7a6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h736a3983883836c51efec45d3a18542595b99efc751c0a39cb40424deaaad79c2ecc4f11a2c85c3ca30bd627db818873c9c1113c2e558c5754a440596ae6d50517920a99c40a345e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d3f92dc7fcb9fbad18da99c4464a22ba28b4cafad2c00d7f223985a931f799b2a75371e09bb5c8400bbabb5704ddbab24724e730d197ca52df845169429b10c1f5ead7c71a6c853;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haefdfcb64aca12a35f12eab9b20d65f0f0b1c60e66f4de2f304f2abc2dac18919056849acddcf2c8e8e2c505e60c59cc3a4ed6fb105c0441a0174f206ee79e395241aea1b83134c6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf278a2b7d7e31bdb655a9c21bc6fbe28ea16e1e8f343027572edbe640ddd8f7f6f4bd8199fd589bef90a6453aa9541fe6bbcf16a30f72b453b0f0d325efd5e7f3f2c7488c1a98db7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h786540b099c3d0f12c3e58a8a1b522bd30b4d0af7ef967ed3b5161f67d80299298d0ec64885e513fe16d1bb3f7e9fa6ec2fe7318ec770bf136e43168e7584cf330566e88e88ac5c3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99a9b5f5c5cb7e16bbd093f6366deecd6bff8358393adefc4785de22f8af70ca583708bb6135409debe31d72cd742fe73775e0bd60afc57d8825c415f1bb78e70d81866ef5033d7d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4527f88e7f81317775564a2702de6106ac541d97ec7a0048e78c855315bd3c01eb74a81e0fe4216a89faabd742c60c5d699b9e11b44bd3f38b282da1aea927305dc8afcfc77563a8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6dcbb27ba548c69a30962b8c0cded2161618fdb0919e7f283bab44ec702c72025dc1da60113e48dd859bdb43eff6446be1a3378eaeb84c43994e3d1c263deaf58c0617162b23b2b6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he09b36fea1229b6666cd50294d2c23a0fc1aea6e158209d0d344064fecd98537dd3e47a38d98d02428181d2d222a3d20f22cfb921d6c68d071357f3587bb95663d5ea8f7c598a3f5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a68ad6eee27e5ae5b57a512c034d4c8f47469140323aab4eed585a0c63746b0c0f70db3caba018bc18d0a31a29bb0d56107e75b118f783d477096756ad66c6a46cb9819b9219ead;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h116241e8a655f216b63cd1800cc9120ee44f59c65286c68abb783d994df8d26d39ee2e1a4e20f6101a7f840cfa8885f8da37eb989b724072953e3ca11c50dd357f230b7157cb306c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c41585f2ba59caa921af98314fa544bae164938c0f30a8ff4ef193413ddb568cde402aba34d142f8cf9915ef2eaec5b55730fb98f1cb2bd72802de66fcb5b196ae371c91b43fb31;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee9c0ec438c95949f42dfaa4eca64a6247194e8b652265bdfce18a942b5e831204790b39ae535813e0171cda8da39ce27268377b33cd116191c059fb9e7d2fc3c97d4afabafcaaf9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52189b3366192bcb7728e2bf67466370d093d7e8a1695a93f0c9bb44109e501f8ff3949e9ca2d6ffadca3a98e721fa0c73856625b538998cf8f98cab8dd8e7c2d78aa2a2c27fea5;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72aedd35a2ee2514912d0925d5d488d5578187a1f479873d425a0cdddcfd87179a5df4b0dddc86febffd194923e32d8140be931fe4525d9aa0d4f1140525a99d8ee90643050ed82d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h977011e7d92a45db41a03d1c16b9c906f249763f53172c36bb9fd47f307d462433c1ceb414d9cc87f85455faf11aa4ebde60443ac16b2e83d6987083af931d8fcf9ddcd9beb04b55;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b9bb77ba49bd56418a81c5308defd8745447474160fc1a07315b3c6ed92943520f25db9fd5cabc9f3727ad91f96e90961bea82b3df4c43433d57d50ddb5c7efd61eac432915bc07;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf0d6f4800b441faa7ee570d553ee3e05cf3f8af3e7107f91b4d2f589436ae3ddcbe4ca95571407b71cf1136edf59aac36d8a2af1dfa59fa5052d1581d1c7c1aa10de5948b6ef455;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4dd51512b709ca3e0eeecbe4ddce5f4d10589f4d7ebe17358a1cc97e457c539a63426516a6f352ec89e10736b3b95f3a701f4215eb876c53deea9c68d42a870a46c9488553b06c4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h880785822e5b6eb30ff302d32a03401b1e62884736dd3a5bdfcd905823c7b874e394e4f6bd8b64e9abc80769dd7a2886f20adae225e890d3ef26acd85592e77b85c8738c261020bd;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67bc16cb3ef9dd2ac329fd59dedcf59947955001ec6591bdcf350283290561dbf7ce80759dfe42361779c2e2343560df4b64f7b076abd50f50d41b90ca1d3834ee0bc3aab06b7034;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd96dcfafab10c90ee470f8b3f4d14ec5e28a0ec62270be95e9578388e112fc76074891229e6bf2f4f785c3b62fc09d729d9686d22a9a71c0801b831f3b04034e57b0c90ca115cd5e;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cd48ee8bc1c04d93e2f66bceaa768433fcda2f1153b60fa3007acf587626fc5dba0919184d7680b8b18ce5d6131cd64d9dc5e4848781fc4551fe70d578ce4030067a369fa9a6373;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h89497e5b96868fb496796a1d0f007d04a5d671d1adaa600623e9acca39f910153382ed70625710b08ba64966a5599de35cc088f4319618fc2d7229e1fc2cc864b7ac6033a49c1195;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4be629c9b7ea764c5bf8cd081624d5cd3f1498cb8b344dd5b500a25db96ef4344cb34bd2d73866751afe58c06f8a2ef2a6ed040eaf78f4f647d6a4ccc8651ba6066874c95609c2a7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1eab17ec1e7036607c51c37fa8f3403906f0f84b631a870e4a4a307aeb3b9dd0227a8aaffce3c973d85c4153be0128124fd3d81384beee6e282325bdbb541ed8a2370817740c38f8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75789db46235d9c58fdd37ab28f5b16e220afac2a84b35e05fbaa7845003939475428a6dd3176aff0a5bfd6ffd0c829efe812f629c5a9e5c3df12eba109f1ef9cc66077b1764f978;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb644763d1905affc65bfa31e14a9fb86c682c8764659e2ed898c1e8aa3e78e3d13f5591c86f92eac8347847b070e8b7012247943e374f7faebcbfea0867fd457df77b8acb84b42f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a835211753efb868861540f55486c29eb2f4f9965183daa52873a199492f524011cb73bed0815ba17ca53723f81f46c83acf8cf020facfadb3b3f3b5daf79a0bf23fc34f26f1208;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd039c5e296dc14f52aa5e2d2577a70733a61aa3b45e36774910c60ed0511f08ea24f0ae6dc15470cc6f18a5e129a276fa2d7f06932c6e5429b5d2637b008abc69f3e4492584e4ff6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6bf704c41a7ff20a6527ce3cbf729abc3af3a7e312e3b4153bf3d08cfe66c91607e10877c05a2248efc8f622a61c8da25ee1be4b1e6830c6094cdc7559d553dedc0ae3d0b80e23a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87709072075d6839db82adbc2a2a99e0bd0736e61e561ab8daad6f456ca419191ab1971bf9bf3241bcae933c8b37a2156f8345fe8fcecddcc0a31611176a0a93fdc9c0c676b87d1f;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd45e7ec1c8291a3b3b650fd3f9518bd7af25c31bb30063219d5187814a9cbd1204a85e60a797b151a4869082859e9e8c3ad35314295e05bd395630b481ed3b62f71267f6195f9c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1646c4cd788d6133001c1fc7d233bcec8bfe98fc366cbb7bf050b9a27625dcf8b45ca620f9ab9cc3bf833207569d67bef44efa52f3aa3ac0163d7c15c846f35878a723bc49f72120;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5aa239c6df0e09f035041bf5212164473c11828aa423a6c0170b84c314ec7b05791c35c5b4b0efe1815ea721abb4898016429d26c3fb88a41303d1bded688ac3c7cf7a7ca27d87d1;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6a9a2eb68f84e664672b4a69b8a2f825ec5841e709f429499be8bc9c07678d55ce95e894ed3fc6d9197b5ffdcf165718b2140f5345b49342cdf5e1a57fdb353cc9f0e4062189439;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd384af565615ff3f3482a5dc894cb15412227fcafe1cdcdd3956923ad952377c83a5d6ac1af006f0c94eaa7cb770f1478abfe404d2204687d3d824ebb0dbde4317e62472bd0d7560;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28555b74768bbeca7eb62a774ee208a38375676f52f8525e993e260831253c6b9ae428135cc8fb73885836fbc65f9be46eecd8d3d16a08598f0d5a7d14339ef81528089a1fa8e5d6;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h461c28f8608dafd7d7caf6592057060754c1744ddacfa33860944ac89db5b3925e05969d94ae4f88121ee7a7a88293be46a9a77e35c28488f6c218deddf22e6ca453d37a518c19f9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c5bdbe748b6f39ab0f33e39394e70f8ca8cf78bd14ee5dbb8648fa771422a6954be57ec1cf34d727ed1bbb892d3438750266b83e82621864a2dd9d3703c4d0e69c57b30fef787eb;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9dacf6454acf45592055db50620174a5d8fecf06d89d2604d07ff30912ede8a787e69c704b02ddd9872b8983da898d911d753466301bf3b756ca3b2fa03cc9392d059e031c7ab9db;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8ad5c07dcc144af81584397b69d60557419279000e7b37c5fa28754fc48bf084780a4f0cb92937d24e96f7f907b56c4c71aed7ea3ac415562f844dba74bad0085cf0e43f4f38239;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8657dddc051edb926c86d33693879c13b72cd5bb1b4dfad954fa2bb1e9aeebca5faf7b7024643b1bddaf89c2e364d102e82a358ec9db005c71ed221ad7fdce60ec3698abe42b5d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd626ac5eb080d6c20290f383156c497bb775e5d7d7d63efdc65235cfb9f5bc706585c852537c4b65efb730f0f17fc6cc3ea212b2d3908a548497f26473ee0eb54b3f0b111f892865;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd50007b9f8dca170297d0a2e9eb155f2b2c79751168a1e7cf92a83245eac7e1a359f517c7609c4c25d3187a57a25a30423ffe98250cd0fed2b85e01b57a2af223323f2177c025a73;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b7bb825e9e2a8b24f7afb14f586c72da2c498b90e830aa2010f0d0408c207b15085fae8ce169506dddc7afaadfa0b7dce650b4a4767b218234d99d2ee3f75c28a2c80c328b8647a;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7938a4cb0ac4dd1302998969ad8e1986acdeebd16838c65cd2112bd24adfa97e5bce1d2e40c70b7a3c0871b5eb6f6ca8669e7b5bde3ef246247b804c170fe67af2e83bcf29a76ce9;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h360f80b6073e5690160ddc74237a30b5a2790e5ba408676ca1044d6c97ceb1cf8343d54eb719dccc91d2fb9b29d8e7335f8d1e778a22bf978df0013ad261dc6943c52903d369d467;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he71856d9293c2a7a7389bdbbc00572114e1bd5a72bf93752851e70727592e6b699fc81b849dd041d0e216fa4f9cdb572910a76100148a0ba05448c60e4ac6dbf71f6865bccbbb7f0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7468efd06a544234500dba217104835554696e2d8608fad9e8ff5998b867feb9e4040f238860d7961bfd61be7c49878379d96c8939fc7bfc3bcfdd125a5fba00fa2878d68c59b432;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h860e963544b035fa31b25ad339a6e31cef068333ac21c45c963a0eb936db7f2277f3f4596dafc5f708e50f899f57f08b5eff3cd464325bbd661b5764a1b03049fc851dcccd7c01c7;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2d5aeeb5b6f68270bb716004afdc7e8aa87300ade03a949f6bf4b4d9d2b2374af5886df48a39f919663ac40a57d2d63bf34f2dc6f38fa09dfda964d6890c320fbb063417231b551;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h264bca87c5adceb613df2fb60098b122c268dda3443dee17aad60da514d3485a539238b04839c2bd88d67181b46c6f2945b4e303b16be1a147e13c79861e694c57e6169dcf0bc7be;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h689e1059d5ee814446741e559f0310dab267d5ef375890a1093af56a84321b3b2df7b3fd0eb27b398f8ddd40c95346fcc0dc2942a3e66c63731351424a8b89c77f168572ec99a17d;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7dc42c7acc92132afa390fff377ff5bc38a26d2fd59c2033d4fa90706b15d4a20ad43cf2487dc0407a887b8a8a60bdba11b491e802255117046f4597857e1d37d44a94dbbaf2d24b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2639846c4ddf0150d4a4d54cb9928ce4479b1fcb25f7ed29220f89c8e2c7b315b8136bb49f9e3f1912a386c7f8f7badd9de8029ee903daf2b1e70b45eb8088c97741cf36a35224d3;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4fb3f6eba6742b77fed50a63405c4c6ebb375bc4ea3d15148ee6a9942d4d4a897e0c8e1a9eaf83da8eb1e260be9ce75cf395bd9df4e0b5e63b4e6721e130fb5741a1a6cde9415c0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9f5c5fe78534cf14323b3ccd9b614c64657baf83ffedc81a38808e1b658c939e0fc0200666201501e81cb6bf99cb56e134e0963b983e69ac8d9c1ac0b085fd110ccacb8c343f542;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d4c12e7f7eb6f50894214845904210769d36712df629f10c3830ae26472101cca139b6f49fb7baeb4cccb6d4215ab770f5d10f5a7fb4d84212f257ee580ed68871ef64865386972;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b3e6f28509c21412efe21eecf16807959231b27e665ab23e0ccf178fc5d67ff90e8810665318a43766fe7a18d760d226030915fcbde45f6e8140f4ebac3af4048007820fb8951;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9272dfa9d174ea8a14e578980cce9a4e2360c2ef59e24082b750326a04b93336ddde22793869783f291e769005b6f0fc6847d0d4eb756729bb38a75a2d8e968a3ea8028a0038ff27;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h284d39aae5a95c9fb8f1e2a0c72ebf904ad3efebc620b9a59e368ea18aff2b5eac7395c2bf6e69f32c940b04417fd8a683693535291df62b71bd9dc53ce1017b3624bc1fa9cca69c;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5bfda02a107e487b60bc8c6a785da53ae07005de6d2c1c0e596a4ce5f552386b4dc2e3ac17ee82e608f4d687a8935a69df1e00502c3ddc72e5ea03f41fe7ae0f40bdfd4744ceca0;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44b3804e8e278c58e30bb0135def12e2d5050b9dcfbabb0665a15d578c889581a1e09a875297de33645fc3eb5d9a22ad33a542bc8e795dfd710f724f04b51e69b682c9a4131bc1aa;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70157e89c4c6dabca0a71e1c37231048c241bd6b3665b9030c6bd335fa3733a7379759093270103be71a1a45c42f7f67b876b7fa5986b8e4c3891f3b0c621605f55c6aad7d074e1b;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd866dcf4e01855b61d2da8622dcc3a7f3b54cf07ad41131c2df84d18df118171dfddac0c4728d1ea03dfbdb6ab5c3de6532c7c762d19261ef544928efefcf890b396dde2566b89e8;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he15005fa3de5b810701d120f9aca8c0a679178829c97064d21550e40e74b995c95d204179b67c9c94e0545a99f4b8614148e83d33e0dad379fd2110cb87b2e86b298f0c45c5e51d4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbbbd3eb73e117c87f9fedde44f4f37b023bad8768278ceb907115de61162c425395d395d20b4044ecf7868a1e4a585aebafcccbf1336d54fc583af74c21271187e80f3bf61b1ba04;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h877130a6dd4044a19c23593a3cbe7210867f2de057827c0b96c03e6eabbaf1ba32beead0aaf4922f14bf9901a9077f228e9bf5e0d9ed27fb15411e96cb2306932b091f4ee74ffcf4;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb300d58cfd7d940b4cfb9fcbbbd156b18ce184ce3bb81d197399fc148ed18812659424b12acfd64bcc8316399bd5bbd8ed3fad30d0aa8f1e6b5c084487b781ef63c2ac8fc3715c37;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he01c39ba5ef8f8c9b2f6200ee7aee0ae9e77217ed9ae217de8279f6a930c4d58e2fe1657e2f66c19181b85eb7ea42bf4c64d8d74001e136f84fcccff27d01d60223eda27ba4f1888;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd6cd1730fe446c393e6ffd4435a3862a9a44935780029e356cab13cfc59d6e832a947385bc62da2657585737a7656baf3f8dceb1376c81ff1ed76e3752b943a14c57b48dd5f57e47;
        #1
        {src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2a9d1ba9fd2ff0709ee03ed634609ec1a9c2633095845c05117f068fd5f81ecd0e927165a68155cbdcc913a34eba50d3db3e989b38fc7ff6e2eaddab757b66fb1d151395d4d9b2;
        #1
        $finish();
    end
endmodule
