module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [36:0] srcsum;
    wire [36:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6857c8dba25263eac18ae1ad54495dfc893f6b6ef2d757fb8a50563622d2dc62fa041eea9b6a5f93b3a41f64f43ea02dc755347db07e8565fcc5e31fccd8f79f9bbb4902ff7a9c95ff51e4fc33020c4a781beb0249482fa124f173cdcbf0da22c5b8ddaabb730d680f7d809c0cd20d5b2d27bbec0e62670c64ec226de7054a66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8357d28989c52434a9e687661fcd7565af66f293af58f68a4c7a98f8eb46fb1b694de7cc745d5eb74bccec2724be9233a3023c9c7fd0c2337b5813c59fd88d3d235be6785168cd0be8517f4e9030ca816eb75ebc2fd56bd41bbf79c5ea994fa7302a705f8ce982ab80f112abc8731173a0560d4af434e04c4add86c586a5c86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f8dce0537c45b874ee2b0c67348c9a5031c5e7757c01d88150a0dfefaddff7e0486750dfbd4be74822680fb221f765ca9cf18ebf42d71dce8a21537afc190a57054551f42542e0e6a8d55adbed4b2e07b0342edae304906655d313bc525ab4456be30ca4a9414786c1a45f19e1ff3dbfe23cd46b8c00a08a2b7550258dd8c7d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15683b687ac5812a472287db789d5a079c93d49dc8f20e2f0535ce2668966b03f5873c1593aa3d02512688a5ca1c7562f6ccd844da5080abc762f372bccc30ea570b6b6e81c9f9286c9967da0fcf327aa0bbd08d537b7e0150d79254adfa88bd8d835cbdfb6c552d014eb43c1833776d87ce52b4e699d40cb4cff8471f380fde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fcbf97188e2cf842631f8414b11d446dced3c9e6b9e66611d7d5b634a2e8860832a20a966b817eee4c0c148a555e524f43cfd0a70b199a07e7fb45f78961135d7e7f71092282fae397a92f8e6a70eaedc9df4f2ed6ae10f34e4f0370cf98da5d5e7ea983f96e7820584d217841d35751f6b52c702ac4d4761ad3dbd45471b26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1889bad77940c9efb09d0d372d7b095fc0d420ea8a5e8f6a580f27c6fe6f0929b1370ae90d5b2f4d7d576382f91cb24bec2ec8a61d9cf08d4bb93c4447a359146b4a12484bd12b0631ad641a734cb7a1829f8534c45ac59fa0391d8e00e2720474c5037c03133e840bac774d1b205d0366110a34b5e49aded4f9c31604ef82e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c880d5e91fa277c1c7207b11acaa62f3455de875b43b1c90a064f1d0c08f45c5ab717745a11b3450ed992301df4657db3f28457c8f441131ca6042de50b274cc74b6d1dbc2e4e6127ca6c7ed6e8efd3a273353adb0929a82b116e325dcfb5c3cbc5f1d1847aa8e80989db949425252b2188b69ab58af9ec0c00c050c4d87ba5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1e9843b1eca6ab70971b1957fa4ab5b2b67648abd62fd08b020569874c2f61bf43ad89668dd9e54b8d3420dc378a4ef5379b8903a490da21c0b4195d2646ea81e650db493a3b0859ece265a1e090bffad9ab755850637e721116d15e8a9259c4abfc41694367ce17312aee313957f6bc3e3390648669823c603944479293b03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha867a7ac0c0a394b484fadbe701464e25cf26bff55d89a8630d5649604bae050e828a69d0c9a238eb17c4c8628cd8f3fdcb8523499eeff6030f65863ae88a6e8ebfef7af151c26cd13b9e7324aad68a566cc49c51385ccc2a8bf01010abf6f251196bca608dda396f2d924411af90df698151d61e497b2dcf20407e6a421845f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6bfa72db89070e9245911450457df587af4c25f45019f5b1a6ba7b7e5e9255332de836685575ea73a28b802899fdff22d815b82234cc0a5b4aa884eb74f7035e2b51f22a2238e20f90fe3177c7ed1b1713bf94f5f8f73708644178cf8f84224c455a5fba259b9e1127bd613d995c96c9002c481317a024e8684fd49371b191f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde977355c94e074e8e5302e5895eb7eabf034766a3343df700658af77774e1d19f72855f25d23f03ad68431b3966ba99f1f72459bf7d32119b281275651a5e2f12eb4220d1903f69271aa8c69b87c38d7713d91f9fe692f14554b528ace7d2c8292e2dfa00c454ae205fcc7e618993726f608a03213aad78cfdc30b171b08c5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf69a89222f23da7a3d36edddcf298343ea0a97e4f1ab7bb72b03fab664d01f9c75057fefa5bfb12c6887a0e587d1ae86dc13c999f5c3f7c0e3b916d9422146d713e63cf193610936e576b165ddb1448dfb48c9681f08de3aa610880aea661552bfbd7769b10d788f3c46d29eec050803ab49003e3325b803f00cac5ec3a45f4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heff42180ed5e76144e95b86c072855fe14a20edd80fa81284108b55dde1083967f3182e8d954b8d1bc9dbde1e416090e906a863a12fc2f05fd1fe835584eb873d079d54c70c2bb617fd70e5d099b75fe43b12f6b2c2e318027523150958e10ea542b78d4df2898cdebdaafd3d1f611abdd311372726af6747a0b219db98bfb23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51258de7488d8480e4208e3d351bbead837dde356d8e7990f255a2c44c8a8cac881c34a12658279a5fa7383da4e0a73a3fa9b88df691b7d070409ca4a71b32a8594079f6d44428c318689b383863eb21f0e2b84351d7026513d96a64441074a8e1d79a4d5b7dcd4a7b56abd4c98825cc9bb3ac1dbe24d2675c167c825d0d1fea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd4fc99330e03d5cf55bc0d48dd97495ed6bfa6c2fd14f53df07578b50e3d102d7d6f27c2bd61c1b22286d9aa72a58f05bc0cb84ba01406bd91db530be8e5f5aa032b067f792cb80a9059a182059d47c5db44d06ec1acbe71c827638c1ba9d395ab241d994932ae17de393c3a9173116440287a47b0961f82ebf6a3f5bcf3c24;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h518aada9b56bc815b81a6c3be86b8977c8a09b598b2fd941ba5aa641160986b7315ea863de103d7d4fc43a01f73e413f2ca04413a31bdcd8d9363e301d75bcaca65fa5b84cab786b3c124b12c148e1fad91f5ca04310821202e313223992c402f4404d611c633f337055876f2ed531c93f4f9fd2c9e42b1599e0d62aaec33619;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffd2f772d0fd6b86726fec680277f4347b3af3587427c57ed7bcb3742abb9ab945a2de87ec4c58617da232b1fb7276b69ecde86d47c29970b69e5c4c76bf1949dff59d98624c920ca51d505c5e4fa8c8ee392c38fe89d431699b37d9c6e63e45efb1cebf041757b56d7d7fff11754714296ac49f895212ad37b03d7dd74dfd7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53f1609c42371a3ace99c76ec45d95946ead4067dac3a67bca07f81ce612810b36915cb2fe11744d8817f6b0368e89d39430579c970286286461dc5776f5cc5e748ce296bedb8b52a3b777a6d8780959dab829088f3db867015ca3f82730357be3714e94f772cf9e04de21bbb0e46a2c6ad839f3d6d21588f6db22e7ec25967b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbcb67ab4c4b9a50fdba4882bdc499475905c28d27ed79ff47d0e85834c09eb5e97c6c75df477b1d4ee5d2537cead18725e0e325c16bd620a108366b71d8c3ba7b9399baaf43327a4d4e02a1a1f1ed90a36421656d749ccd879d77ae0a78ccba722f9a8ad7c4e45cb2f2fca1cd2a8ad54145a9e3fc12e449a4a6124aef7747189;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6de821e18d7eb014208e6535f41035f9a13e1a1e33f4c4d637bed944ea8d7934f12bbb9ab44a3829f8420a5623a9a6e0ac9211d2bf7ac83ab9d1f6e12be620c6fba007def69514bff307de5a9ec45f2c3f1eb14082caefffee5c2e2603d2b8921db38d79d8b8682981e83abed72729ead4dedcaecb92471600560ad4d9abd9b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9150ba11c88f729322614deda609ec3b3df6b2f883741ec35930cde5480b72f74ec98cffe31e3c088e79605e7880c14b7f8ed247f91a2f45676e1122c369c2488368e9a44a751861954ba21f8225cc1d1d060545e50c22b32bc98f6b5f25cb67ecc961e3a39bb2cdbc6f894c9960b875ac696f7a6b649e43fcd61a0e3d74d7c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h279cb686df64d350ff4f8de5e1451316490fed4f1d39408570606a9f90a7797450cafed30a7d68fd78792149bba56d8d6097d2d1a9dd5ff50b1432399bf8f29f139435fd1c88a3bbecd877a7501b6c74dd60853584272fdcfc14e63219179c0bfaa7fc5bbe98313063e548c696d07fc93a02b7d1809bb8f6eb512b42853acef0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2b5a1d59681b05191ddab868cca85ca18aaa0e1284ced41189cd247cab9cd06a42e26bb847e2a8ecf538641490272792e6f33f85f8a45be5a88c5c3e86f6c879704884b527da470ca88b4e33b9f4c94aebbc14dce5e4e5d6671fa4a7eacb09e54ee1bc82ebaade457903590f984a64eb6a205528b5fbbc70c7574c057022cff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ecf55ed08faa0d868945fa5505e402ecd908d36b65ca7515cb7d1f9efafb3029e704218fa1807b263d5764e2aebb557590811f5cd4a9a0d6d1c8d6b616f97827f5d72c138d62d7821fad8b5bf0d3b5199b2e520e9c142087a28660dabe2264e6a05a15038070bc417c9399ec9982d1bc166b40699f980b26cc89e7b831aaf45;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h833703f03be66e301a4b16ca72e0744ff0aba8ba42bcd2f40b0eefd44a8cc25a4b4ffaf8e2940620b0ca1d225bdd7e34fb57f49b6e67f2439e9aff82192f3378f4932895ee8ac0570752639a292c6bd2e9d91f44a3c13bd45012be83902cbd267ff6b6272540d6e17e92ee1b9303db83420e175576880d8a68102fc7ca6df7b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7fa3490bc8bc4fb1fc8a7e5d129c891e19b4d3cf06e882551432e26f062f1cf10e00945abf65c5154b725cfb8964a0d35fa897f0cc7a9816d4cd6e197c2324d3a65cc6c3ed713dabfb82791accd73b4c3a484060af57b0d7a790cb19f24b01a545b5772e0f0b9c20a77b48f780a418db11f9f6aaca86c226973d5270e1a0fed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h627e665a85257e164db129f2dd396a0ebb64c79fc0ef64443972c6388c68ccfd7a3687735d1384a9a7dd0c81f7dfef42841e4749ac9bb56635b272bba0ba452bb1674b86cf5020326d46741f1109b808b52147e712c33f83a9fa7aab735e7ae4ce04bd76ecb764eca710f236306fc128378fe98f090397fcb4e3c3a41df079bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd50db5b4643209b33ff168aa56d29fd448d6734b7e09bf3871b9efc82d0dba7ffee96472858b3c409400d61a33f6dd63ff5ef8b865377d5d321e330287d300fc9597e56ce49659f72154250ab775818d2ab118c212bff5715a1d2720f3de0625d83c5dcbe71f3f82c01d471ed446a50d86c0a12272634df46a996fe67754018;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h384933dc56379b17f8c4184f4cb2e1f48cbb358ce687b2802b5c8195b71943820a067ad2b4919389df2f5e120383da44399d12c638b9364ab5c4ded828d73cf60db02adbcc7ee564ed95a053633b99ceb02698be14e2779548112239bd68f21502f027b719f3eef60593159668ce8f1fbc95d58cd91971e406d00c130f1c3325;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfdb8c4e6007cb0ab7ecd92db93612125ee470f13b6a68e01bbe9a338581b05792f835d9a4e8e4d9a47d83ee9c532cf8c0a8cb7536eaf80ab7a2d67456fec5c6c1a076dd83a7b45bf84da8ce9209a4115967f5d4a5cb3fd01a119c47075484914cf2f259839ad87a0567c25da75c0a57c36a5e67d5a0646ad04006c9df2e5c29;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h372a909b1593362a48aa15a2581905b7f73794bf237310fe5a24ab4f49438ff4d72e60cca9425311fc2ac678bc4fd6836ea708225608eaa76a9439bf441902b786e74ca0c8e136729837111dca4d8a1e3f6810285d9ed5e23c763202dfa7fe591c368b4238b8e7af0d6cb70d2c01ec952661352a8d46887e6e5e025fd577c5a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69e44b6f56206d7025f71dc75c40a223c20186a37cce8c7c7a567431d1e6df226c95a5b3144f8d073d44763130dcfe7a3f13c275482867b3e6ac3bafb79b17b73dfec7ab8c3698879ceb63f0487511a80dd14e2d57f1b6eed35deead8fdb633009ca4fb666323444322e1903a1860f3c3e3123385f79aaa4e0876230ade58d63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8610e17c0a2b6fd73f10f4c88674621cac4aa13d93db02905bd2ab47d53920aa8ab27ee53cc7e9af22de872068dbff3d442209f3f5163bedf8031d3063c7b7bc34f002c4c88892b691cb6fb58922d1218945a27cefea5abbc0a2531beea3cfb72d50e3897ebd1cd6d14c2f5aa8718a8eae403fd1262cd28fd1fbc2651d37abac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcebebbfc475f0a569abb2cc327474682d08f2f4c095c2644872532f80484e0ee507bd1aecddc93b328b7bd7e6af3f3d3978995e0a2a6b04b0ef179aecd1b94e020da4041c4354288cd1139b1d45c0a17b08b3e10b4d8b0825a8a868b46398d720b357b9591b4a9564e693d2f107f4652b91170310672865878481120f91d13e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9b2ce9a258828d7ab55ee446efd8b12a9213e89fd59a7382cdc7340963cb980a1c96b1638581a952e7224e022f2a5c03305de884b4cab0d614c1839ed48e6a2765aab67cf0e009233ba4a2a460e371ac1b4a706e7e2c08984fec1a3c8470077ae9166a98b8eeb7efc2a4697c8aeba803dc95d2335463265dd1cb654bbb65a86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73b480d20f080f56c54da2534d7458fb76f6ce5887d714280b8332704df8d9aeda862f3b4d171e2b862e6271e83f47ebbb0e90c87ee29f7462e79fa0a198fbc1d276f3a1acf1912a9c1080d0dfae72013206e57d61f7752e8120abf884305d9809eb59becd050deab3924200af1a099515cfe67e71b0d2d97447672380ba415d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ad1d17dec23b77b1d9bdb912f9ec47d4bbc0f74d96ff4a158f2c19a88a91a13d7085eb4ed9eaa2f9c18fc21fda9ae55257f1bf590eb8cb79cee4ea193f29a353be0706fb9f4a02444ff23c9d8aec267a18d85c470bd4d901e3668f69eb5b1b324ed57a74697ae29720ec2880632b08d60f4836ba2fd4d06ad3df5b176c0ba1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6991d3be69976c34713f6ff3d2d52670f539265c2bc0c72c4983c869d4de2f95bec9e82fed6bcd8c1b5e1e21d3eb3be85e04413b294e63f38465d9eac52ac704ca82e93e7668b5f5e3d45ab10c91de11d1e385d9b86ba11bcfe9318514a2404027b85419b6f7c3d234f53d2a93d8d68a17c916bd328675fbf6d6d5bfe029a2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95ac87550cf5356442103ffc32852498f2199b58bbf71284cf2c058ab551cfa81d4e9967b3a2eb2d5bee86d5d02abbf2cf1d2deae9d3bd3a41caee2809e02f8e605a740707300c17e993576e8c45bbe733229d8426a8c4de6e6fa814f48c7687074ee2729475c561dc1129f6cdb185ed62c7737c2291bc26f49be007b2b633f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5435304004b920fb7200af8e378f825bef22b48ad8840fdc565cd802a1bbf948ea948891801da9835d8e1004d6d997aa8bf84a32253806627daad68ebd2b3a59996089aac383c20e08ec7b2fe6e922c8e1bb3ae9be6ef6e587737e1025d0b3ef7a9c68975ee2d5e4da04388e9bec2ba2f760735a8f1888278dc03a63a0ada8cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9780bd0b1d8ba7a7ef0580478f3133db8d3f31c08077b1c1c08ca4db73c757ec0e69b66f611067acb6afb8a131875e1294c2bddd55852b3964021b816fdad0c10a0f7854b9990de97a8f7e1cdc480954fdb70949b3eb84abfe10be19703cb67b23b72e4fdc5552fc8ba553d7b4318d850fadc83f997594f6f8ab20e1b117a511;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba7d23277aa618327dbdf5b539e65600a64ec2a3f729f4c91337001bc72e3867c969ec04c77efd5d8cc79e405dde397691714e3f88350f5687afafd4ee4281c7f64c513f22a793fa3ef4beca9d0298ab649740f9c366c37c53826d7f7b25c249871a7b429f19a4269fb5827cf2f72847c328b32dde515f1a74d6a1cbcc93974c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27cd72cbc6ea98421f4d3c4a488c387563abbae9708374c206770c96d719e04968d555ca840c344e5bcdad684c622a9eaea000572ca4ed6887db418c6bb9051cd57964b685a209e2ff0c684f7dfa11d1186d7b49ba3e4aec5b10a9f3b46dce5b31e29c6c9eb5effea76306433b692c76a45f78521584814124e1e2e4882c3408;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8583cbd3941310b2fe9a990ae2866cd2efa8c8a5b3dc76b71171c942da07df9c8e3a85df87b063d674469ffc3f5f81336c7e797b403bd02e6137ab64aff68872a090862e6b685759a7c96cf3aa0b0a48c00f338e651b4feb356e951023a14d2d4948328fdfae3683b5cda02908c5a7d5a49b17e7d33df0060fe22deb5f072751;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10671b108c8a572f5c2accb25635c283d14d81a9939022032dba4769edb2554c75a1d0c0b1bfdd0b4a28df47f6ace023e77c1d4addfe3af7b277f55c8191460391f131ce45154a82f7f8b3c3f6112ebb4ea3fb27df6691cf2b61294aa6828f9832e652c0e86d89fef352b4f6e62974e986cbf99d5cbaf22a8885383dba3689d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94aa9cb325cab25aaa620198ca597cad3cab0c7d0f126b5edb4a114630775f9c56e1e63333e4837c130f85c65ce8d5f4659aac747537e3ac7f12b1078906f82fe245e760d01465611cadc8acdd6bfc75bb959a9535dc13211ca6825eff8f01eb899e9bbcc419cc2faa499b13d5cd0f30cf879aa74b75c806d5c0ea6ec0c5940d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e0eea4143bf9e2b1b0d2a0b569ff1699603ebf50599ea4f6545ac566c2aafc5bd6510dad525951a1954c6f1674543374603aaaf7db22c58ca110879ed6d9c13add5a8dde4ca0b44014d7b3dd2408a82660a3a70ebdf3ae7d8ebb4c04528087e0e94c96569c66e46a9e8c48fb52c6deb62bb435dfc2bd7fbd090eab96a7f7a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h571b9c48001b9b5a4071595fe9d606ad45648507ebfcf5b0871fa199148f521d47877dea01af87d68dc1ec3d924d7dd2287e113c59df4ce9c921b4f61a69f868b831edbd02c5159728393c23608df488641f8d86163bee288443c0ea12ed4f5752155d52b9309dfe8fbbf0d8a896a16ff286437b877e9e715920d4d7dbfb7e93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbef2daef9c277ec7b441f343c633595c760e978442c5ba4e38d09f988127c5984afff6949b7efe5ffac41c665754f1a03dfe6fe23065c58b88a346e2edbfa0df42c47e5103fa4cbb663a7d01d78e9c7fb114be22bd7f0c5bcff71dd2d513fe52d57553960c33d76215728454227d7645a081343fc5aec33438e89e9121592a2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h275ae282a21f2f9c424a8ee5a2aaa0521517e130df0763d66d0c51beb1b7f5dfebdf44088396b4e8e1df49e76884223dc8db4847fd0c239f342aaf2e637d770f3dbc90a70acf515a3422848e02b08f5384a20dfa06b65e9c7bf5356d0fe2fe3a7e718e1d99603afc0046f3b9adc7bcfaf6fc5f67775047a354d975a31b61fbe6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78df9095f7abf4f4aba98df96eece210c93efedf37e11ba5dbb3ef1b2ed6923f2c3f5290decea21715bac5a16c4e018715b3e7a6d046b7243e18bf7294d85fbd11df9f765caff414b857e99a5c433f67655d16b769ebdc515812b8a78f045f220906e1ae0f922d77cc36d782ea91bbc19a0f53e0167bb5d812132134f62cba19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44df87803e1e3900882cff281b3409b33327524ece2ab6a2c9b08d026f5bba6f9c481de6b70f6b0a43345ed5791c680e533dd852f8a85400c2faccaf7a0646fb35fd05f4e0ab30d4f6438b55a55392889cf3f55138f2baeb657a297e0daebe3abfad12ec80901b2325f6b1fc123cf8de6b6d703f01fd52ab9a34b5735aada39a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b7b0ea6659a4446c9e48f290841c7cb679eff36b041995d2f0dbce482afbc24397eafabbdd57e989d43fd34cc0a083bf30fb695485d7b66f07cd3f6e78726a592942b41dca19fa0f3fa3e6fde95dcf330d09e38ea33990699e08d45169105b475dabc76a732a087ea152ba55ae37cd31d6d41a301889f023a948e3d642fa640;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80f50a959c3afc774b2f26ec4b8fbd40d1e672bb1824af79a72a105b56294c8a4a8d64572c25eadb4b3e2a2d4b57eff57c23b0a3b3c183b16b3dfdd2eebaebf071116350116256584c76bc063088e03f2f8192b326f1dd889bdd4090205d7ad77752a33f6d20b6c4d3d72371c715834455eea09f45a051492c6c4fe3719c8dc5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf03fec5dbc3a2b78dd852274daf2d501f4d81d5790207894e772173fe5933c329fbc82caeaf010b7c8b3e112df9bfb374336b664bb2cb0e2f3fdd4688ff5f6927b6951415d26fda081c30808cb5cb5026f6434d0e5b9167a4c5c333bcc90df884a83382f8c67f5e2c8bad0b71cb86125566791f3e3a4ddc6822c92ed9774bfc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79493c1c5980f72216ddabd260aa6c46ddbdb59c9bc42bad383520a4a6f7291ec9c5afb1992da6879beb5564aec0c560768e895e52dcad995e4e434cce2b0eab2195895cdb1c3ced811a742228c2c37f4ef026e3997d90cc07932fc394e10521067b31ea048fd30ee59c881a19307fe45b73840bfd5dc4d7ed8c882686ea14ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58265d96fd5c8241519991a4214ca3b2417032dbce171960cfcfc589a1df699443c51a7cdc962f3a80d582eb1a07b19649fe6653802e064ea608f0ef22f6372c0e04374390e2fa9875e76436c503b44ad156e1722fc460be5f86fb72fcf3ff742c0434f81714d775633f1a1c1ae843c30381d22cdd599bb6c7c2b40e50303fb3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f05fa468dc7f25532243057ff607e3252259db6b5af3dac3e09b3fac78b0b1ca3de44c094435373e06f5a933835749d837717ec0b87dd92091f9b8cd3b9067eeb7d009189c216877b26cab6056208acee9099d8921d9a5516686014d916f6cf535f4cdb48ed2de22e0d2cc3985b2fb98c38a66c7f6976815d35a27659ddbc70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4294d45c6b68f35d907a9e194b09a9bb3f602b19bdc2296e26fe33386b383505281228053c096ecd1a5b1ed13526f2e1e71295e58f8f5b388faecaeba1d89a2cc4f67ed16722e389901394b56cf36abaf8ce9b1ee183a84b749281b8a2d0f56744ed2dd2bd50feab1d6a0aa387b4266f370fc5c4b2c0728b9659e7df3fdae3d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h938b66339d7bce868f073de454f9b0ac426c897a2bfb7e6f2056515ee6b2d0c1c108310fbbb241f5b4d4fa37f4ee4f9fc2e6938451644362caa22248b01fcbb57030806c97b465ef9fac82f4c6dd0ced44f4888365cccdb52cc32cd3e37d09bbb181705c28f75a4935ed04f6ce0bbabd8171f21a4ad89f6e1baf6192e882398c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94090a1c59f040b74582b6ddacda17a736162a1bee13d7f13be7a28c5c2cc011c56e143e6d36b9ab1bcc8c87f18d22e862ca98a295e9b40ac2e8f7355eb29648cdfff8eb84ea26ad4c0fa9d7ee0c7fe8775ad19ad06be8282c54bec0937ed5e78fc8e8bb641bdb1d0b2000854c97d3e44368d4f6a552f1db527ce54ca94c7bd4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e8f8100a95d9d9bf61404cccba02019172fd93962011b776b6265a74d7f2d44393431cdfc2dedd3c09693865cb2a4783e476a6fc108326ffc1c9c61277168757428501577bd16fddc8069782c003155ebaa6865f81e647dc1be254a8145cdc558c91738c2acb1a3795e917dfbb920634f75ae9f4ec073b6323c8f45b015ae28;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h754a3c3e18fad9f0582c2ad0471d7693447309847f90a8da0fa8783bf8b191aa91d84d811c36fadb3bd0ec3093d75785110dd49a58e36a4d005546282843a7dd2879a48af460a3c028b8138f820c6ec99d04d11058d915325d6bf9393a518222bfd43e183a09c362301d24284297c679a7536879d83b09ca956f2157f8476f08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45f485877bf51a5034e090c36a3f2f58fe00634df5a93c96df7178794139c83514dcb006dd84c0f85fa1c03bd525746d1293ca62d299807673f4b6c5c5d89aa8d41a9341ee8b66d7c869fb894f86fdaf515e91ea7512d8f31bb9559882dc141a6bb3b3f08db28b5a33729a95ba24f5e149bdc8355775915d14cd86e335fff65c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d61975e7f1c13bf6a2bc1ced7fae1f717d77eab70e03b21ca650fc9241309bba6eec01022611cb4b48f55d39b89cfad3def491270c2191030617bfd0874cab588a49fdb7ce449558c58a1f21d89eee2a05e17ef3c8492bea74f686364b35f8d777ee68b7839ad28d8660467f08e90f273366744c234320418a43e70fcf0c427;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41bc863c1fdbaa0a87b51f31476e2bb9c17b4aae054877b8604884940b161d620384fac65cfea8e44248f6bab620a74af101728c45269780edd46d4e0b748a770100d76e87e4a59e4da53e00923553b9039eb2e6d6b9eae5d213bd6268119e41e5779a7ead06fdb3644e1215861a64f2a2e7b3838a62f59c2344fa2b2c259f1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf95614b5ab1e4ddfb44d5d800536f98457e530e5c998526156d1df0e6dbf10490e10232ad56d46ac518ff3d00ec72bde2b91399fa6d557b26dd8740e5fa9db4c9a1073f900fa9a2ff7ddd0cb735e6fcf8b08cb488df2faaf24d81b0b5957cd1555cc78cffe857222cf0f7a35ba2d82893a3b3d2f1e5bd9761894932589fc5907;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd51c9203c9616648326a48dada540915d8bc0141bb8c81b0f7a43afc3e3cd2610ebf14c38cc41cd8eebf3544ac86cd0e6f30ad4719dd4c105ea3669f1f5037a6ad8062b20220f1ec5c7f9cf2c474c57d5f060a6974a9f5f89418a5d05a20c5ea7fc30fe05345c46cb3a54728bf7531d97b3650eeecef345f0d983829ed7ff421;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebce24641dfe14d93368299e4740e373b098a4a8a134d9cfbce373f8808ee53049ec35357162dbf9a9e90dd4ec9e8eb84a0923c49c56f7e7756f80b14e8f2722bc7be0e879ee8472455a66751bac9781ad41b77f35bc7b865dfa73b95f9bd57d400fc391f667f31a4df4c9e135af692456c6bd01d0497a8640d75b5e1cf2da0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e75358204753a1ed72dd43e6002508fb7b5cad1946522089e36f0e7e6d7fd6c613855d8b4e9ed6ed137aa55023f32583d141a2ddbf14bade990a8882a5515beeda1a0d3dc290e70163993370abfa287a08f8c5b394cc1de5ab3fbfb751412a43736dbe8a35c3f1e3f4f8abcabbddced1b29caf2a6f0a12250eb6c98e97f8a3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe7e1258174c99add99b72ca4c7d28cb5537c1710ea2d3a3a421f2d2cbc7b2d817f5bf9d32a9b94f1e9feee27e51b400ae6716487e724faf1c13670abb1aa4dfbf7e9e3e5a1be6f700facecb1aed6430665e1365c6289e53c995ed0bd6e47937653139f746f89e3c8f446f84c452cb3fb72c35d7a9e0da10c1a6154b4e0c84ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d41f4fe5449ca71cdd3c1157735eaabd7e238de0a53384f78cf0bb3327183aab01094225e8d165a0c0def2fa738e7fc0c5d606567859eb2ab0623ae0368a486fbdb144d235f8c69fcbc58f406a62eb089aa9ba95f81d3ae34e2885496d4e2e7b76bd32a67e19be220117d95ac39e0d4375c92dd10476c7fcf25b1dccc2a0d96;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cb5d337967dc068f960171862118567b742a63a9f327ac81b46278630a3cfb8ff830edf42a1f215eefeed980cfe2ad8d7bc7078622e8a20ba968befdd67025954de864760bfd576247570fbba7be073c081e3964bada2ff54339d9088e0b426f7a1396a8b6b1e861a67e033ad6c7fc2729cf4f00fb682bd868d8732a5125788;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd432e1eefad5373d2c2d067ab65200b1c5552432a8426cd33762c5cf4e27ef9d958cf694fb7835a5965fe2cf69abd5f7ebb9f8db839402d75efdc5bbd70efced57aa5093e0cd991a895fddb171e7cc8371bcd11a123d3e72fba42eda36f40f87d9ab0a8a3486ef787f235eb66c90da5382df805734aa5cc3f36fe6b02e7ca6e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23279b39acdb61e639319647e8e460299fb4e6c9caf4be78ec7e20a18614e5a51215cb62502e83f1cdc6b762ca7b0071a27dbd86f9f4349b28f2ddb33ad4416714b6fbf08319abec5787bf8f697f74a4e3fb4a3027aa3d2b3b0742c532a1aa936d52200466d170d23f85e78cddaeea6dc4b1517fc53fa4de533c9408946dab62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fd4c8756d3f7f7e6082278ef0aa4dc266133d3f87f7df25237e026a192e16eed4599dc806c521c7b0510c4b87a912979b78a40be51cefe03613ba498ce8f4bc2846d86e6850f1a14a290ab7877a1c096aa9a1f5001e39a300b40826b57ec2c9990b422f164aa16c5cb45ec6814167e8a656efe2ddc170f90c0ad81232d16aee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec00fbd2f1bdfbd93774c44efaefab9e670fac1668080dcc8b58622590a78aefa154fd05fd11fee4692647088d550a4733655e627c2e8b417be33554360d916e2284bd970122f73aa7176ecfdb60395de76ac20435402ff5eb09c1a7daf8b24214b6f00fbd82640be9f4bade7982bb40014cffe9143605e65c3845fa9dfbc3d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcca58685cc063ddd265a9d0f41dfc096b9577e19aec7003343f75b9a9d378adeccd7434887d73c85f342f9bf04a37e1c9c2306c93f489aa09b96f7d748204d4dfd870b869c719e3d571b4d3def583061eed03b914eef6dbae5de2f018a9e9da6271502fe422d52f35482aac56289c0287773b364474b1851be0f1faa610b863;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e683b76582fccdda7c5403746a2d4cf106727e0d7ab4b51b010ad574f14a75d41b1883692b503fabbb49290001ee82cdbeb8b1ffea222d464c654d41cff52482ab83366b1b5c873b0e79efa92ad0d96380c72b32dcf8a6b86e4bd3f413f030e4525d4103a47877b7d29b7e46f12ec34bea43be1eef2d5f7e7f69ebd71b5a93c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31141dbbf16169c6cb2ed1408b3b013d51a88ef412e622b086cbdf6c3e49dc493e296422c63846fb3aa1eeddf179a6e0fba516edd3afc82151f31e7c79dc93da4095aa804735a54a8c43e9aaa6ee6c5a5f4d5c313f2a0ba0d40b4a126bbf54f461217a7ff2a7f6aa5bf3d0082fff0609e9a748354849a628e4808e43fb13e811;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf52139769eb7cd016f0895992f511b0070f1f3c1d4e11f08afe398403c73a779d0740b53e379abac09d43678c96fab5ccf247b7919d90a5338fa8b7dcc92cc3f0ccd6b8e2475c9c0989ce80ac51a90e158294485f2290514a35abdefa6624978722ba1c6c6d69ee3a68ca3b52e9ca13d2bb291835b9c87f0a327ea9675aa8ed8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bd5983a59b953f9a2cb7c764b0db4f87ea5e75796ac87561026bd703414eaafd897ab19f6002e9a06dd8eb86e9c16ae2f78fcdb9047852ce5aee60f58abf303567c2fd89493dde6793e73e6f2d4506080f6bdb4ba965a44ab9827778cd7b5737a28ec03b9194b8f470f92bd01c5a4082ab2d41e1db61eb79c8f779d189cad4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h568dc86ac6e0f00a89f03f4e17d14c7369a4d10059bf1c30130accf626815e122649bfe076156a8cdf5ae0986f5a447cae05df61963bce9add8012ff0b5510494b67e4c6eb21f97ce4534f224cfb4d7a3dd36491a61294d7e9bccb9cfd949f1f5093006e6c942274d1db340d89a4fc45d82fe24167abed49a9a99d0c77f7c993;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecd49b3120416820d42f711fa6d0df86541363b9507460c1cf73a90eb7aef2e936518a9982b2be2f5ae6b3137c56d7ff4ddd4e38c0166b06ff46f930d71a12b368e6decb03e1d447572ca0ea6266dbb4f024f6c201d12953e9cc6aadea1b4dd0d167551b75fd2a8bee328ca8e52f19585d925ad90d2afa54948bd41ff44aa548;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7adbb96ce803049e9501c41661be3b7718546834d00ea427c6e12ffa2ff812793255356c89b3a21338c32410579662602ee6f0985241ca4578ae62a12a0185ab2c48fe875cdb18158bcfa9d55a2095214f8ff35bacd2c58a96f2e090fb5935bbd19536baa04c26b2a7dfe443aed2db2d76418c73b97e2e147c8e0674e020b1ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb071369a07ad7bec4d0e753e1a2472ec35c3008e4933b3f1e7bac1e24e3b96e7da1c47e7fc0b0b177cf3a49e6745b0a6c0983bce0fc9c87282a1b14a5539bdfe340ac4d12c0665b714720af9baa7dbf1120338c2ad42d317f99f5114a140c2dc0b0af822cc9d7f6be65a886aba85894351b8f71dca2ef22259333526db185380;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h359060f24590af9273dda6acfeb90434db8fb743a7bbf49bb04c9ea96e3f8be09b81b0468ca104db31d98edf8cf1b8e316a280e9ff4d9a012d310110b305bd0906b8634f835b7f45d692af097f0e91f8289e6c72a28474b4476394a069ead9ee492088c41a7221b3aaaf2f78538a48c9c7b849e93436ef2253d6bc7012427a7f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75856993079998677fbcd80dbf0eb92e3a2fac3858ba82f09d3d53325ac9da4b66a9787311eeeffc33a1aa484d5523a21f1f35cd1b2929cfe7df08026dc49614fdcdce584d5b84d06c295d7c37903d6c07bbcd705e2d33186912dda366bd02f71effa9e01d3c1ec23d117a49c298e2a1953d4c175820cc54f83b6a15561d20db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40267bbbe84f1dc7d33bd73582230afe37664ab1c41240536382c058dddbca6e2c1e76a001bae447462b2743c123ed654916638d320c17eca0446eee10b963f747bf147c1fcd3808eb5463fbe27629a7c2bb70a9f0e079890caa48668c3a3bc4d39a20d8721731c92b4bcd95fc7a885861cbb734525b974752651990fe287615;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f211fb401814ad94aac044def295c0fdad1bfc64691a97f4931467201ff3877061b6fce09c8107a43986b1472a768aea078a2f7d22a992b8003e6d4a1b3bc5347a3cb152b5fd723379eb4b430a8fc24cd809b76414633613608a44b00273afa2404d1921d0d7fa1967acfcadd836c9ff7461f36bd9371ac4cfd59cccabdc00d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9f9f103319cd935ae04b0ed52543c71b727a7c5fefc50e895a36f340df1892d4fff877707dce4a44fa6bee804aeb2fcec501d700642f90bef9f446ed9becad0c66f5a110ce39280f8131e362b6aa20e918eb26e5e80b25c6dc2a352dab3d283729475c60d37043ec762dc97716aeaa5303f09263ae2f80bf116ef859a7c611c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h597a7f447968e7b4f64429ffc3beb99fe81980b64e78a6d6064956ea2955b3098b4847e39cd0b5cd4c8ff48954dcf83a6d2ab7fe918583c78f118055613184ad4bd65956e7d43c907bda0a1408dca51176dcd53fd0dd810238021d71aeff711e3b583aac3f17ed3756935416455978171940b522e124b1c4932e4b4d3d1a8696;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h426380defcd5f110bef79222e48263103ed55446ca77623d0fc6473935d01e6fbb3b35a52d20a96e52f7051babfc85b172b586503c59f5dbedf480e9018534f372e553b8d2179eb9e304dd1cbd91199bbccdf36454e7dcfc77cba7934b15a4002ac7682f15eb9f25a2b745d823b68bb0a21cfbe358abc517b8a678c70cddd660;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53425a60ad377a87aa4ce3e5ecc38dd1c6d2049b942814030cba37485fa1725f47cb713497db7d62d60912ab6a445c05afe4e38fa9e054a86c86bb60749680a1b7d502a021f52af772350ec82da48491af4653ccc4fbe134982eaa0614867eec74e5a56a25ff3f1d1df904a6c11fb39a814146caf85753fca994d94853d96ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d98efb800c251301cfa53f140a334649e8aca925cdb8d16b54a876ca27340fdbf2baac6bb1d6ba54fa6b70002fce21bd11d3c24a7ba5432c2b61046865695bb1056d5e6de61b58e5b437b90ced05fa8e3fe61a29250272bb99c45aa09c22bed45d6ccb791eb6421a635b579d0b6979f7a92145df2cca82aa0b8dba2156f3221;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4dbfb5a53d144410be232d3a687fe0dc38e5938a1e4f6b0593ef3f83f3880f13827a824a79da71cfb3b82304d4b556f64665c59a5301a39049a599410391a5e3bcaed2467ae9279056bba42cc2c495eca5aa56d6085b0b5589af74e540f1b02764c24562b158ebe766c150c3d0be35eade58aa048783a61074dc1820ab04991a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14e80b19adabbd79944a1a4bc4d7480114fc9edcc559a7b93156695ef0b4e682d6b6166171ef3db8715cfdb5f6ea3d89196226373a875cd9196346ecdc7c3b1247c493403542daeae68ecd16bb1ca1b59efa445d59efebe82afbfdbb6ae4f3a460e518a8422dcaf49619aa9341b622ee8725a3b5488168e93bcc7165579b3fd4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h343975d129c7b96ab5ac42bc53f8959ef9f7717b99ef5f3e8d12b1ca205fc27a53952e439c4a38ed5466060c0e4927d94da38b94b2e087bc95ab5076cd74c928b26b6324b6ab7384976d38d006dec421362385b2ed1d30fc714832a4293cdc9277ae92d87eb8b8c75800caf95bee25faa4c7d811b40b9e8c26e61179c76f62b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6906089cb4959b86cc467a0021df192dd10e35e4d5e2c4e202d6a72cb02c8344045256be71e931feefd5bf2c811f5eb53c7e6d778e616497745b8fecd4c72c68c7232552e33675b778108be934eb07682e001c2edbc935c0e3b7057c18d4aafc367e7b36386288cd1bf0aeadbfd9a6529265ec646154d0f4f93629ad64d4b1b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed819ea5783869b0d1ff4efb9f2b646638bf13b3eda1f724c35c92902651ad4639316ac99f6698c8552f28faf870062f0bc96cae27c73f5e1eea99a60ba8638dddd51b41c870ac54a3774ccfa324d0514332251babf8fec9d4ef1a87912efcd75722545c86687352572befc6e3aabe6ff637fba8459a58abb83515e16b57acc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b35e1a284590a5b6293ff80556c4cf411b1fb93b07588d5e0a9674ee484c93262bb5d7965c3a01a65820010f9d6184170925d28cfe06fed724e8afc0403932710d76f1c80003cb8675c2d568f3baa92dc50a86363f3cd9acae75b4386f4943a81a570cc2b752a00544138f86f1439b0caaba7827eb412a9126d1ae19b2624c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e4b1e57818517bec5e3f7d201b00e87fccc1eb5bc5d7ae6bbedec1129b1d6fef243dd6b71b4fd0aba55fc47640c69e215f69d813ba09e0ae6dba187de73940135170814c0bdef5c63638632601c05de205081a39c23ba1b839c58fbffb66b2f7f20c378dfce8799b711a2ddb7d3c7cc1fae8f4798af93ad234c46496fa5f782;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c6e6d6a94aafe63e00526c9f34689909d7107779a2d26a2a0f6402d29105239bc42d3bcebf01f49d4b561773a55140d143e2c4ccfbf7aece110ffa32bccd650090c78bdb9113a37f81ea3987439448037fe2ac5a6c45f9fa5238fb3f4fc4b256ad9117ed1e30c69f2eb678e71282c7084e265499b9889b2dd9d216fb0b3ceec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5106f24703f754d162d781ce4d6b42d022daac326a829d3d1c0b4b023b40f54b5c2e91fa1eb5d2904a70d40747de375637d5e6f827be82eb90bfa7773f547848a1a2104eb2ec0861e1ec2c091cad7853120d3409bc0d5600a9e93d072a6631965873e0c0bef555064f161973573e910158d9fdc952ea6933d5c8101ee7e14043;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb3fe5ed1ab81b122c0edb0fa682aeb6335399e5767d1880344c09767bb20b1c86b2723e6217c53e61ad6786c01b5185dd4fa98b112a35cb686c5060b67626373f32afe273d98190eb63c0b6c6c8bbd2f41dc3ff57cdc232f617205a55516878ea4b9f3efb6ad7f1c2d2ae0b653ac6656ebddeeee3547b1746c76abbf6a92251;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb41a89151a7c79c1bca168608c0ef1d3973a12caa5b77efe9f02d7305060cda395201a8caaeed6f28d22e50737897e19424058aaf47d30d18f16a347020284fb6456e4e17bca2bf1a95bcbb06b5756fb7c162b79be719a555ea4bb374b6cc0a49e78367fb756c6a37ac6e37233257c78e3e169939b4e896a5712c0ef618b314;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb0c0e248950513b2506d577e60790653ddf9f9e7e1cfe4e2221a8e5fbba7a35f94d0b490d5f0480d49d0f726e86f2029d3f6e4c8e781343dd5b6b7d53fc22be4f5613618860de27b90464fce87614b11575e7f2d474263386c4cb34f946a9afb2ecb7f9f4e5f11e9cff1b065436a790a718734fa99ac2885cd8eec88a1b0b3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd158db767372c9b436d67f00d3906b67ddb5ddcabdb841d69bfc81e967833934a153612778b05bfe0637ab0ca61d2d234ce3a8172c6486e273745473230c2119a86afbe7cf1cdf99edb1a8ea6a2abbfe67004509e4adeda59aeea7a9341f7e8e16a1573b60903b2cd4a694522a3da58694c69f761b8eaae92f25cf60775d3b1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed511dff281c2e9720ca12a1bd5e8c0ea2a2c9553d4a05bd45010a1a6a93786b9baba760e08ed386b2b2d88dccae5aa50b02a3b0d92299fedb7c82a2867c69e19f7157a16edfdfb9c3c081eaef69e179b653b546171d5a7b3826f31a9991f013d12539151a73e386175486d85b09ae755d266148b2b03c0e7fd2747011ed3b60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1097c625d172267153edfcc5b0d6a7bb4b9bcc2d0c87def50f1013bc2d1a5c668010e3b724a6e83116a7ebf091d487f8a4a416944e29ea466b90cf13ecb45ec3328b0466e8c20803ba0b376a55db600c1c6f1441793e31668df128f7b4875f16c25738981c0a2acc750534b26acbd25d5e45d94e13e34d74dcface714a95f0bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0c4ff70911cc4c737ab26d8e1ace4d27bde3c7543dd0bb047efa89bb3bdb99048aa89cea03565445a4a6871f615d798173135cb4d9c8a8fc65146fcd72b115ef71822de13732c9fab385771592f7e5667e2eba4172c7aecee458aab5b9d3876926f7149cb4a4c153ea862ff3eb3b38d6e370b46a3009e34e91038f33d6a594f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f2c2efd997387a4fe8e4daad7124e3c38c09f794422f31774b141aa47f0d6e97051ed9b7bc4b0af00a19307a7d46330b6c20ef774377929a5bc5c26cce96a2097f462403540f01ee8148233d84681ee835eb63b83ab07178f258a48aeab8dc44f9f959560e7e01d86d02b546de4f976837749742c3d70f25d484ab866a78151;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93fd491d070158424cbf99cf435c7603ccd965926e2b12c804d3507d1715fc30f6bc940e8886e19875bd9fa6c46ea247fce6837c185984205bd33aa33e2fe607a2b706db8c13d9a94011dd161a215ae5a1fbdd19c93ba4d7eb1699636ef505491fd4d5898560c95731aec3ee4f5fdb1febb57184db0d8a803841b88dba17faba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7a466b83ae7d4fdf585e4a36a5940f66d4a9f9cc9f351bace288f640d3aef77ebbcb971e0010eee89250c226a91e4815b43ea23f5a81b2b69eae284922604857223c602b9f7cb0aee0cc53edaced8111031e77718fbfc69a8f462533ddb3cffd681a5ef01c32e00ef1109810918add621c0562dd74283c3cdc074b74520493c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha77ee302988541eed6b08bc005d38f657e378528476be811bdc21e6d094fce3f2c6cec12876cc4ef1346ff3afb2aecc4641c82de41f45522e8ab15cdea9c835dc21ee9b3486cf11211b72a77ab9362b7dd587e88912bc573a6c3f22131a582fa5c73511b2c990752cc88da85943c1e2932e9e54ad7b5634b546552a780e938be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61526d5a4cb327a554c8f3d484e78e4ce64e9d035edc458c367bbf3880b3e400f587c28647fd082f674c801b836c9fcf8f3771a11f0e735373bd9fd747128b2d5bcbd1267942a741d6442c81d6c30b5b01d9e83d78f7f35ce68f4aba80dfe5c730e4516522783a7eedee2025e760184348eb1d9df4379ff59605703aa5b249d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ea4b0ae3c396e3c929a45409e19527326e0fcf5b613adb6ecf16403b1fe18262021bb77d391d673f7c6cfae16a4b9e62f94e1dcabcf4ce7f640c632c78a9df7c001cac7fa8061c27cede8420a64db0e55292c89400a45ed2fa158f87c235ae15a7db42c19a3f9df20cf02e2c71a46d1d35fdf5931d15184bcb03fbfea18b664;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ef26748f12116aa453a2d4ee1f598595fabb757d20798ae3a0d2fdd64e51778fdf4b9f92a0ca3575f09d658e9bd633b6661b41208d46c940ffac53a30a3c90e885307fdd864954aaaef8717327a441854971c14d7cb5762833a4415da18c2ada63598a1f4cd6e3c0ae6237a584edd28e73291aa4f6ded899fa97083ad2d53a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e10083532476937c96e13ed4bb40599fd8f4284a5276eea2eb0903a43bba51c9f337afd5038881f3e0e3320d53d9df84f2acff2e02831412753d8cd9ddeae123fca011b73f1af8a08b9e56ce20b48adf04a210f70796b8a9b04a67c299757bcb9de5b1d46f1358ce7223f778ce37706705db20ee26b8eb25d858ab3941a576b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc30be977fafefe8ee3da7149c688b11edf103f96afc7d8f4ba8644b32e4b9745b888f24d3008ea6d65caceb19fda921967f3d6799c3568c6e6c3590554079f32147c163c8efd22963a869409fb11edd077ae7fcbbb43711c05d10f9644a529178d2d844a4629a3fac457ab08f124e5c169def639d604110e13a8da8d7076536;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66f890c37bec5063abcf7b6ad47afed22906937616ab3b3e8014544871bcc597ef6354f2163ab539925e1d031f4b7390e294b3d5e6ced64fccf38479122ed21f102b01406959f1f5025b2a13a672c04d025feb92108bd962cb5cae433d43bb5ffc0c8ec78414bb8252f6571782b90428394ba94d3976108e850b39b6b1e2546f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90069cec2fe8aa092b77a425f1b6c4448a315aabc3f20297e738dc7a257dff66bbf6f9547121140afd074f34fe032e1a64ee327d0f31ec9f19599a9e2c9476d13ae1d49f7f160d1fc3e68368747574f5b7c9b2ddb96b7f78efafac12e6aa3e949fa1ceaf6cb03386d56bb73d61b93901a449c7088afb50414efa49e796c01d79;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h448141182475e47198b3f8a03724a6ba390b9380383ebb5c28acb0e40236a106ae4082742638510ff1dcaf1267bbad8afd7ea523570f9ba4201620c07f2c08b713049240052d2a350ebf51218af221bdb0b36485f2bdcbff8427ebac9aa7bf4f8aa4f81455446602387b8b6fc5e068bcc05f363e20e7b5568694408498974074;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cebbb7d5df0b9ff8fbce6f82064006c808305e4f957b92f8c96f3cd0ac989639a31dc288cbf8ad40e0cb6e17039fc7b3c4d84bc3302b6d0487e3cc0197099c79faa24b12edd2595a5226ed8e1ddd1de4df77726bdff413b230a9b007aea7982fdd0e911d779e7580e5b14723895a0a4ebb3d7a00cb60d45feb559546a344bf6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8506f6555dd36f59408242d9b12dcce1d328d3df86d9c79377e8ea4e125c5b5d047552fa3ad4b4ec55e5bfaee680521d08dd1d5d264e3f6f31f1ab03d8722389937450027ad9c9bcf1961733752eaf38fd438bb0eebe5ab603c44c8a2b70120c961abdcd49fd445b7d9e5f26ae67bb038cb9d63009dbe4b43516d1353a33dd92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6dcd7367477a552447a38d34c5cd09972fad144b46b72792d7f1962bfdfbc2b75fa0b85049554c174aab802e2da8d9d1565f7eabc91a008f8aae72166dfda3c9f4c210190d49f9505613b18df7efc23c844ba8a7b42f5707f89bcf89dea170378496d70bf0ac15b1dda0b0d3594da0500e046e4094a71d2b1a078d6ffad315a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c4c46f92772fd88482b6db48e43ebe757197fb610102ef772616529b4d6c27c2fa7061435729ded5f6acaa632122d844e285b93663a354b1cee29b56c7caec165477a56a09a496c520cec4350b9238582fe105431ff944d5322ae4233e01b98c46cbb6c53ee5427dfec3598dcea8d4dfe0a5de9f1246055fd9e1f287ed125ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d86ea0a6e2c7681d59a2afa2bebe8eb991716f6e61d24ee8b2c1e75f02e2579ee7b4b152260967d19a03ec779b5d7a73293bcf5023011a9d8f87caa4b6babb16fc5b94a329b9c3b2e7d1379cc98745e91a5b88a958a1fc2a189055ce07b29c17cf7fc38bdc1145de112b3da3fb060cbecca3cb07db0bb1c35f18fcf9ff3a30b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb3b1b246afaf6d4b79b1bdb8bcc33ee2ca108348722bb0d39c27344e4d802daa395be7ac9ae1305d34886ae4afb4ad4d5ca0394140ae7ffed95384a44b580ad0adb4e6fb139aa5f57cdee49aa053320181ec9e0fc7fb4b8b5e3f33a0b48bd99f0e8d94ec968faed820b76488fbaae75e51d457117289306b9a6e1ceb7539207;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ae60219455691d2954a73694ffea3c69c21e3b05643a094aa7405374cedfffe2562f0b08f9e77dd64bd2bc2b75a617da41ca0cb0e6bcba089d423d922d38e77c787e7b29ab1afbcb70f02989bf7313e412ac49f10e54a8342d82432a97aa789b944ed638fb16eac8cbe0ca6cb107b75fe8b2ee20b5daa6e955a5ba72c0850bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b52bc8f8807f1c391abe09943d5d2f2cb270352d1dee8b0e127e79043ab3505c338268ad7906dc0ae055bb70fddd0a308c28cd08151ab586ccf7094246390adac57b37a8a37ec42e73922a8e53f03bf4326579736c208d3acbe24328d2e5bb10ac94ecc54f4e53a31d7b10c2d93ab433becaa903a4c4aea3a19a57b694ce99c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he47e148f7de03c13045bc4c62c90722b14823325049dd223ed65879be46067e1578590234ae847b2e6c4cb6326d738b52bf8340bba8a8b8458ab0f4376f891baba0ed24f8a7033adf2ddea8844f953d571a484f28377d4e0d81066175d96f833d4d5ea923d45cae2850fa74ce0011fa8108a441e2e384c17786352988d6448e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h291a329347055d3cc3d0d833f1c214bd2488a493d749efba83eb71d6f25d0d8b2b95509ff301c22c1ac96ce8e72816194d42522f903324d4ed2dc9ad742d6b16ac195213e81d978a9a47c7264ed33c056c5076c2521863cbc393fa92945aa1812ef0ef4c5fad1c55c9ce7a3c3fd5f09baa0d0f4dafecfc2486a4d47cd204852f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c699c82c0b33ca085a07ea890144c13804e565393939489c54210786f6062cf5ef88d3a290151969dbe547fb8d2a2d8d082a4e42f2c27c702bdd2a2597c4752fb8f1d4f433e00f217ae886bbacdcb0db0d770816c19ecb9f46e9f69280c8e7ba01605cad462cb9daafdd51002fa3ae871dae7038717c5f53c2f464d5538d5cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h858e64858e98e5c0d1fc3f3945076da478d901010a8e959553769ca64493f19714bbc2baee7206e78d92183019e7b197d7cab36a6f0c5f619348d90f3148ab50918a875898d880e456e38437b8df5c5131f5a56344c85f5429dc53a171ca94be58949dee14b5843cbd9511bbedc588dc365c2f58a3e3de7ed2d9bbc95101abe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f4ea23c8d1683ccb9e546924fa2fb9c07a909cebdad5925189abc73c7f1aca3ab8c244f9498af884cdc0ea1d1b595b605a68c74f35a673b0da3f69ddd717a07890c52ad48cc072053ae968129d96f82acd797401d562fde3b69ddb375f697f5f1505588951816fea27554a96ee24e75f8f647ffb9646081e3036fb926236403;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7de3b570dc046697a893e057a84cf13d0d0aaa1ab41b0bdd2b421f385a2802bb8ae0b70dee2b6a2f4a37e9480d68db9596bdf7fd30d514a19bc380eef0293d88324a0b4a9c6479a1f283c5ec6afc748dddd391b45e8b3061a3c0e5e016b5eb2194652d8699996ee84c1f1adcd67bb6b2d491f31ff577ebf00ec8322d054c0626;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0d2351fa3914477ec3d5da43839c08277409c3d7660b25819d2337acd4d8e0d5329f6138b87647859a3049f412eec2ccaa2c5e0b53220a8f3928f2aed4a23db33e8a51fb4b2b5bb01710752b4a40d18beb604d58dfefe4cb074c127679d83e59ed878faf966fcb67472b1388d43af4eb3cc91fe880efd19e8a3e5c8e2695c9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b65c69940f34166d4c9fbc07ea51a43d8e7f6fe890fa571223b6b48ebd3fa808ce7fef9a28531217f629689359c667760454de72d499a30e602a08ee472298dfab1676b7797fe8546db62489f11662da6a95d72ecb5123adb6ae5c5781f2af3f898661b68e13b76419a4181914b73bfe85f9d4ce74c51048cdf53eb5ad1426d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab8b0e63b3b54de9aa69d0fa2b3a706ddfbefa0acd502eeaee920f6ec8c729dc50756148402f497388d8593b0e14dc836775964a6e67ba6706604fc69f2496e527d1719fc456ad0795577f588197a07dc30d17a56e3b66d810cbfc0488d5ed7f829df048ff32627e5000bbde91c4ca001b5eb5f7788a0f6fd9d5481b34d4a283;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8bb89079ab00469f96aa32763e93daeff73581d495b2a79ea68628092a67c04e6a816663a70212c2c4c537d47d5e2bd20e2b2d05876b050dd4cf3ebe7e05f21b0967be918ed8c4a60cd75c90c2d5498a63d3f2ec0b3b794bbd09bd55a823bb531aae576e3a3c6a11db90df11abcc539a6a1d7867d80457e3b7368b5a4ec504b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd708e5c91ced9067d270238e3a622f0db82e08786dee2a2668024360eac670b085a6ed707d57932b8e52b3266a9ade59592ddf004f8525d6b347f05c253fdc04ac3b898db8ff29c9d980d039df2436a083e4be23812eb2a375c04fedb08ee179c467d06cad30ca1a7a36bcbc67aadb6f5bc511a2c9f566cd03ae5afb7b03cc80;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74e61755c1a47bca27ac02a55cd149a6b600ca4da2a0db992fa1f7ae06c59465b98eb3ae1433d155dbfffe5be3ccd55a1d458f087bcbc18007c2abf5c9e6ea5ea2d52674706a6fa45e3504dd18dfddd3c09d31e63cd1191f8c726ffd0e790af4aa3abcec4329351dcc2a587743120aae72fb574659bbe5669f5e601d5e9f67fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27ebf49bcf4700f85f326d815204326ed7e509cadc5ff17991b92d3a748174243b71ee72884776fd58ae0812696e0b157f0223f00fd9800cd2a16897fb8a6591bd15f77d418acc263d6a3dd0ad2a71c9df79014ef2dc68e4063c4c57483de785728eba9c1c9e2b1744bf635610d476d7e596814a21a005212d01b2874b411ed5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h990f3bd25e931549a73d3d9a42129849d7414ee40e10128f91f90a1d0280ee9d23e285f412f8c7da0899e8e35a4007a71f15c0ea74799b2e017613aa7cecf454f82c5e6cfeff31af7a8ebcfe97613946ca523ead0f4b8a6bc7a12aa04306e3d0ca847be8aceef6db1aced2c2b6fd138742a2443d84ffcd4f254a324ff8f30d46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0f6aea8373455683a77ff916ebffb3871d3a0d3437377889b56dd751a5fdee36e3589c2ad33bcf584282aa563c7b1a5a83de113e24273cc8fe62257306be05ee7ee319acf08013d323742b2bd11fba78d257d315161565287bc38f1b5c42807d37e6e1b282ebc3be4cefbf9555cef0d75fa919a866b0654cad88688e351e9f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94a19af068debf0273f1af7fab8b6b4942f11ec9c2eef7e3d9f88dd9369b9040406e6e336361832263f829f4cfde17d0415bf219a348c87b34dc2387700c5cd1b849c497cc9371a517037ef75f56c5bad44b432f6bc5734ebcb790c1b9ede0e8bda78780426796f4c754f2bcb570500bf07749cf241748c6a11b396d95fd4915;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h619f7df25c2c0bce50b3b08d3c4b1d429213105cebc753eb1e87d9fc5de901092cdbbf1e7d3a46f18ea3cb97786abdbafa6f3aabf4c297f6116af33076e9dcc95929640c3c8b86680ae1ec298b4c59f72c5a14a8d9e8eca29301cf4379cea046d99203575eb397b2796aaccc9b984c2c706538b7b5e454d08a11cfe3fccd9da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e6acd398f94e94194543e2c529e7112624dae6c84fe45f03675d202da6988a0db439532cb030b47df611c6d0c70c3010fb84e5da1738f2ce3064e9162f54f64343b8c900a7f9d831981968f2dfed73907907f6c9080d69e882db5ea7f84307853181d57358a9915e771b9221057c8311a98545ddf816cd35f29b12f3b39f8e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7dec395f0e3cb75a6805ed8acce67524ef33cb9b2964e626c191ef8e76c4875793ddd68c5cb4d5a66caf0de410eade43fe0d99cf7430549216f255e3f8b468a52024ba2a990b06e6cbf6964c1e4311f0e6125333c19d508ccbde400fc6f1c4b2a7a507aa0d4cf55422250261d547c0c027197a03c8f3e9ac61e2bc94a912f31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h636e5be30256d55007b6e84d7ba51a25d40cfbe0ed3d88bd2223ca5bef8964b8ee349b97f4577083a2c86184d66c02e1f1909862b163a802ad332e1b52148c7efb2f22c948b074c75a29aed60f8b27b00180b731da7a7e05ff92751a8d38bb137b4d4c40dcf9d146e543f3a01b568deacbee8d67232c38f34450c6ec711dc544;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57a1e8436c953c7bf12ba12e5ab600e70205e87661ab9fe6edff7cd0651b789761a0e366889f99bf18d59034fe2a6e85b27617aef75b2b5fc679d4f058a97eda058dd9cbcee125a359cc262228d105c745a010fc1b3cea4e62622bd7c7ffb16c5715a88e403c8e7cfb10f9b33f849e44cce5079698cfc126c7a0508c6fea0587;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd415c2306518a127b36615e28e43a74d5d995896406a9b1bf50dd70d283f3515bc0fe2c4fe4f522ac07224e9dcc16cc2a37ce6660f00507115ce8c1d8717059c29e9e3fd0d77192d371b85a6259e5f92c44dce6215ffc246c95afaf934873657f955b18692200c97e58d57cc84ffea2b1025388ff54425f313249b757defb374;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6887d65e5827873378f14311e7582121531d60409a4bfdd51746a3cf6ab344ec015d2ac03fd1761cf9ec7ef02acf8fe07dc6832d59220b55be87851ddbcc63c31c92e187d7f376942b7a3089c7118935c4f73057be307aa524e2748628ff2c099449c1aa5713ee461b37f80043732990b01171df22c3ac881cc7abfc406f335b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf09f47dfb92035ddfe09215fc5ec52a1013175fae99acd099c1db6c8d3a06a6a7b6d0737727f1ec69b7b0badd51bb4b7b8528bd54b5ac06fbfbff3347a43dfda1194623c4fc9490dddc55428e5d8827b1e7fd712414fa66851287935608ef64c4e57b62e9743854bed6ddea4beb97f34b487930247a739ed620e0debcfd899ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87ef128966b14e5125b64ce5c8dc5c76579b3ac508b8d9cc5f395b22f224f8b97896709214e772a0bedb7e4bf41e847aad852d74675a3aa7b4f07c7dfa3b4aa122d5220a1df0cbf8b063a414149b761d61c7a90804b957ff0a29ed1d9e59b0784213637e0defb0a8e1a692519b1f92bd975d8f947bf6efb12b8b837f723c3cca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58a21b78c8bd7ba35be1a93bdf8bab076c5fc724be93ce2a17dd9877ece9981521edb9fcffc6433627e26e0b163036f01af505fac8268821670cf7a51ac1b2309c0505b02138333acdfaf080230181a5615bdc37419256ac57452fdb25b68e4dd45a6ecbf3a75d66f092b0abf836546bc4753195c568278a6352b299d77ed4c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h239e5ece1801d6ef04923f7ec5db797757406350715d3413a9151f6bd68d18f3bea2acc843077b1ee6f9c12fdc4d96920542da155dcdcf208d4535cd89eb0b2a2d1a58a8319e76ff1b3ba1b3ada68d750e62db76d363e9d91652c5d0c3c757ccc273ff8b131209dcb00db9e553f897c84a376fe0be599f8e53b516e6f23193f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40d1904c2c636d2b6fa08511975245c6eb8b51e6894fbc22859b1040486480cfb72ac7714dbfbda706da2007beb159d2fbc6dff75c2c6d1ee2aed10b283b4c0a9572d30d7bca3484cf2c61a3261cf8053ba0e9ca5c7707d508e9e90a22047e93cbfbe469aea5cf3896fe22b1e6cb2ac609ebae312c04e3b0d07811b6cea0b4ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c488e113e88614248aad9fc16ae9376a896486984b58536a1f2c700d69cfb2bb34742cc05aa6381503584b54434b7b400d0be6789550ee9ae7d69ff9902629a27f94bdaed1481afc96abfc1d2265f056b5d278f8e3ada372df521cc3cb6162d1dcb7c35d9ad124c4cf3e5cd982eabb97c8d6f173f883cf32f589f530966b0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8b34112b48a8959f02573ce21f4810f92aa25fdeb645fbf35e206cd37cd5ea0617e85fdb4b434cc5ba2cb5c7227ab2b19e6af0ad1f228496037c8503213880f8ad26f952d72922a5616b500e98a86af61b11b4a8eb5b7f96fa0b11993fc30f084d41ddb6eca3d94eed449ae681673c6edbd241ca830cfd5990fd4feefbf6680;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde3c50093a4aeebda7c9ee80fc4e0d445229b34988865faa7c147e551154350928eac4fbb095dfb687d8a0a131f4c1acf8f8ef9f850e7d22891fa02baf22bd606a9e574e1467e95fe468072082bd41f1f8e49f2efefddce2bbd26f3adcc8a9ef1837464f9dfbde04698ed0e21c23bbed451a461e73b3183e37dd6454c4f5eac5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a56f5715f90f56ae780aa1be6745de9abd39b73a0c96af75101e5f3d16b6cccb5fe5d930f05736be2e3a2ab2d2649a7c01eb63c3abfc9ba9e376d31bdf2e0557f1fc4d6cac02f5405ed0f617cc14cd87ea9f1604a92bc5c5e9cf33f5bc2366c6022c0e3c35bfcd01524da37e55ba034e64968283ba94e9c642742f7ef44744d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h900b2ccb1c6bb32a228f93895d9cb706344d84ba0dd119718738fe58f5726616e1ac5df237bee2bc3f1aaf669069a3c88416c12d658900ff379b75a4c5ea9a8b7fbeffacb7a447959179bc4c4563b2d2acf44625945e4ab5e447c643e00db23f34c78a2790f6af28587eabe443df465462da5c0747de62172d79010accaadc13;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5bf0b5f31d10e2054ea5af6960ae6e2c0c4daf232841dbcef697044ae559849422945387b23d342c87615702039cf4facae303117af1cee277d1904bcf370500d987cb11005030c4d4196456a93542684c5d4ef20e7b0ff855b878f2ce71bed69099f7538336b7bdbbe9746a6f0b6f4345595abc6f2e817898aa4772448f83c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb56765d36f4b6c68ff9d88ad0c0695544eec5b9522ef7efc5b365c7cf88c629bce2312e886a1fc56f4b26fbb5699e2dece315664151b40334a162914e7574d3176432656eb071cac3b9f475b3d9b30131c8ce22ae57f33e637d89e9c6248e13f41ebdb30df4c0ddd93bc664e6612504b826761cb7a732dbd6d315af2c9593da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3eddee338d16d7e767086dd03f83908adc90a6c1609fc3a66332b46f97bf2daff2eb7fa0ff6b8b97cbd1a5ba02fc013804749ec04090073bdb61aa5f6016059834ed393adb477efa8b564aaeb837e01b3d9bebe6daa5ad1edee2a2d8e3f33707c3bbbe22778a1a1fb536560cb324e5dfb0a17bd413ea971c153ea828fe44ee4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54633b4548ca6f2ac05e764a93f0dcbd0fcb6c9986ee9b7cd756f206ebc340bb03ab6d2a772487c108cc5bda50cfd9e812a549b5504576104b74ac3c2d56463d79ce0716b9f51960576cbdcbe7ad302141ce559c01ec9a63ce4228893cb821445f02988b9b92c804af3fcb214d89723cf103f640b4732519008f8c7a09cc5e76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b50a0262b9aef9f78d1ff05a3e44d6b996b1377cee6d476ed256aab642955293242b35e9d94ee59c37f2160385943c9c4a60b2adfa080eafc2a048e983117396dc5535ce8537428700a68f79a230395412138e60dd6a25346896f8b31deede4ff998063f201ee1293bfba0c88ec59bed00e6e3a13c0c7d1ba6285778adddd91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedf2bb4a7bbb8d85c2980e23de6508ed1da0b1a2617c9e593e5de5c0fd69c1d63443cf242c92a8518515552bf0315e25de8d6f24e111c37e36c7628be35790c354f619f0b5914fdf20dffdd81399ca255eda006720d802f6a65d9e83dff244e3946ec4c839f7dfd5a01cadcd030460bf30fa1bdda444afdf9f09cdce2ddecb9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b6b4562fd7878839b3971eff17eb247a05912b1538bf80ff1a06233715d39f6658f67128b3f5c06d957617bcaad0c0d683ff87d484047d6053b1547258a6a94ca590e0cb83a382f1bb2a67d47e17e673d90a6d1150464fd240b6b815a0b2b5561337097b7b36a924a9665a7ca2a01d4db582441150d61e9c8e95e9ce1315bd0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haef494fa5f3cd2504624f2882121d27d544c10b073bfed32bd432f7f4e70b56fea013fcdd3b1cdbff2114727efd18443bd896c02d00f411c5c5d7613e5fa6304e2627dfef00841588c8d415fd603b3f11d0c9db743b9657bf7aeab0bec90337a9b69aea97eb8213f5b5fc32d65be99da92c303c79c5f9b4b1983d15cc230e7d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a5c1fcca1f6334ebbfc3ab83c375cdda975e0625304a709f4e978d62869455070861ecf4abef41b57cfadd4dc8dcf82ea544092c2ae607d2ea3157bec82e7de4cc5c8d2b024c9fa0fed4aba6c8808667193b3ddfc9c14ca713bcd8e85783db7fd410cc86495f3ec202ef58121ffa731fb0402e68a95a8c60feaf566553164a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ed996b8a657f8898419f23356311366bbf67b56413060fa07637e75634ffa51addb4bc8dd83ab32d753a894b1f3475b45fd0d823f4539f15f998919a0ede4e206ba98b9aea5dc51677c3f5cc31f4c4c57d854101ea22792765592c3b054b627dc77778e0ffca39b1a01ebb2a3d843f55ce900b86dae41ba345ff70467385cca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9cd3995a87367fe1695e53b92c01879c5e6682a2b58ba149d9742abf8afb1535d4c0a4640a77a325a09d6530a6ee720a4b730e5914a7c4237507d18cd47fdec167da882c9f2648b023088ffbf9aa933e49f98efb4b9fb87cb243103b327e7684adef88fd76627d2cbd666067f71bd78c282d5ec83c418ae74ca7a31e51edeeb3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h706ca3a228bea18fc9c07e4ace297fa7c25239484ee5a699c6e129c68f0ce7939ce1cc3fdc78d062e6b553a2ff6fd65649d04b9915e8609bc5880f9568743d27d0575022cb2c60bfe9245fab4fa10ebaa562a769bd1965233f5d5f2a7b1e40a4688ed124ff63ffcb24c9cda73268cae7dd0386b3a78709514ac018aeb6076b3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19230a45c4a49d4c2973c2e6f265871b62c279027e28e241ec5564620518ced6812121e0624aaec67dea1875a1ea1028f6812f8c34cdd6e696705fd519cbeb10e890cb184ae688d0cc9580e51ec0755cb217d2db7f3486ad345dde262025575214a9557c57af37e72abe8785d20350f9a517ff27106e9a9023f53cc271c3ba15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f7a78a46a3d4273decee67d874777817b50384e62400da758696ec285f25369a7198b444ff22bccee6761855ce812bad646c4a5fcfed629590849bfddaa6d5c306cfbe2535aeb5a8fbba358a175c4795b1ac4b6c7c7df576681a8c77537690ac40fe7c5562f0dfecd629ce3cf28a89babd722c47d046a032c26b71d40031498;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1298764c09ab3ad5f04ef9f475caad54f8275d29c85a677111811ef71808e3ce869df9b8b17bc912dc787a7450adba18ce875b9bd48b4457419a49d461f03625fa78be88bfb0a4d473aa4a9b80a0542cdcbf95fcfbccb6d6363b1471d549226f82dfeebd7a37651caa8ee40569657b47a93435b84501aa5487f43873a8358aca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73d8275daec199b37e5297f7ea5a76481fce6acf119e3b06374bd3e28dc7d496f3a6fd8ce10d1e7a106d3e1d0d56bd87e69b7b3f1c9b2d0d966fc480d8a9c2a36d6d03d6fbed32d0aa2412613e4e0b164039fb18ba4f58f287a729d00f78f2e5c01884e1fa31958096b448578f49efb3750ac032da8ab46d64444a9846b68d61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8200d344aadeef23c16e2a377ef4c5a58b8d91b699a9f43f33fa93dfd3a517e57dccea9aa58804d9aa9fc4dd513f5d60d6fe9858ebf37dafd49b2f4a4bd4704252b680f2d69d99a24849688ca348ff08f13a3d60d809e1b9ed7397ffe93aa90ae9b502a0100ae4c885439e027fc14592accfe28f111643581a35e3749ff97ad3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5fe124ffb1fa24187683d6f8f5727a78ce6db7dcb3787b3d2910237c053c9275e02f52af2d377aba5d7f618fad531d3779298c89221f39403c6de40ab0461226d8236990a0c10645864b35a919c008014d44adb26d73ee0c6d7399c5ba725103ecde5d76a5bcab7990feabef4efcddcf02e8646d0074988b173ae52b251168f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf23d6c4347a0d2dfec87bbb4569eee8e5f898b3c2a29b0b2d1d52b7875894c8e69f39603c77f4ff06369aed97f059a5cbcb5893625d9c7bce6eaacc7f217bd0b05c5221065d4884108779b37cc510212855c181e9478e21479c6bc486901b633aed13c90159ea34b7420a2299519e97b92148cdb5bb28413606c82518c8ad8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf509615f653f7cc5f7dbbb25bf0dcc60ff718614a4941f9a9f89bae67a1d3a66acb0dfc82d60982358f21eaa2220ab9e6cd28cd099dce0d9b94e1375eb5b910110faedffbfa929a720d546681eaebcb73cbe11e6b47b84a8f601df0760aa0804b1aa4a0c42a84404f7d82889eb6f340ae33e9ba140fc510b4dfe6026fc707fa0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53cd686d8b4270d27d1256039dc23f6478d67172713feca9ad0a5c59ad73cf8ff832acba119bce9e040426e248ed56b03ce1f7b415b3ba15f27e272367f8d803ad3fe9c7769a849ec1992c6942998611fb7c937450e6e1cf492a495de744c216ff2d7460f7f13076c160bdb625a3443422ab0ec41eedc592466f7738e6d7a032;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h382bb9899c5ac0e7b83e735d44525c28fba7ccaf5b777343be3e72dfbeabc6bb4d91574686b68b5b51632fe9bd3604b2cd7f1c4dc5cd7c627dc8d5505c72af0114cf912779d231e94ecc9c04849edb00cddc3cbe676a27d448e231bb1c904bf58ac44a1ebd8aaf4ca5fa961c176350289d8368c27843edd70b17abe13552e726;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8275c831db9210298c2917f98ec1a8170effdbadec32df1df7b86125f0828c5fe8ab508a5b607b49bb203da0ac2a6a5ab881a72a1b2bd52a09617d2e6bb0d1e825c0f3d54accc91fb4ea869496c5a352357e035e6f1e5750dfcf5bfa4b7b912697622c4f02641259e785186aaf7012f35ac2f225cefafd93d394800076a02a1a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3bc6595aa07f547535f862bdafb20b0a1232b2e7da7a26bb2bb1544c420ac6e304fe5b28b9a7c44135f806024a2d53cfe12c6f1a9ab25d02c87d30e9ac0f37e64fba274214414ceba1f9cc5e63876448a079e88f55bbb4a2db0160438fcdcd076269b30db785a1dd662f7f2053c71cab6b01278bcf71b62c9337cb352f7bd4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc4565f5b135fa57440c975f10fe4aba6be2e51d161678ac1e9c2c1a4928b549544302fee1f03fd0c69846ba3540288df78569d4c75e3fc6bbdf746fa60eb47a7f5e6aa428a8683ab0d4142af9ae4cd7af33eded64066ac6db55e099b1112d7af6259f511a5ba4fdbb78f47640b9dbf5fb748a336a7e98f7effd63483f8972c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h118a3da974ff8cd4b89be173e63786afc0ea29fa5a02cbe2d7a9d1eb076852a982c2e08f75451a28ae79edcac973213605ec98a264d65491c87aee9cfe5f9b39b2efb12a44f4b48044aa944b8506799dbb24c4c8e1c7db4cd8530d037498b9fceab7cbf791a18eb37e53dd725ba3d638aad31a54f3bdd231ec1ee28e80912db3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe82652aa1771977f0671c747a3d1789ea32ac556e5f69c0b07f846dc1aa1e860aa9054d31e76bead4b0d68b2f9b02a0929e3ec8033a687e6352a70c21abbc255f528bd123bedab278ad6f02c0b3177b544a22b4e296793fb84811cb58f7db605eaca625bcf552cb2fc8d41d840a3635bd01e99f5a411f5e4021b587e7695ba0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf2b272110cc2b7284692d2ebd3cbf6a2e2a95e1f0c88b1056ae28152d6533ea5dc0a3395fc4798fae934141a62e66f6c9cfb74cd1adcec62a9e6ef044c9259bc81dc477102e7f196e43fdb4d6e086fee75e082ed2c9a1388a5ab24e17c8889f94914933f6da37be946e4dd5ec6e343ff8c636157dea0c334791849bbd199b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha59d0f326abce8ad45e0fbb893f95e493557af9fb6d146ae60c578046089cc9e2ec0fad30d540978c8bf79cf659bdadd725a7638e2c157322d6e1c975c9099381b9d4c375ca94d0ff3ec8de87246143891b2a3bed2b2c39fc58bbe18ddaa3b6532e0b11dcab9cf14aa5d95c80f714067f0aef0e68a85c1ed1f4cc204eeb62d85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he26f9aea1b7bfa886f05fc867ae4949dcefba8235532a7f9700744786e7a094bb212fbeac67082fc84a8d4daeee9818c2f146b8cc1326e8294719f832364db386df6b8c71ef0edba938d490d30a9897b8ae9f3fd5712d171f36dd2acd64034bd21213b6daedeb9572a21721dbe1ac4cb33ce696b2f221730571eefb3d50bee81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36eee20cca8fbdbca5a8d6c4a4ecf74206c24ec5ef2d6688bf492ec77c1858cb81b17434d93e6d96118d6c0efcfc1c517224ac93211d4f8a1f9d18c18944f3a905d1233c57b28014448c479fcbc419e78290505fc669a15082d1fb10fca5a1d0836a8536a472d49b3235132fec66409893170538f6ad1b9aa3293228d50f2c71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb17f57f257224bfa1148a8d58d2038544ff936f8b912998428dba8ab419bd1053890c6432c3c24fc5aa37d61c819b6501f26752a7414afd40e219db9fba27ed6fd67c22a1df5909b4aecab26fe30b848eb43282a480d42f1d387951f3c97eede3e6828a3ef16811bf2c10b950d557f45670a688b26f5e7c28b5c35b53d68310a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c14114b4e364161c7ae5caee42773a0cadd07fe7b6fd5b50c159213e9f7a9dc6075f0fcedc96cfd55c776731848d8d0fb01bd53534ea30f32a1ccb35460749e0003219a106fe00d97aba0744fe38dfea8c74a47f00beeb5615a3711efc2b5fbce6a357f8dd316066a83c2b468a2e699fbffb55f0d5025fddcebd95600de0618;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h380b87dcb5d0586022756c1e2f1737e0c9eeaa5a53334a24fb2d1eba9de23fb8fddf5fa974dfdec11aa0dff35e6cfcdba5d7628328248370e4768f443feeccb8e259b678e81251a1ac4de24255bf7404eccfa29c4853fa16b6037f2a4a9f665457d14c72f2bd57ed97ceb0907b05b2abe7e16cd67ca84dc67df0cfeca8535874;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9221b6f507322bdb0c09c8fa0f81136d47bde9feee22afc416d70c27c355b216fd39fa59666dff16cbf98a49333c067e7523a452bd66d8ebd6c8327d13e3a3b5d93cfff2983f38755e932c2a1f223fccb6fce20960e2d125dbde99d5a1dec9916212bc02d7050388500da2660114cac67351ef5a2032064ce77556dae0c3ce9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3261156dc80a7e378c18cb67a2490ba3582eba0130504b577270e32225e937f336465b2d2ac367beca13ae7cc8e8048b58e729bedc16372c35e616d5060efb737f93b875662286727e53f5dc22c9e20ca0b38ac625241d0802de2afcf0d349e20de329b6741692882398ae9dea7a7f14a4ee3b0e75a5c9dfbf48574fd5b617cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22d92e9e0a35e2774a5f676b34b81a432cccd7a40750b5aed16750ffc836b2aeb3515f646e30c4804964e9ed45c3268b63ea1a576493f2d553768823ea8707e4bcb95646155e460a010fbc9e055c5016ea34de576ebe53eecf05fc81695d90526b84e88a14c59feabd0a1599215919ce37af06747ecdb727db23f59e3cba72d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha26017ab63159f4025c8c44370c89f7db38336d2ce45b22ec550d65cbd256f990c68ee736876b3a16b0f33e5d2c6005ecd7460b14c909bac3e9141e62f95f0c8c62fc4cafb870e1cd18193b9140154d60d0dea5018beb7e894b7bc538528d7312378f6df08ca36f9e20b8aedaa876ddb91ca4e6c57bffb8981f555fd9fdd3ca4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d0bfd11e057e407e0aa93396ffdc3925155a2f23186ba5ff7a818cc7f2f339d705672b5d32ed427d59d38aa07ece13faca4499953700258fe434ef23a8683e8760aeaa601312c966d3dfe9f0d0b29473fd664d5873f654ae087c0a180d0b67e62556f5599923092fc632fd6d4e7f245fb467b4dd963c206b0f5749bdfe85bfe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1e1c7907084c2ff525273b82c81f9a8373cdf1394ee765568dfb28c10e94a1764705b5a84e1e0a23d57751f96e299b21e116f96339acd70564df4fd14aab6e196464503a3cf1a02a6e5cabb883cf28d56bd49dab285008815c94de5cb5ca9d18393975d04f24fd32afa4705df72c2fec095887672faad3d62a98c0ddaaa398a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76dc439b5387b99187b21790411fac6d734925528c0f4d12124dbfa7da71de6931c375ed3f3a9ccbcf76558ea81d5f6ffd1778b0f37975371b8a0f1da3fb694f1bdd89ddf35f4a867783cd8b63eaf17ad86901ba93276239638eebf0a96e3ab8c42bdcc0586c02a8e22155f01fb85dece9d29cdc17df94fb35fb67fef581e138;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h125d49cdb990f8c0ef500580e943a8bde4dfb60c55bb69f121935a196b8e891d4ce33af494c20cf929342ae982f97dfabf738f7affc14e77bf6f2c9f6b0931c8f5c7576d66bb6e296d7c8e21040652ad423a1d1669690f800778636adc9939323133e72dbc6c333346cf82610fbd0c9e6a248258b201d52a406a829e10ff936b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22cdb38c905ad5bb48a8f92b6048aa6078418b617ebb9ff0845f442c22250a033fe688c3ce5f3c9a421a14dcd0600127a1bfb916a8c7f628d45fdff0f010e15e3b2812f54319d391b64cf3d92cc900f2f9ced4804b2db247b84e7012ee3604ebe276547f14527cd72847e720ebf0d18225e713f6ba412c8e286095f0dd9b865e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89d49cce54bd7fbfd0d6b0f7168ea8542024dd040f9bba972ef15c05fbdd28cbf3313625e52233d6f3abf423c4f8d9fcd0ba86652cd10f7bfaae17052a9cd37cbc56ab23fb53807f33bf585f0f408e3321496d9ed7135deb9001f4a7628fc1f08a478a7eb587cc4c92582cd730de8038aa383eeb92dd1c5afd8e752d9dea2bbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3e882511463ff011d7a390e59c05fe05f1c8819350bbc69035c26d91ff9afae94043b4a0c26f871d697bcc2238a9268571646bab717d28382e08b7875885afe484b64c1622de8cf43d1305f4428d50f2929dda709b2e6677eb88a06d08ac7d04310ea8b34b6d135244c7d5e1f4894fc2f015b03e6b976dd221d85e3e7da401;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h516bdb0c8b7d7ea4ebdb1117b2e6b147c7ccfe9614401bbbef39dd7a5d9ddfa711e2c17982590d91d545fb18e9c5e46b0815c97ece503b886140eb63032d7f6ea9fe5df4d9d957760caea6afd47b9ee18a3554d091d17f5e049d884856ed00944b5a3b4ce817d70d0430a4ead4e3ad12f224900cc8b45196ac6cba87c57dd963;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14bce40827e12f0f35a0512f44200c41b2a0cf2ae5579217b48769ff879f9f9893453887a48a0c023bf6b35b94cd7ca67b187c16bf6ba49a9f6b8e2505f36ac6cb7ec666eb5036cf65978ffc4b8dc69c6fef130da9c5b957f2d186b6d308a28a0e977a2c597d088767d5e67fbff31c995c33ec72c8d87542cbccb5df922e28ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdc61d318f45f6ca947aeb7902f28131fbc72c23b2e2f51e0daed1985e83860613d1d75afa273ced57a0d432d8211856ce5d70a0370d875fa2afa83a3d1ec3f6a53979d3edc15825203bb6ee5d094c7551f7301fb6b67a108706198600bdce625d65d89d94782fbd3d1122d9846b6d4a11d2277e6dd6f9b4bca7ddba8ef95db7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4565f53c5eeb79f436204013d52e094d220e10fd31e5370d341fca9c7b825bb1770a14ec9fc428f10c3f49dd0822a4299af6d3830feeb7b36e7dd103afc05ae96d53978790a5104a8a59918e445e6f91651795e15771e2564198cf56d674af23dddaa43a4b7181979ae8d7154cc4bd229e5313f92d635f7886ba8aa1cc4de0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e1c7be250facd74cfb22a32b1f968d29de7cb5cf0f3339e1be1333a00582a648109d8a095d7f28ed32b91f6c3efd7e110dc999c9088c5062ec8993bed5dc54995eb2967c0aa07a545801278ed86cac5fea8a43e4e4caef2b1032a6feea4b6c89863afd17d2bc1e9df32d98371b46b0f25336182c638db0d97966c1b6a7a89b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5dbf72a2473899d4f84a83c4d31766819477ff332f75560422c9894f66fc917fe935ea005318e0539bed7cb68f3c7f007428a5037b1710b5817fa82a62d6673d7c6474450ea100582803d6fccd7df344d4c429dffc9632f2121cf59ebaa466f24f62ee7ec5c2a4a6702c2b5e1e00ce90396b51cacbfac8f7ef58fb76bb23892e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4ed539d5b8a238454d249bf5dc734e9b15693488118b60827591004cb3af01fe56cb6df86751d58cb3d1fd690037c95bf823d50ca604765e80abd8f2d3efe8675e400337bd7f9908ee63920ff8b0307aec74e06e772e5afa23f3119479e1ed4ed393e81b6f07f58c744c174a32316830f149ca3db701daf82fba056ff5a8c67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc9441b1980bbcd383b41507e9fd31c99d93fc714dd7cf39719ad68b1be7d523e4a45f601751754f6125e233f24d6cdd16d7f7f373a89600415c261f8ef59ec0c331e0f5179236554eafb43c27021dd8266a50ea9679d3bbd04e3e0be016232e315653689c625c59665ff4c9df199dfda0d523b5a77857fa2bbfcd8726b30150;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca15979dff979f3039b87e7f47dd3a5c9835340c6d50534c7055fa613f1f3b9700f188d77948117b40671c743bd446d6030a021e64ffbf860a2f06cdccfc90239d842b52661378f13646e1aa3d68ad44ba4e2b16085aa3899adf7c361e715c0e8e3d1e3febe33baa39c20aac69f1a6ad54d6cc2f8c8a7d3344af3bca5c2e446e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd622522b3cfaf06da8a89c49c19c5e786117fe6ce13610cac330b31e5bdac5e0903d1b40c8099b7d9c09314e6612a9a5e40a810a3da63f4d52bd3b52429a4b97ee4fbfde2feac522b5862ed6b6f5dedfa15cf62d824178649de447bf7d6cc28c4ecf8cb8ccbccf5059105250d31cd599b53454913a2e44a034c77a7ebdb9c437;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2416c6099130c31ad72dc7e437bb7a22c1efa4af7c1f9fab18e68e33f88d9d6a4b11a6e350efdf4e2d1e7e5dc1c464cebfc6b54e9eaff0c2ceca558fbc9af78cb9679ca2e3ec868fc1bea31ace9ef6337d687cee02e59dc360cadf0fcd151ad2c99bc9daa6e1a7471bd667639fb3c26f285966195e056638e70934cc895bd866;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8aa3981e33ca3c94830618697e5934989ec900c997fa8d359ea4b3cdfc01c92509052725dbc9702cd822b1553e8f58d5a6e7976967781634901e0451f44492945617520f34ed5ab2493131a8d212e5023bd74f98002026af3c248676a77394bd49952de532fba126889b82282c74c235b65290820f24d6e214c4adeeec722ad3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2de92d23ad5ce56cfe2a7c16471df8cd0e4546e42508732fe133c2c42cddac249c712916bc095a80f91e747979b4218a04db72655e766f514026cc6e938766940d90fc397266bb265d81f92a6e136ee381acf1a745508b3300012b8efbc52c5555b5042a17c43069a20b4a3d333433b89ebbf7eb1ae5b8d1c624d70f1bebb288;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h948df664c31886622b2f9639edde5e45f4022b44729a7c5c8a08551fd996515d0ac7033a276390db9a25802234cc76a7c9328c52670a05a2909f86dce7d9de32b04af5e5ddb716e8f752877bc87b66925642ef22a316ec278c1e6424f06ad8a6e419d9b04e7b5185b49e79fe9bebf862824f45115c44037f56470186faaa5f6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h240b7d70f5204bea3fb0b5f3a1660292a67d4d2887be315094c04799f0f13cf1a01a507bad0b38a78d5403cad4f072c58ff1c6a8a690965c4cca2015daddeb546007416717aa5c6f0d0ac4d1e2f0db16965f9020f034c931f28c5952c3f0b3cebfa0e061da0ee3643c35393e21b271bb712eb33c1957aba70792dc4ae35f0dbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadc5f6c96eb587e0163a7a208e97704f74373bd28108de951245c4274324e2d500027b77735ccd5714c4eb9409f901a89eedbef9f81f37c4049e8a7918c1ad6ace90635774a28ee835d7673bf3cbdf094a5ad4d756456b1de1f484b057a04c238a3fcc53f6133c5fedcfedda29262b7b2a615844a270b32c318db13edd02863c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54910c9faeedf5cb9458c53bcca5e02cc256821982d3186faac7ff7156dabeca90b92532de8700264a429fe46d6ec640c56281e5fb721640ec9498935064b3877eae1a75cde7d8f5d6e1ae78bdaa14d3d14ce3945b83f8cd732c4363ebc4dec5f46e06cd1ace85906bcb338ca2de132863ff179a2ef6d16c36a12ed7c6f5d10a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5f648719eda490b4096ebe72722d4cc156cad0d001c688347943bafd45f42ea64b60174e075982deb5bad6ba819b47c278ae60ee110083899281ac7f1e2e2f5c902051334500066b4719010f3129ad899d40ce4ec539cb49874d0a988ee02cf8b9aabe943869030178d4323b083f3b7c813a8be7d4a1eb6ce0b4051c218cb31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ae82bcaee3917854278d893dfe3d16316dd2e5cd79a64d624ab654294b68c2887c9209cc56e12dfb6c609463a8c6d4ed9feae79de11a9e8fe10d16f82f2442a9eb813846aec87caa590758c2aa857a449b06a85e3501ffc29427066eb17169cb4850dc5d3c4fc506bee013837d1fbe9da14c1afb7daa923cfbdaa9f54738397;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13dd1bc630d001d66314b243db688d4e51a1461e3ff922dd575da3331afa15e201f5a3ffe5bf13d44540424f54514428367122864cb67ffd4bb5c3849872d93ebc8c027afaae2130fceb23d68d9302468cc8cedbef7e6c85b8df0361f6f59fec12029adbb157e9e257c4cb4c13ee377eff781150b183aa31c22d96f624f7d4de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ead64878584b8a2318087bd7f92484fdadf798b15448fab08da100e5f76c517c2453f9ffa2b919791911e4425c9deca7e46e4480fd6fd778a0a91cdbcedf1f6d39687f493b4e7042d93984e99ca2835210ecc5c113ce4e6c34aa882985cf6a02413cbe16c50cdc2890afffc7077225cb2dcfa6b9a895e9458399d0cd4053a65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6517f5b389190d8b36c284b8e832976762402760c4ee72c4429f347295fae3c475b4d89ec7e3e44249a2a2c9de9e9d06027a21fd546adffa0d8f153aea99f23477bf57786e75327f404988a4c0fd691f80501563bd635520865f65bb5343a9d2dec8bf5d2cb1d5ffc3c54eddcea2703b8aa998396b180c313f468da43a10fd62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb87cdb67a55348c90f03096fc61e5ba55b40f2121d9794762ef4c13d7ee0737fc14da39793fe8877913c3af61dfc7764b05fb306b92593122224e314d7280a46c2e0d9a59e80e9a0f48c0127cfaa0ce0f2a1cd48968fb3e360e6ec4c44b23d11a1a424d4722570d56dee6dc17af682dd9f561011da6f0bd37a126133bccdb977;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he608ad4491039c667d2234e4d8ff8f5c2b0424af19d365de60524d0dde105d8e27598317d84cb4d23f9f14715c7f13a5c83d10381d4a76f535afcfc5469951b474c81d0746a63458fca052653b242637ec89bfef8c021e27195813c6b9804c90eba5da734cbb03671b26f6b0c8c7bb8e37dedfa300f7d18a2c4939cd50b3c8a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h925b42385fdc01062a6e81090e168b10613c33f002d258889e3f65eec69d9fb82ed56f8fe092b0ded88f6835c80831e13e0efc7437f63107057ec0334dec0759a966e50670377241af468179c5dd995ad02845924cefb15f11d82c97f5cbff62dd4364a09f21500bd5b92efd78a575246f3820bff509c209422fc0efd7573380;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fb9d53d113e9e958af897937923f95966e8117390e4e67c1bbe927078418b1fd033f1e7491235ebecfab30166e3cb8a351d895afd4d95d24ec9eabf5d615d90094f56f38255db5931a17ad3df94ad8d2dfe6856005012af1a0b37052761e684b6f031d19ff92c2686617fe961ac5dfff4c772e6e7bc9cd2fda6f36f2c8343dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h278d186f01987ef1d4e9c3037d47c8a63ad590d848b0046c140cff8bf9b4a837eb4b2f89c2b876cead2d882d7a0f46607ed7ce73145e995fd1e33f28fb4e673ba8741204c7fa5c215590053f65b44a97b63fc17addfa5b5900b05610b5d836ba4b75115133874bddc0806e663b96a0a10495820258ffd7ca3e21810c99420388;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc46263753b88ddf599fcf5025db222fc3740484a3dfc668179a078d11e0faf0a2e9fa35ccbda5c6acf4fc61b2c5b206ff04b333d75acc31df1e9ca1d83b38eec0d566d1c812344bcc3bed94f5434927209fca2e1a400aa4d51c94d4789bb162521e716213e8e7a9e2bc78175bcff9bb1bddd57ce8ecffe86b7da15e059fbf06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1a0e0a7fc571e3a9e478a3ecad4e39b70e26fc20094e5ecad6bf99e25f2dc628e8670580355d04430dcd4b61b5fa076878c8057b0307ef5c00975ae23ced414eda548c93a6fd66674f635434f83318d5053796d95d00ab795bbe76f99310ab47b4080223b8d72d14b647decb78b45a13b1ce015a7b6777f1693d708862d1289;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1087fd44b4ed9a60a24399d2409f753314c604f00eca0ff4c71ab50a39e353db839676c1ec9d0b503a1449b1844a0e96ff6e67ada93185a064dda7b4416c5c3465b9b7d0ac8ad0de4e10a7af30b180cf385d2616133b9b911b2ed51adb0e70a2f3279ed1ce9ae51493c759220a3ca0e11ce3d59e1b6679d7810065c62a5227f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f437ff85c191b03c8aa6305210d6ed41df75c4938d6c6674961746e73f5e9ce90d9776e53e16620e85cbbe2df5c944f2f7112f98bb6144f493c6bdb4370208942cb8cf709e29d4f522ea527a0da6615ac680196302d86658f7225f37e24f63d284a179a29c5e88b1bce605407c5b8517c916093c87f1933d99d3500e9534a5e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37973f0304f179ca60c79870200060441d60cbf8b7880ddaec0dcbd7f558af965355e5b652195a37c10fa7fd709dab7f6f5d0f9217e419e06cc83a21d2d25627fae0e44f7d3e43b08d75309c26bcfeb5b3a994096d42358f4d0a41ba2b189613fb8c19ce8c0f0fe8aabf037f9aaffe9cb0e258058d2b9aa65ca676b7bb49564a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h450dc22be96bfda186414acb57cecd2e36b9ea3a6821b6158d83a00516ef5f840cd6046d59acc521f65c94e1d40b555c49fcae4aeecf02b4af7ef0f90a509213d7f6092c680251386605edbd27ba3df1821a1df5f31811caa9a26b7be0d5bcb2c7ba0c230427638868fde801a62d5ff95e9035053b503c1fc1ad18cb53a2d699;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b0b9ef4fefa4a407bf52294968318ee4daf3a7092007fb4a1de790a84425163392ba7f4d49e29aa1db258c6cdcab17aa459e876104b71de53dbec31821370ac7928358afaa725b2290fa68de32bb1970c739083e592913ee0ab1c23a7228b33e52c89b028421978c1bbf4b917fa68915e9ac7a0830efa93ccec4d51fea26348;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2697e03ee7b4ad8c7fec8c30a4c422ff0ca2aed58725b29aafe3eacba7bd20c9645005f71a6a86ac2063d9505534af85f01c16523aaf2f8d1992b413250cc86f1d84eb952b983e7ad9a1818d087735855e08276ad2bb00af483c92c6dcac66902eeb30a25af09db0be3470051e9026a9089422cc5018b92dec316a802fb2c01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h682634e1ac992a1e38f39087624e3b9374461f906c15259a85d39fb52e3327ee89fb2e7bc58c2babb2be859afb2058938773eeaa2c70ade56373d222029393e1839b529e6c2a36b28084ff5da777120ca0311a3c1ede9c0cdd907eab52483687bb7aa78a872b81e4af61eff372431d1e721fc4817a6104e5e3e9566bd400b1cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadb068d810355fd8e44f2b5729c83ab0603e29a085b006e02dbef1aae6d498b62923e696b4ea303d5c6473d923c7dd24b7b201d3f11ff1277623f90db98be20fc39267654ba1c1e9d95237f788c411a44bf4f955d9aa7218b510b29e2d0f06f8792dff5559f05064feb0e0fa8d2fe08f55b2875ed7d2bab3b909d069144e7893;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h678a049f29ce0f7279720928f620387f11cf084669948389fd65f9216a871b3c16c08e8544aaaa8567ced30d616431a6cff033fc9f8554906d6e746da76bfaa7cd5b369fbd4e1d4a062ee4543ff6f9d8c93c39901f6709a8d49dbe16cebdbb82998896531049c1be741d9d54cbb9dde0e58db95c83f37d646068d6cdbbc875b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b6a7eeff98371e39dbb706949fbb29f2c6e913298a113df3e23a00800760fd7ddfce899bd29ccefcd76a6c9a065be7be69b2f91325f9e16d220c902a7b1d056481813a9be7125b49ccdc32f1f8198376ed8d7a2faba2890ab8048ec2a71b6957d1a235662ef5d2bed9e4630f1dd703db0ac2038d18b71bee93b53e5bfe60bbe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f89b02f19ccc94e17f4938b195afcd0dacd1de3f2fe60bf820e93cc0081c91a5881341dc0e7c16084abb081499aa7d02af7011f2416c07a88c71119f78de9425042eaa929ef572b115a5ad3e15421b54b909bb66cffa9480e5ed8c73ebbf2143bfd1464fc82589880199577c270d046cb15dd315c8508eabdeaaf8bf742655a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h835cd4da752323335b0d8f43a6c31a93086575e90d40a5f3a7d5430a92831466f3cbd72aa70ded0b07e73402b968a94950a7a0e2134d1cb49a0c7e90da37dae5e33487ed64e651fdd0a4d1ca380d5a3b8081914c6753861e10f0b2bb1a4b6846ff137ef13e19b7ce1719206af71d173e526f34c6b5fc12868e726ac341c75d88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b80b16af59709714df0de03391a2ce895620151847dfe1563348178f0bfaf01d40ac8ea4c9c82d38b37ee206e20d4a1ec4072c1dcc4a329db3142e95ef5d6414a789c2390fbeba83d36fec8d866dda04e0f7930eb97662d0b1bd635dad110ac06b3f9d807fe7ce1efafcda70b72d140e99100e552182b4a5cfb962d5d7ccec6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90457cd2664eb2ff36525887dc2276be0f68edb846adb95fc54fc35201311f5f4c1ce029d6f93dcbe570f9787e86e3b4fcbf306dbdce7425df4d8f93c604b4ea3d108b6dcfff1f83874676ca5471590c4c0a8ff332b4f7cefe291da99f8ec3f765a4b829b79917305c4347b287e7d08df2b1c38d1b4dfb3151b3e9fec882a790;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb400d1e13b0c59e77b58cdd5405904a5a59c3f77db1877e73c0e9d02c1b0377c0fb1785e475359369fbd9b0f2cc093a1a9dccc01188f7644592113234309acd7c078fcc7bf859ddc18e4ae3d3774d7434b3c3089331ded1deb13479acc7dc73b0c66957492a2a39e9fc75e3f28b058e1f98d518e9224f37ac2f41177a416881b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb993b2fce657b1f1fb183890b96369648937609e5b7fe9bfb037d6eb29779833367a5046d2c4fdc69942f6f73c4408c4a7328da2513b0fef42594fd9f492eddbe4b83e8810cedd258867a5fb97322bfe5f28832141b43df8c5d369e6ea9b7c6181143d37037be36be83c7a3bfe8c765cfc22fb77ad212639a82dad874ae306a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h176c2513fdb1aae2a523c9643fd5672082cf1d75462212ffef17cb2d6b6813b40724a110f0f720907d3ebc402e6364a20c6581858e9174aa259a9ef851566c96a65c77d25abf6c9e020bb86b9cab6903e1dd63ad071f83330448ed178b1b634e6ba550cd98d9b59d9f6532213b5669f3d43b9de9e8a255818fb360afcac7b0fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h604a71b359d14b59922c40dd98a203d439c66e445078a3fb3c5eed792a83d4735d593a14f66c5fe5db79f7462fcaf2068d1562acb4e4e613208b99a8733b6b5aed5d533304c7b4da02bd3197aef6b6fadac94478f84df675fc1f278b0a024e741f23ec1d6556dbdfde3591de1773ee9327e3365cadfa9ce754b1f90b7e01595f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71951d2a1532e246d3679e1e8bd955e18188992b99aaf892386c762ccb80a7239ada04b790eceb91ff5a08212f2302991afdb474382207b9ca59bff126e6a3e53c443e82feb9e824c5dade5f3bde5cc6495ec9c1b675bf0387d89a86b5a75b6b5f29fc137603dde11e99f1bbe505c22b491fe53284b31c4e7b0e5d7a7ecd3706;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69e9862fbb0e0a8d573466242a7d79a11f6bdb1e0aff083b512b3a50843ea444d1e63bfba166842b521530be31de850e4fa3b5c5d53bc95089a1ab186f517b3a4173e268ca48fed92a9cdb220229e5b7416f04001d922a5777099ca94d0664f472bb2ba4bd7e33cf8d1139f843e8133701d47e22b4f1c598f80bc1dc8f6a4832;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h455e9a672dfc935657e1fc041a1a636db2dcaa72e9d80ac35d77da0fdde4736d7be6532425782ee7c9d3ec72152b7a45379ac4dbfda36fe0a034d9f405f0d0d37b6a136084f3cd6375ba4d63cf245912bb2dfe56307c43611c9cbf5dd4c4c8fa076b0b8d04e8750d2d951693cc69b9c5398c73f5d8a33c410addc5e72aacd2cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c98e6483dab6a84c6c9d995ca3a44ae62a285879d40958dd0424b2c11f1e5fff3d526cf3855d09496770576ea8a5cf56eaaf0aa8e326750f80cd23d8400f0934adb22aee4dd2a1248859a0f096c9e74fa31a05e3c7546dda435beebcc08c41837d9eb5ba3fe6d001635928147fb91c9ead88574fac148ee302e5035b77d0b16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51db5fa7ad5b36ca701ef5a52dec5ddbbe5564f7dde7582f8261d82811af4a68002032ab625264e780663c14d7ddb6203f25598deaa503e1c4a8937c98282f14936110019cc07b277249ec1b1415b2ea4ac0ca5f61cbf1b89c9f964537d475e123dd172ae46ef992dada05af7a2f8202ffadacbbd1ba724920fee44e3653498;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dd8d19a6647e8b62468775790cd2b33ac462a47373302ef36b9ac8132c54b6d2af88f8e5d67f86e2bc7e2a0ab15dc6e0172946e6f29c077ad9fca1b443349e9a8f353a01f67b837e0e2b17534737ca16d395fd29787e9026690ef42ad09a908ec14181ec11f72339390aeba3c820b9809446284ae06bac1ccba766eb4599cbe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27aa9f269ef1ee754c824d680fbcfa55194d5058abe0d16e03409ea99de0f8a87af01a98aaadd23d36d492d5f6d632531470c5f51d8f302daefaae74256359b1731e29b772198951a3feed01e682d0a079235806f74b6b5208df502aeedd50c28c498378dd7624691745dfe82a6184c96bd720e34e4b2407b8cfd561a9fa35bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7af151f4e81e0a6a407fad937bfe204d6622a2cb87db7bea97a4aac23cdca9409cee9ff70c976a16ddfe599f2fec56347832a75ebe5c3e588ae8b43e148d32181b0caa157a21be911e5421e3b6e629d49fe494cf44b7dcbbb3f691d5679eedc8f2eeb9b535d19dea863322f780e006ea0343310cf7afd809f6fffe72108366e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15f593e922743c995ced920f84ae6399fb81beee794cf3d746ff302c5961a4ec8422931772f8b94bdd8937b343abca6e5962baee1cd673292c7551fade6242a5a6a06c478f7d42e8859f97ebe2306da4fa00302bdb8be8b06b030312d76982b995afe455a8d6136712e58a56c05268f5112d7c4f709ed4b16146c28fa24a7ea4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bc2ce1878cc5f2665311340343fe7647a957b1b431465ca091c088f66024d3fa772998792cfd3370c62bbd105f98cdf2ae253142c1ebba029efc496a434cf2a5308cc7a894263865ab6e879185747af3de562ec9bdd6e7213934f12eefccc6e6e73ca5aa7359a0ddd473ae39a0172aaeef8fa599d3b549c91fc0ef149260b3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45d78945d17e6e3f6dc3e3f7513bb0eba0aaed7b9a312bb0f14598cdb08a3456b01bd550e31f26604cc25cf6b52705ca855a338ebd2f5e516445a1411d35d4fb1128006893b84d4d3c4571189de5fa277b291dfffbc649332ee67ed7e329b63d7111e679e9300687c125315446b29b5a2f66a583199e8ec73ac9b6fb06e697ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f35bfc436585d5c346b1e5753e4a00cb40417811764473ddc4714cf890606b0ce65517ad78087c262221944152b11ada96ca44a6b2cbd7efcbc456ab73c57380753c80b16130802aab3c4a91d948de3400014786d9defd9f1b40ff34eb46243baacdf9f995aca14c960a09de0abce6d7b0d74ee846100db746a51b4fa2bea66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha246f5654052ba44f42d8933615bf68b80a9989d3d3a38ed9747c1510752623053209eed40178c8ad833515b8f19765e36bc0db836a5e2e542407bd55e6d20aa8f9da04e52234e52fb1429d3fea3c362763379301eace530b5c8b27ca696361a846b915cf89c9a2c436064361a5fc76e053a1b750a48c4c1825a0e277410c00a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc20ad05a1abfcc2163faa79e0b7778ae7b9561f1949d067d5682fb083639c1f1eae54f36626996c49426e7df4db39e567321147edcd4b5f8f6eb9a2fca6854123b9e5c855f2ae48f3aab634823b185519f87e524225b3ef50e3aaeabb889d85263c8d25d514e39c1d670d4a70814117b9462ff752e2bedf80e03a1b488aa28c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2dd067394746df44cfd98c113625ffa42c1a93257f011fbafaa7e8108a031bf9f3ed6cf482e9283e1fb80bd9b792f75276e2b04ec942331ac1a68a12b74ccf3385fc2a774fc6940dfb648debc4d11c6c5a806f1dad5d1736a9bcc5c552457bef13923b4cf088807053e240f4429e956cec3508e4e5c981e5b795a345a963d0f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3859438e470adb4ee34e44aaaf052e6e66eb0eb02ad5fce5456d7d61bf99989d89ca4633eeb5882b0a6870eb657c2b5ca8097232c7e1f79c37dc134130838d831fae25c21c1ef0013a924a3bbcd7f2ed275b133a829e8a2f4f8660177a788d81e634e3565c436c5a6106616e7a1788c9a7ee2f100c63771a1394c584847228fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36ebd3499e977bb401246d937f3de87915f912ede1e8ea67c191ec6b689d71cde81790401170350fe38c7f18487e674967da9ce742782ded26b0c90bae53180298c1d7510815157e31ddc48694cd0e6d57185c088f0247374c0466d4c89404e09e5f53c2b6ebc4bcbc157f14e395b54194d357be011e6cfa58761eb3aa0e270f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65103baad38801d8a89b7dc32fe5360e943e79c49a901da75c8d7834db3f1f9257d02d21c171e8ae5bfd9e61e01d8d0dcae7634d3cdcdcaa75e16f0ed6cb93bfde76a45adfb9ad756232de77cb58659c59d4995b86dc08534d41e4e925b0d571fb15087e252ac029fc5e37a3fb72f0c666aa09e8878639d0fa50cf9ceb350021;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3da8d7a20ae0f985e89249d5c57642d27031d5b9184c98a0bba0338d42e414c885dbac27c25910177d0932e7d922b54914d539c3d0fd6bf6482a810d560aa75bab8b84b1eb06322e93215ccfd95a57662debd323e0cb634ef5c1352203b5543c9a3bd87917f5fdfcebcb83c0d2b92312dcc5934e323e9482e79cad559fef27a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21d804c5f6ea37f0ad145248770479fcce84ba6d23278194bb754f108837a78c7b61818f83d1425f1375832f9aeaa9eee876364c4d9b5946e4742b935bbad967a3ceea59a7f9a5630b613df2ad4f99f63ef89262e0e7386e26aa90d1eb0bb8f5fd59f5ac17fa368015978c9e7e09c6abda88573f22dc82f1f03f7281b80ee43e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17f07161616cf17be00a44749590cea0048f9347ee5b74b44426c9f1ef48ea727a77a7a6ec9780217717e2cab1fdd5d66bd860aa9227fe74060790c8b5a91f89523f5d7a6396798564b87eac1de45e195b827b56ce4340e6d11f27488132c4aba564edd3ed447f32e9b574df0e501bb8009f5e04f2853046f79bbaf4b34816ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe4bed9e9970aa02a4b968665574ab9b133755c1515171649bd3f1a27fa97d7ded1af106589369731689253220ea89bf935128348b18db676d39fc305f2da0be603a9fcf122dc632641a334fb86979467cfef4eb26cff4a5a1ae4856050d9fba40ac5941e5b7fe6ccb031a812c8e5dc7270a0432cba91042da239432987f7828;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e6273e1df29b202324c594dc2ca99d4c2cb829cd2eb9cb25238bee435a2048267038f76ca262eba960d2f3b1e409ec214d4d05ca1c889b81754e9f86bc2f8dccf44b90f82d189a6f8bb3ecce783fcdbe5f9f91f0669f917bc7f0696a07fbf9a93a103494d4115abfb9823ee5b0965734d27cb29a1edcb945d6c5a1ec7744004;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h395aa5636ff3d357c0f7224204f259cc024e633f30ddf4d9b5a29703f776d9d7bfb2da68f296937f123e19d255d434af374de8400cb9c9f553ca674b801e6d0a0c0d8dbcd6891a1e3638eea9c5fbf9deef697964ba05c0c3b538f109c3e4c730e3683bcf6e2d107b2d944e40bfe1b9752d03784ca5eb19e0932040f569890cb2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b8d35cf556afc5ccec610d33fd376ee30f817898555c99e74a6b18e1edae9a73f20d3cf792cd81b5ff05d269d830e263393ee22618a64847c874567bc7481d31f5992ad1aeae9cd9e7e881ed99d52d855c613b3cdc10c7af2e7f6082ce7a1c29045885183f39b0cdabd84f969f7032241131965ae413639e6860ce67efb0f0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b19d537394d56621583ec42947f2489978184c7cc788374d30718bf3917d592239230e0aef06d4fc959623c879c1f7b9b3dd40f148bcf78a3b6c4dccd3c7edffe9ce2a1c3c215121bcd899e36790535900cbcd32816cf43f50f4453a068f56ce14e8c8abee450cce7b05b65a6e28bfa84469b060daf1d81ea145064663a730d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26055ccd123d53350a5aab49d1aeea95a886a28a4570c10a7abb0599bdb98703cb1ed3207c6407f25b92800d82754b783a4e418febfc63272102269513aed39412fbd952a1c0981c4b27826d2b3c3ae3ebe21d42105328e26242c0a1721727fc95e4a09a067b0cd5c3204aa30a8b1835f85047e9435a4436ac3c9176516fa0ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4b8fa9975ebbdf2a3ddfd58d8ecfda03966a6eea6d53ff7e658bbdd33df4cef12aef9c8a89a4382c02bed22e0f5181ab3ae9e865c434937868b9d3ebbc64ed98fe1e801710f7cd4b2db6fd6ee9355c4a3ebd1a2958989975b00dcf9de45d0800c01b9210c94251bc9d17af53d4c780c6cc622d292d51dff05787cceb4245ce6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d47528d4b2dc5667aa2bc95c8e446c3310c99849fa9f43f88b08540375f678a3fb1562e30f1d9754431692dfdaad76e09cc9def0b4f1b50003b3e30c62632dece023313f32464c4516689861f1617afb5296afe81dc95a1007e7f4055e87e2dfa78f0e89ba366de9f5c6c8ba280f46bf0478c2da63e3305399fef7ca04e382f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h236bb2d926acd6a58f7bf68ae65f5a952b84fdb0fe3332b012027347e62fcc3565de0608f8bd85580169cdc3cb10e8b63a7e9cbaa30dc250ab0e3d452762dc8bc1c7a3509df51202adb1a5dffc9f3f06dc3e5a59827ec7dd20eb76def95d5f268dad6cf0a6f73741d09678cbcf027a21513520aa516a16a3659fcc5bd917935f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2720a0bb73fc43d43d91d3a369f53901fc93ea4c58fa5baabc0a9be6cd67f8d889d0b6b5365c0c13041b199748844b7619c25156caff1890a9bfc57cb34e00e54b0707205d4ba55153fdd009b8ec9166fbbbaa3d5431f3e0663f41f7d5c83882dff8418907b87143cea47ac4ad8fcf877f33a7a1ba4bc091ae2a04776bcc3c65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5af8ffe064e063c24ea892b98f1ddb96f993e1cf304424b04594afce024a57b4a8026f444939be666ce38e22e7136a656a643736cf278ab7f61b670cefb6707bee2f87218ddaef1aefbb4982b88c91e6ebf9b58a176a959185b3d7ed4d90a05db02fdc8e00e7b1c2a43b6022ba98452b0e4560c6bb8ac0e4ed915dca56ac3ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22e74ffd5bf512769f27a18c45abf4d509d143b3e00c55d94fc9458e8a94c554d1e6de4d0a454cfe25704554c47289acaaa118493c8a6c4f1a5757c81b5d68c37107e5784a958843b46c94e1cb455e9a99c0d387b47643faa917722dd5745172c6f37d3a9226f83d04440ea50e3f229647c467f2c1f57eb065136e92c34ba89f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94167e217277b3bf34bbbb17f0e8b08b63689f96347b81bfa23f0d7f3421d5a0d08e2af4c41017e989893ec7918665543676b28b61336950288ea6bb437b1e67867bd882f70c3689eaef8302135ea237cb5ab25752f7ccde1d26ac9e3121278e6c59a3e3ffee63b2942e93f8dc4250142a36ec6a1f134fb1f085d4afac7ba5c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h189f2ad956bad4d1f846198361bbb6b50bf8c6c65ec985cbc7b567bec6191f83d3901cd3364840916412b5d5a4375d62e80400cfd760c042518173e9ec99bea4ab4d45e25b1c3cbca883a1dd1079ead2b711f10de330595baed25934ce437879dcdedb667c573996e9d31bf17b49b4d81b12494307fa353a7defa6219cd3bddd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35533484e0b342d227194bbd698c3dfa391e6cd5603f846c914dcdd1d4f80fbe293a61ac5b59822940784b437bb621b6a351c30e140907670e468b50ab4d3f05abdc66f58d45b79c4966b24812acb1c7b3912ffa9577dabbfc179963fdec77d1cab39478e1adfcede3f478c0e445c5dcbba76bacf5065d730488fef16def82d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cf4e53d4f19ae07d724c7a50165c95513d436d4791506f18c04231011e00252c1187ca7af5724f557f0c7e2e56ac2848980e7c17ec4a2a88f06550f389ebdb436ae9fe2b8d77d7a83ac7bbf4481a49c972354e84397607a5d5e6810f9739850975938891896d9b36728edc3d51ffd4d00ceb1a8705b4d7c59d8b0590bc60c11;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfece0121085553d01709cb354bb3032bb6a840d7adef6a9a1891ad866e33936b0573504d1be490b95ea16f3c34870ef5e29333584d84c3443f0271ac8eceee636cc5c12c81f758eb099ddaee8d113e6dad9d0599fee47c36d8e6f8386a554fbb911576c47994de9eae83d313c0195c2c75219985b06338d9f10b6eb6c592540;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92e4575b9d8cc6a62b73c241f69eb087161338519048de213b1fd1a69b224f32bc4ec445bbb837b370e4673ffeea8a70b053fa887583d17d18ea7f6309777926407fb3200d1756bda1f3debcc5c37d01b3d92fa0741d7c3ca0a5fa2f8c000975dd42cfb9ff0dd48323a88efc486a0ae7e0e51ba9f804f5fb6ece9c442544fabd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b2ebedc478561b3978cdd7bf9bc0cb1c180446be52233a48dc65eebe1dd720197a987dbf015571d823fc8ab30c52f01cf5f2174ae73b6e6ba6ce4ccf01d23933dd763efdd39f8649ef32b1c751d2ed1e39f5638f87339774d0dcabce9bad95a2a9d9ac6b225342145c35a86109c176be41ff2a5ad5097386a7f3695595e6319;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he53beffdae8a9773b6d38e00978534dbb934e52c083fa85d96e7d3b5f2db3de2611368329bdfd03e8e797b07c7ae5373c1f88e59099fdf7821409955c721d505d0af70c6e79f70259d19afaa37b1cf58e797c994b0b88cd8c998dd3ead997fadfa8e6e2ec7b6a7bd10cf23e8d90f8fe9e42e7667a5c212480d401b2c8aa51192;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd05cfd65f5eb257a9dd7e252516329f87de1f59cb8a9414e096368647e2023fef98bf5d22ed3bc178c43a95835de14da3cd8dd14d8b26b04ee155b8fc6f5443d94f405b411e0cc0c1f0cf15cc3ecf17d9b2ec104206877e247a6dd29dbef8f11afaa941243d7368ad87fbfb7e0eff1ff4d63cd51fdb3ab50c86eaded0aad0850;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h297c17ac5f3d7c3aca72d5a96dbc936db4c37674906194ff0946fbcdeda9ab8ea354197480b6e8fa2a575dc754fa3c120d2e4058a67cb0aaebbb848d242ce7df57fff95cb7e4796b49eee715552c21c9418dde5a3865ab15926ba22198d68d12901823ca70ff13cab18ac1f72c13dfc608dffb0f3db7ada2d93b66e72cfef5d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd72375bd193cd5a549014c4c5f5ce5bc613c7f27295b29965fa5964868f7411fc93e3ec1138860a0ced3fe09a8c1ef30692ca5dfaaf6d642230902004077ea16e6249da5049321b52891e96d203a67df7d25e22ac9ccfbdd85e03908fb8697253a256bb12bb6aba30b5338ee4472a1b44da582decf546ea80b1c62a5e528272b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82a158efe05f12bf317a063a153c69303723cdc3b86a16c327fc96d33c0de820d855d6dbcbffb45a007ea8c820e92aaf717daae535f4f2c5d60ccbb8354697952b48420ad15b5284de20e24b5c6c8cb227c366a7dd68bb24a6828e47aeb7586273594634e4a7e01b1e8137db49865c0384966bfb2ac7327dd26c872314835561;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bb843753860d94801d3d8bddc4f4504aa8020ba00ae65b4044e24a6e5bab6cdcd33def5d7390ce814f29147cecb082b3e2793463f2e5c104e96d2065d0e5d5402fddb7a3ba749b6cea9f22cf1b16d6c38ae7777e24211151df633d66601935cd3784fe5c5b3f2a7042aed91fca0439f418d98a5f753f2aaa6231b381d15ed2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a186286ad29805a478b0f75474e3db7ba559317bc3df70f5891657b1d6b6a21ae3bdb35041d4df78e910c8a03b3d4df54bdb80cc5ec8077ed8e91f51e61ab290990dc473795da6f906330a417d1c64c4c0eb49ffc70f5e1260783ba62b5736fd8bb6a761b660191a23a271fd9ca6b8522665fe94db043a77b18ee31b398f538;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7f9825ed6ac36f01a9f11025a12c09b2f310ac8b0ebde728e2f9c897a2e3739e10541cad28693f1f88028714580023fb3ee005e204b15be5cfaa6807264f3fca48858f806983e17776d8abc5d95f95afcee2748d22b17ae6ee83393f5c21d90a21bd4877711dd7e02cbf04138998f98841620095c95c6829eea5b0b28e8abac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c4c74e978913b19626af6b5fe8f5a27a9790f9ec89ec9ee1308e36d3e47ba34cd166e645587542298f38a4c88922b3b3afdddb5edc1edac4a5de90f37ac9aa6bbe9485a6fcd7e038ee198236314dbb1117213f04416c3bf903e023df656e40ed9a26f3770bea3a4aa85b7ba2fe20775802b0d2bf8310764190531002a33ebd1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb42cab392d0eb3e4300d42f001c8c68dabc1217c12c182b1b1b27e444508849b3634020ad44831bda66639b1c6bc6e37a722e1177274befd234d885fff181582afa5c98b9c2b4a8f39c275e93b777ed394d22a68b12a30c4ec7495c76308aa69a96432e8da8941a9d3c4f760e4d7766053b86b356c8f6645bb18138fe9c92cb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf65f9db9b8d42252baf87adc760af884b18f9b2615bec96acefd09eda2ea44d90d5a8620750cc44829d849d8544269b0fd8f7a57bfac7f48a50d48cb41e58a0b410dabcc9bd2f8f9ef1f1b6d19c37a6a56012d3e3df3e855ad1a92c7e220404443e9abb0fb9cd64125ea43a5fbcd63ace25cafbc763b6bcf001782ca89af69ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b17db6b85a64b8e78d01703487db37709dff9c2d3db521039701afde716ce78b7de1a12da58e80b9f7ad951e79b147dd2c59a3493ad2ce905a0765dcd03a301f03dd72b4ee249b47781a3a3242afdc5e60872690990c595ad291e4c58bf9453fdf6e2c45815ad49cabc84ca61434326a254138c022c2056b5e7663c20318307;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a1ea38be28704a97c53d92800c1bebc98485a2b02562785ee81ae64f8da31cbad398ff76fedf80050bfdf6e1ba3bd613578743d05230be0141aff0c7eff8e1ab63e347423b00a3d02dc1aa4023b76fff15d2739f65a932655b87f5d4566d3a223408d6ba2f574f58d56ff0ed60f2f7d3ff8705a2e50a2239108524e6da90636;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h122b2a0d99604b7d9e7d28f2c3c60af5b41b4e5c35443af41521df9f0f037cfc6151a5140a881d4689f951874b07b19148d18106c72e0cc373c3bfc581641cf2562873b956f464d7c543a20d9f8d3696c297001c6708347280b24643c1a1836ef22288b5efa3b7d965859c5cb20275429220ebb6a7dc820684f5a3feae2219d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b849f7df3a196a23e64696c5142ce8b20a820cd13ad0b66046439f6d4dfc02dbd1f2512c627f86b59b3b2f38bdd4fd3d9f36e02e02a389f48ee4c004fdfd6d5d7aa2c1930c78396e21b35045c783aef7a40d7d7610e16c6d976e03e9a49f9d37fab9adcf3236f038d41cb3f57e4a37e9f4a7a3f688be11a9e8f0986e17a927c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c21b9eeaf320917490b3f7732e90c950f41cb742598fec7108a539e88f334515a7dd71d317efa11d7216b739c621065bc782b33d05df5aa49c19fe45c294a077e3695a6e5aa983fc45bb96c6f931f32cfe929e2309321fb05f50599ab97e3702e66f660da33a5d66fcfd34bda010426b71fbd56a25134aab24fd73ef34aaacd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd096931f1cd4b265532130b2dc4c6fe4a8fe0b40fe2326cf7647761fc214bc6807d6bf86750c12b094ef486b4b865760b47027ec1174dac2fb8622006bc2099b043f924223aacbe532292b117f4dde5b2206996d54ce597d386e23514ba96bca5e9da98a77f88399d7c840a6a2f8b5d8a4b3e772d44394d6a27b69559934493;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bdc93311f516c83c403f72b5a8609295d0a52044dd0d38e504a07639fa51e199191cbfd6d428e20bf49f375bc404de2dc86f8b5b1f91ff9044d46789c5289b08ba7986bc2352c9d115c871d7debd2b43f7bdd272b08a69ffc38bd7434a666880e77858d0d890b4801d3c798f455df555d1b57331b038d50f6d40fdcc48cc0e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fd54ef269bd545bf89a59f111b677904438b26a9a6223a09b43358f9a1f177c04f577ebefd7047cb5f4f13c56f22498993a5ae9946125a7cd0101122dc9e961b83b4ae19c4ddc8e45abe1822bcb9f72653dba596eb5ed2e8003897cd6b9214f0c2e249053d362fbe132541074034621aa7bde1b9591dc05130ef04a728caf99;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3956a0b5b66738e269f2f147d068071152ce2daf9327ee7a41fb3d630a04a384939ee6dbb0756435779a7e22d572417098f67e3386fc7a34836c06f821e942f23b45a7d954958ea4c7d65353597c88ceec79ee0e946b6d019995fee12b8c1dfef174e65fd8c646461fa09c1b35e03f844ce1011782afce47d1550eedc546740;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h203ab4cde02a779ecfe40d0fd08e37acec0d8eb7a4236997dd899658888c1a7766fa884afabb3b0d101c728b7c28d05cfa7a184a3fb2ad2c8c92d93fc1c70b0cd82b51b61d29f13ddb00a271bb5fe6687eb0d24d58e2181136bd7484a43d6105dbd5f127c9127527da36ac048f083f09bcd20ae84e5f7f960ef33f4b88dbba6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32a3bf9d8b0d7511b707c56a657f267222f785dc816cf7903d639dac28c0a13080f4632d83a36e8196e34288c4a3de69d4d17fade0878d23c45c4b46cbef57bb01760ee23c3ec6f0a9b23ee453c66e3787f0eec76e2885200d123a7c760673e4f3fedc95e99ba1e0d845f13da10b86c803ab5a2b9cb114a6abca94af22812f38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf92e0ff6a9080c90a510bcc1fe3af67d24c7179ea15a70d4735e52669e241937df96108471378ce5766fc8b53d6b3bd02005dffd82243a2c2a038cfb65f1545794694574e1e5d5914babc91c18ccc131af243454298efed7a8f2df6e4e6c07a886910d5d10a9da50f46b2ec4a596624316017456bfdbb8dd40ae2a7bbb1684d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6920a68f25df967bba60ba8e369d1e4fe6af37359b6ee83594752c3ab090f42fcb74a036c332d6b4520226cb07972eb2511bf1da3e05eed64cd01a28568a6f4abae3f6f984e4bdff9abef5bbefd9088e7891937ac37ce989e5fcb01b023ef9c1d5d3c4cce6d3e0f0cbf02d2478755b695ab2312fb9485651c553adc95670491e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88e6d15ebfd02bb2f045e122128adab8bbdf41a825a2afa6319ac929d31ecded7a7d6e4cda4c9bc43d78f81cbf6065dc5d7de70dc65eb050e52da6fc848d4f2a4c3999327141be0cc4bd4e1af78b185b82ccd4025a45fcf147fadadeb1620ad5d9e81f1e0f0cefceeb4a071fc3f7d81bd10dde69d7475f961f1fe3c4176e1be4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d91c2c393de4d0052ee0f8bdaf1b0c430447f01b0111ff2337e7f510847471746967e25f607bb16a13603ee50ff34290d5c93934c0b8a648106b499ec64b1f6b3c0656479413709a66332dd46e82a896b4a1469bf241810329eb1456216cb2bf03cb5a98df243cf4855fb3d6a9fb1d11950b55fb85379b5b76a18a0d15c31f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e27f41563ef30f078282c477aa4de0cb147c6846dbd91ee3ac1fc9bef94ead7adecb66baa7fa4d8806cd147d3ee04546fe9d5e60ecaf6c9a07216c1fe2b6750202ee4cbfc9a4f86598ec890cad7753f95ea2a0cf4b6fde0d24d6b6d0c96b5edf42eb8d81e2b2b8a1fdc67537a7fad75955198808763711a7512b4c7107dff67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf839f19dabd30da3fd5caae5993fda23d9f6bd0021aa92cb717a73923eb0b5934c9305a163b2e5928702bb7029786023110216eaa5e370eec17374c3be3b66271e3ec9455ea98e2af1b843f1089db709820a95162c136761627d13367c724ec6c96b3608974deae3e837081b4bf59f707176cf59e6267de0510e168ef79b1d08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b402d4ccbe0ad13c6c63211d30b1d07956158490f0fa5865fc277d0e66b17cd9d82ab915b1923380befb0feee6d5aa6aef916bab5dc4c7c93209211dfd2ef163c722f325a9ae9b82c095d98b95b22fc31c7b5df49731ef9c2d268ead41b15b60f86cc34118bcc6d907aab09860f1a76c80aa4e1854b53d4d2dea6d0ed3c1798;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cd5c168c785324938f964838cbe5e8d5360ff1e4b89717dfc13d63111bf97bfa3a013045c8b7aa70446a5ddb2bebb710c1bd6bda3f9a28c4c0f34f6062be90be6b8edd4134153a9ac5ca921e9e3ebd423efef87eda8f277de309a243a649bd692ab175778f3c88e4e6f714c655c20a1d8b4866e33dd2e9b6bfaf293f4d63921;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5c6ab5b4a4f191f8135a2fd915498d909a3691d9b5655befcd8ceb3cd1a787fe66766c0fe8e440f9bea2effd0edbe860951ab9ec016c09fdaba0daa4883e02e04f736a8db003209423593825cdde1cccb9c5699d0b197df7d3a0eb4748281c27f97dcd7e3bbb333190c80a3cddba0ec3cba9202d4d5aef705d934fd849c954c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha68158cc5fac445a616b80f004c826eb7a4bbf505e54fe52c498a5a6efa80433fb4a177cb59a2784c0141315e5e2cd3a6700eeb3d7d758a6c655061aecef4e4692dee1b25312f893a6355db7dead788ff76f5dcbc0129b483abd4eae8dc74b9b19d720a81e3ed76b8625d9861bce059c6933db61d625261fb7c0c2ba7de96fdb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf216a30f2ab14b16c093b9fe047bb4d2a03be9136548b0b8da231b6d44537883f1546b2736dd0cf09d8486bcbbd9f135e4bf3379fc7ebaf8f1cb6bd588f0e16398525792d3e71276e5c9ed5ea96047c2b39a656a5cef92c8741bb84c4e4c08672eab386dfefe1714ab20b0d5e244bca84c6f4cb8966fea2cf9634d5c845a7d83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44ab22d6b6eaf9fb23d1bddaf9729e2ce696ebb90f0e38cbff50ffc1606be7a9cd3fd37b43da043b0f25abfc9e4daf459d0ad424a890e9dc6334b000397c40d8a1c21a824e8ef460f4252357a47df73556319fb178d36944ab56c7299862760656f186289131082572914e57ac2ebc6faeba0ebd51709376a4b12980119042e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h100c0763c33c41fc12386cbe436fc9e59d6c70cdb1313115c4904df4369790344592b74fa163b5428ca06629bebd81ace514c61b4216d79a1344779c54b8767e6a16b969f8be371e5f1ef6c3507fb5a698e95d0d8f7748c71d2832b18a936d77869485e083b98812777c0e15f9e657e465dc171b5ff466075ff6584db8d24559;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cf260725d3b12052eaed2fbd937e7024f769ca34b020d51191b054aa722bbf0c66faca1b2725d4ad3e25c00070ab826e8c527f1144429f88cc008c61e82d74ee47d5db6e909562e2ce56b8e1ddbe75c8f1d2bdffd39de3d7447e04a23797498f954a7b28b942b4bb3ca74864fd05d31330f5bd3bf92828a280cb410a65b9524;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66722e02c72c6b972b3470027c3b85669784ba18578792b1e040e6da615f135f228cde985cdf0973c798da2decb1b3e7e58917f05513e221ddd768c0a57ad29f33e23f4eca07730c098d029611bc507482f64c6cc6fd0657bb9828102901b946557fff82f3ff543c3254844f61c3c4cbb35c52a262536779fa26eb32efeba779;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8211dc3d965f7bd3898e918d5ed77fd3e30e9fdcf7f034f7ff121c82f8320d71185135946c686dddad0d15f804c5330edad4b7b97475163db5264d9e61a6c7d15f351c0d254dee93edffb08dfa6dfaaa0c641a279a055f5136c9c8a987915dc2d4acb2949bec2a85085f1e030361471922ed9b02d57cb24297825a9ba42571e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31985e55b1700f0eb592c9c3693b0fbb65d1f71b1c72aa64082ed0f58462babdf7aa63160d36cf1bc87b02271fad40fb897b703d91c2d03c6d2d7dd57491d8ce5a1acc4b024182d27a7f45a47a9b636eaf002ea7526042a033e3f2c9d34409121ee86386debde1049d77106b9152ee95d720d34e0f1155896dfedb483fa65b9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6be4f3ef351d60fb32a3ab08c234c4d17d638f4ea13ae9267779c8c2d334c7c9554b6209c9a0aebc7fa6625eb19483420ec13994f524a855cf3fd1ffa3ec2fbe06e92988ed5b7d423ada64f3faedeeba634f80fc954e56a5f9b1c0dbb8636d5bf0f270406d47c07897bf889f56dc4bdb28c1967dafb5602915b9770a3037d0c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h990d8608c6dab56fe0ab5f77ce4fbf4c07157efa5145b432113cafd5539a14905411b2d4714b330f9a02a8439ca60a101ae92d2fc37472c36124dbb993102df3c6feeeab24010e836e691cb965a486a4440e3d23c8e384baac4102f912400fb52d31c3edee7bdcf072e87be42e955bcc89f8e99d0f2e45e97d4751b27ccf9f65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10866f6d1bb186e147be4848445b0884defb73f43dcade5890303f6912665df2575a6d753d158071ef99d00d46b3cef49078588f1f99ade44cc1ed55a3d2518a97c76fa46564d3b4da6c3e8caf5128d2884547baf82b433139e287649c568a15c94719aa7ba13fa1087c9a2f0d58f86f10c66578b2d7f8c5bd3d40980a03fb06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefe954b5526cf389a1fd195130ee82166d55f474d402e8097814e7fc8b170d99428fad798d6bf577b5288fe8b6d78f281695b1215c15ced3d0e02b4cc8c117606f1746c00a8ae04aa6fe842ded21b0fbd3b334edef3ff2f6e56b4ddf95254d305950cde27aec36738adccdc15dcb532d57d9295b7d30bec3a6357fdbc8778cee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd65dd448f90e61ece1adcfaf925a604153c9a7777f9a592cfd62ea6330ec8b2b7e2451874303989b04e56cce7b071b819863d0fa8a09d3258775446cd53bcdb672009cd3a670caf05af97f6ee2633a8c30d4d53a3c2fcea23739e0685f4951c123bc6cc9e85dbdc00722aaf0b8d24a4b2a313dd7e4bc6bbfc106dab02064baaf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd09207fbe42602da4a1bd60a5069f5a830729de01107daf8b2bd0dac9cc5329fe0e32b09c1df18d96cb1f5fc5e71a4f36d334186e790d8d691af53f2654010cb269d020104af8b80fb2a6d5599d509c150e3eed5a09e0c85a7a3612df0e844626b21deb668899e5136fafae0a133dbaf265c6dfc24f1402685d4f39297236713;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a40279a5dd7f456c5fdcfce535cfcbd33ae877a61f509dd998564e4f1cc077e7a356a498fe941a659ca9632e2d3fbc072c4a14630ce612c3b1f0a3b5b897abec7d72324bd0a5226f75e2c1b54fe44cd28d063a8fe480b27a7cfc641727980708cf90eb6e6eb2441f7e22d2c3402b18eed1c072a214717ee07c7d22691e5bfd3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d049fd09cbf8946344d9e2d64ad7dbb3184ffd654343f430357b8b68a7241a96f661b7fbbd1cdf4fcc9a253a2bdb29159f9447bffbf9999ec55049e5a6f157897984304c92808461f3d9d4c320531277dc214ed1dffbd9f205740452cf4c393e3ec6ba23398eec8ccb684851045cb17a7091405416f8c7c88b7fb1b2fda0f9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b0609f0a91cce964d021ce9d7f2b2ea99bdc8df5c0ed4de757a8ef576780aaf0050c4f537d61c11e3dd18f067008280a0a7620e0555f5bbd85bf3ffd493cf9be09575eec8b8131ed51460d98ae31f7e003e48616538293be8489fe30c5d15c7a9562082091358dfdf504676e3aa5735e136f0b62d0ca397843273c856f1d9d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a2615625e99969800b89248431c1cbbd854cb3bdc8a45cdfd88d260df6d5d5c20381edb9afc8b2226853c518b0473eff7dd71fc3581e46942957f1a7c99e4d90ffe68b0a10e5473a8355f559d3a92d8efbec5b8b5468d8fb7277a8a462a22ae8010ab362fd74932833446199d1347bfcea4e9102742ce4ed751e0be9d8a50e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf11b0c3d346466500d8ee4ccbff5ae72cdd0e7d22e06d5e6e7b052bb202449d0ee590b772eb75f2ccaa516261dd219ec0e74fe75189dfd3268de346b1a41fa9d57c6469adb0a213d3bf5c0fe508d2dd12dffe5f3815435a87322b8636618c54395f07edff0f0adbedf31c3557afd188b0ab1b722a1c7370854c0e1ebeabc021e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had8c1acaf20eb95aee0c0efa14b780d47aec803c8121d9da2ac0591fe70bd80290fb03b2b112638b5d8d20dd33fe02c26ee99a7b47dc3b8132a98723a09be898e7adf6283e6aeb0c317585e3daff453739d4c1e279071f7673d2534b10568a321eec22c5ece856852155e7f05fd89312362c6b27d672cfd594ad72b706109737;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haadd93644e7dfff0340402d76a35604ba0d72be9b67681334765a43b36476ade8f9b39767eb04e21eddf816910263ebdeb4bd3efdd8768e4b28824d4ddcc2540097d3ffd7bcd063c0af987b512f886f2a72b3b346db3b1520b7ec8649ece1d6676a73caee36dc3af9a613d38b7e3e77913e9a9e3e2c70c533e35f2877b4e0020;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8af25b48ddb4a6d46ed12e37a195e88402e001453c91263192a0dbde4a10521bba28ac144addc3290f94260eeeb3b6cd2c95a3eb2caff005b869a7e4c7989198e6347b487104c41cb24a59afc68d644a59dab6e36e2b0b59022969437a26c7e97e0189f6109a0ebbcd3e48e13c19a5cc826edcc0dc0a8c67849458b4082e810;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbab3f4dc2bdeb6b1142fdb06b7402f4dfc25c7d7b7a2cbeeff0f631a85bc4882326b82cd63081cfa4ddc2688ca09b6e34e6e822f58360101480dbeb5b0f954deb2cb5311edc5fadc68c75cd928a1f210615cb6a2b988b29caf05245c019d4d3ae280dd30bc90ab801f0c86c2dc2bf9d0c97b384c82333ad129caea600bf6f2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefe546a4cb2493fd21f537eb6e2a37cdda7b509720141fb50ede19d71fff49b7919f1998b118182faa109f97ac568482c9764ff65f2c79b5eeda57d859f732a77d09f53b554bc2446d682faf8fb6bc13ebdf00dac8092f788f3f2931cf91a5cc897a172f6a2be184419b6ed46bff2cf909964c49b3647e969c4bf5e1b77d9720;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d9b8966f9ff1b4a9df3b2fcc637fea8bc57e9a97bc9d8ddd495ebcc21a6f5acdec9bf713d4b140b4793b47564564d7d4facd7dbbc658538c7c17bb6773bc337f196d38706c0e90eb0fecc3a95be85801e9769794bc55d9d953cbe7ae8f27f17eaba92f09c60318d7ca40e90ff29e1af01353f3637f1676dd64a4a101c19d702;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h288fc807454b2d14d465a9a771daa64f63f22fd2e976e542bbccf101ca61fc6042c933a95fd8f94070bb63556dd00700a234f8338ececccb63fc6d0a771056983f33bdaf8e879bdd63b65931bf6e0b8236dc729ef8868a2a9e2b61ce012d148501cb236c5988da29897274c6383d6fac0b79ec39491929245c661fe577b69458;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb21ed5bc9dfdf829780080b03449d46e4f9484206bcbd353d6c4756f2037145cbc9f528efafb29c0c7f71af5182af3d2134b8c3889ff0cc7c2806ac69643799687411832788a954885dd87ee2fdccc1121bed2519ae4e1edae147ae5f187e584e697ac969f51f123f7260319cfc67f804d7b13aede17fe34210d74ffa3d36be4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f67dc631235c7eed7802af8ab9ad590a30b598234acaaac576765e61de8188656b539636d8b06a9cd7e52c542ca6e7fa50915696dfdab99c22c9352e97d9b6fb4ac0912be024c4a02b5f17f30def7b8fb80c486380cfd597821539b0a713589bb87743698a3ad99f8c9c082511abe73b0ca2f44a29d9bb50e3d0069b5c2355f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d2740b4fcadc07da59ca1fef008344db87ae72b9560f35ec448b48d7f3acbd40c592896fae1e8460f0cbd8322d834c9968fd10aa3a424f99cfc2cadfb04caeae1fef890f3f3932b071418f9d9a86474125f1c4a4008522343ab3d56ec41164e16680709368ebdc2e2194ce000c5d61b276f447afba3e4f09157b4e9592f82a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf8069e8aa49ef45283289070e7213542cbc31bf7666a9f5e52cc217be7d7c5d3e0bffc955d89571316b598c1407104916448a8498d0a8c6b50330547863419b86630efdd25f663c8b73af828638f20e585c521231758fe77ca8cc73d692120d25ef8103158436d97477d7f6317ad27c5cf58471ade299c3fb436029437b3a08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba7be1609d4a3c9285ee196a5f9e99bbe207423494d17f5a7ad118d792594dede52ad53cafe4c04898262da7c1419970666e95f9ed8aa4261a0cc83b4fedc766a4a47544982d0a848cd6393de91954cc5c94862ac4d7d5d19386ffba277317afd587a2b6f498791ef69ca012883f89a91b8f35566360a8575eba11659780f325;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8367860027a9bb3f185d4ba063f993dc38a9bc24d392672a7d9e3a686ebeb097d1a206fb3b44ffa557f025a827ce62a359266ffefd6888917045ee0cb60aad4a2da6e4ffdb9c1ecb63c4b90694e98e05f38f49afee620e6de1badb342ce610cf8863db71ec1c4aaa9a70319a0ef99ec0c40d0ec5c28b9352de4d372f41fee119;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26318a23b79576b96237941dbb2c644db52885ca52c8bc33046ea5ef89e45341571502df84f0c01e78089d98019e4e5120bb297b6fe72359817d3f3c6f01e62af7bce40df4d6187a184fcb0ea946332daccef0a91f49bf3fbda0687678ab594eaa831124952c845af2a60f17e0c40421c977431a23be4fde9c35779cd7e840a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28af481e43bb9bd5486bc16f105fd8b776695d9004fd607852f57483826ef00f29137b6831d040aace6cc539e92920538039232f783dc3e3b6da427959a6b45fc5405646a1d5e31c70b154a94edc4c14331145a18560f59053553338e44812696f1fd1bfed2eefcc60f8afc6f461f4a1287ad3b311a29f4de1d58f191ea1e742;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3240510d54a0fa6f96e8562e36ecb81e38a0dc09b68bf2cb4c4fe2733903926b1662cbe6981938f4a3c671dc819fb1c22a70539f4db9faef18638b4142ab35b837d1ce76aa379fb4199fd78147d96bacd63839f3e6daf6baf97711466af24c532ca32e9bf5d4b3196ac9a0761f52285749f2be0e000d930122e2f2ca7f1124e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdea3efc46254f40e0ff66bda088e9de352a9596a7029496639f61eb184f72526e46bf199f2f44f447d48fbdd25862f22d900dbe366360409b9b7a2c410914e24d19044dbb86fa98fdeef5b184e5199052b94f85fc4074c4469e2c9dbe97e5a76698fa3c8fe0a136d136d5b7080351619468b4701deb69a3385ecb0d70aa0e21a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbca6324668d8ae77a6a5471694730f6f4f1e0dfaae8085b53483bc7db6444fd69236f7c5c6a93140aef21e07fbd933b72690df8a4fb905cfb2b7e766b1292e46bbd189f33985a6049238bdec13a14403e5ff62e83efcc9ccbd83af028f16b5f92885187e559d6aa63f423f93fa1954c30f503dd2afb4c7764601aff4ea822b9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75a5e97391bb61577afc4b5aadae0a43c9bbb8f04ab52155e30642854620f5b4b245e5e1826838f527f5ec28260743635321cd42a5b46bd442cd4160d30685142e61792250c8922b0bbb1a6ff3f3fd8e353aa0581b340fd2e7591040d52cafbf13bd2825a8ff17744148d88844393558a9455edaee8f3a0a66c02afea4ee5b02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a0681918f9163bc0a0368e945be409d554ac9c13b3b4cc83dc393dd75c9927e8b56634e4d74ea5119d377a0238b0b0a84143a48ed5cf7b8a0b0038132253c23917dd7274cb8d2706f7cc745260fd222ab43d16e338f499e28d1ae37ba8f592b5d9e9ed7088280348b2bc67a912dcc678dea493f8bf4285d86957df720c6ba9d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9109845aef55601e7cb90bd9a9254c1f8c99006d025d44369d85a2e65befb85b7d377c7955dcf7e95b3c929de7b1b2ff08b591d500edca68e96aa772aa3ada558ab770a354dddbfc12b87a4766c60bd47eee493943e291d1a337608e49b94aa4f066573c3c83e582dc88e640842b6c8ab6ac3e9cc1f0ba975815ec87ecb63d92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb769bc8a9a264855b3efd866322e4f936c62bafd22c3c9359405c3e3feb3e5355dac8a6050e91a9b02f0b4b462d0079cdc9309e1bd092026acc6ba7a1af402eb32a220e2d7733fea1855bef5b23b844049044ce7fd3f23ad0c9d2186d7c1c4ba263e70791d9cdcc99cf1e5a9afc887931f18b9f795775cd1203409d616c35c97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3704ad64d270135227b564b96d21e40f9cd9fba9de1f22fd7d039bba07f22566326379c7c2046ad9f30dc00e95295115674300c68e9e60e8017554d9ae6cf7d78889fa4d655e8ba9d60244aa1c77445ad1eccb25769550b10baa1b8855019580c3dccd1eb56a6170137243ee1924c46deb3e5d93e4cdd6c5eb84f8c75643f09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h575672030bce06dbefe35eb1fa1d61b4c8e09f31d690d9c0326ccd84499c2056cb40cd82ab82d87b3cbe1dbdd09a9d50db550e337e70c1551f8bb1e6148de68dcdb2d67ff6a9e8e56b5b2d22f238d1c0d80be7fad197fac1484f7ad9a2ef8ed857b9650a828473dad64d03fa2fc12d30851321fb5bb14024d020db2e0a1f8e4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a72907a945b88f9db2f8beba0c74b112fa672c1f182ae6c4e383a630c1c65bbc7422e6f385704ce84df677949143ba59fb53385b5b096921bf8417231a43845e41321d492ea786a3bc66d8684c9331b69e2ca8d7ea0f045ee9b2ef8546baf19e64511db71fd7b646f32fdde04fc72a24192dcc8f6099f092339e1d46fe655cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f502bfef7d2f2600b96d10a9e8a5fd7eedbf7d246c267fa8f1d30b62a736b570b7c19235b7d48d3f6f9d149556ba15173699a45dc54440833e6ae7571c039ec9c2c62f8971666b8e2b5b896d7ff117b063549e982c6e1a2491456dcf0a3f4122bac411b0038454af34025023161bd05c443bfc8220cc50315f8c4a340c477ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c685aab68fe43c51eb876bdc19334422543d9ff9ac58c6d478eec836ecf2d89003db9976e852f36b074e63b3e50a4166f853020f2defcea7ec5a4eb70208960cf89c0a7c30c549bcac174879270df516a9732ca994cb1d84459a4cf9ec05e2cd3af66a6f546d704356d095001b5191f32cd632088e71986b73ef4ea94b9644;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1e64666998f5217f515662b205fe5bf951d2b3ddb4bcc212b72df527b1b27810a17b7c72d6c5a5e99a61152b8ff32fb916d14933284ae3ee832f5e3bbc2da1ee7d40d610490a164fee4bd4ac3215696912b329310fff829d2b3724865aef368b7454756d57bedd225c7b11ff0991e767efcb311eaa4479ba8696b0a57f79a63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b5b234ff47b93231c3e10a6dff30a29c8dc565c519da21de7f722261e903c105bac8f0c987b84a753b7c46bb639342c3256ab929dafcd0edaaf020610fdb02e106f9c36e35eae353b756031a9aa13ec6847971c6bba217295261f776b5b618f200f1eb4506d9ab94adf23ebe2eaf2c3f8e9b095aacf7684ad4f48e522a5fc9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1e23bf3726bd10afd34d183097c2659709ec8645c5f2fca57b9f903a2d9456f171c1814523109234cd971ff2b189d78388c8120bf9027fe5cd9b9e23e8cfe8568f1c75a5820fd18b331e31e0fc7ac1dc1b3246e242294fe422acee48d9d1711ea6f86b2f0e93592e6838928fdc204b7e2161a1d97ea908af70e5890172fb57a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf49c08955ede98158cc10cbf953b9e004e7016e011504188082f0223b6adc9d8e02a94666134df765e29d97f7b070c604fe942258fe6224cbdf14ae118113eaee67c5ed30484205a477ef3d0420c068c27bd3ac4cf3c67ce43b86205080b6811afc8da36d15d979817eed892c7437acde2dcc2dfe940864c348c25b80a785b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66f45ef4b6a2395d573da32f501448b86102e744de11932a574e5e28b89e1845bcd905a330c90ceb11b898fac7c2b46e05bd18b81fe01d85ef347d9377c0940ac4aa9c7233dc40483b6821908d79b51971b5630e961d06531ba8dbd7f084a867b2250a879b2625be09a582ecf922b8278882cd683e8d695310014237fa1418e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47e770afde9e287040c9befd43482739b00f5425957f35cc90637d00984b117263007ca1d57c69f185f20ffd3ffc3cc79b0083598c991255794930eb9e0431b307cc2c5bc9fd7997ee644693605b6e9e1edca64b703c3ff8f745917998e639bdc4b57fe4232bae7450dbb43a1a625f12ad1bd4b63077cc2bf5b779649d133694;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ad0e0f09035b3c0378a83e7a05ed1de9fabeda71a2807932ef6ac5fa023267ca6387343bf902217f267c7f353c85ef8f9f87e1bfdc8ad8cc124ad54ecbfe3bba93e2e8d39d5d903e3ea37e8c0eaa630d5e74b9bf4aa8788d385ddfd25327732d800c2447eab3ca6f0bf12a7419787b4b8f665d9dbed1d376baa1793d39ea297;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h758ac0bb5acca4023fa71376ca77a89544d7cef3b24a73fd556227bc096d6d8ffc96447540dfa4b7551f981a711e51d88947ca6978786fb84415a1c29523dd923f36a1371d0c878b43339162a5eb1270db7792073bc43f80e94063345560fa34522f6f2b132b8216f762b11e79dcbb81920b3ad19d0cd8bfea6dbaa4e7e756b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18369c2245ed9bf8081894879a4b7817998d9e267fd3b37c0b1dbc18d254f1597ca57613ae6b252944895d028c554123624f29f54c8cdc87b04172be2efe918f35079c25ad660bbad3c9a4b2c3b429ec0ebf396012aa2ab7316cec9c57e98ef0502e6bd20c079dd975c2060b75176d47258f28fa99252c4771c0df9aec73a538;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c2e7ede6800f2e441a7f293dc4bb5f6123632b367b35c8df24e967fee15134b0a7c7fdcc821f8899fcfaee6de4e84c76355f831f8cd84bf6be1bbbd1b431c592644d4ba25d1bed221f2e0b5bdad016339bcd4f2920e84aec8ae692eb65b5750af857c968b0e8510061e2b56b743052f23b353282974a6b27a5691fa8a116b17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64fb9b086e80fde024c73ee0a1063c123e2c6fb4fe4ff5289d280a239e4d4ddaba0e0477f6a04cff3ca8f2188505fde69e997e0db37172720ea41b05edfbc00e5d47074ab3377728b498ada0646ddd5961bbf7ed16b509cf60c022b8797fecb5815fead7028cbb6bab2d17f71ee3fbef54f4a4e2c3f3ad779476d6ff78f51fbe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62e6ae0dc5d2bda36a8198ffdbd1059766b61a5ce0321300837ffed577bd1e2c514f6363d8959361fb36fb778355cf7d825df5bedfe989a0d0b10b0785dc4af0f53af9aa3ecffbc42f1c428d4da58cab17529650de7a716bc3833b59e82dad2b966c422b9d3707a05e7cfbf94b55cd6bbe510f0fa3e1d5727f05cd4ac7969da2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e25b7b4ee9ae3c482bb409cfecb06c9434cd91800199dbfca09923a4fe9bb28a828798431158e535f4cd031cddbf50befeec2cb05b44ebb5f4230bac86977632461341ca7f4036e59867e6043d767f1c96b74db23ff0383b83ff96add79d4bcc627cc37960e3a3d889fc13e64cad99bc57ddc0112d6335fe011e27d78e0c184;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc487272e0ef811990f7c20550872c30cd9962c4682811be23f79f45e2e7e0d5d68b0c4164d446c6dcfa6cbdb666fc49665ab2b0e380f67a6a67719e2d18f09cabf71e455a7b5949fe84e74d6d981cf9ea45aacabde01c2a16106746a27599a29335949421e00e606dd1c97ee3ca2809fac155b87e7d91eec2a8aba9f74125da6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42635c70e6a5407c855b40fbfa0229d98f0184cabfd172db4e5500df302db6466a70cea0e75e15c3b03e83a8b4bf8cbba7bf06e3e3799bb04bd49eb6681bab77205a1afbc1919552dac99f8a067995a540e6d1e9b60fd8aadffd876c679e9eacb3e2f3c68e88851eebd2420a4fd5d8697297a0f90730e5e2d12e10d7a451215e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he222e19a57c3ee13416001d3e61a5ebbae8e4df866a8aab51813617096b888e1c9f7d35f9290eb43807637edf1dfee233528255a64358ad82b8df3c5d2653c365e93130563b660bead324bb197844052c3183ad6af31155e0385cd79d20c5776a03ed96e4511f8dce9742b233b8669a280e8b0cb8c4a425dc5361ad0389cf1ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ff148bca945bc790ff72300425e2a6dfe615fcde3de797b8bd620d9d1c21411d7697241208cb2aebf343bc8eac8ed519714d92e4027ec97ac66083fe658ae0602a5b019019da26f667ddeb5691a53ecb3f2694ebd3f55c6fa05d128010946dd0d62ae2755160b178af65243f0672c76434b0a9e0632693c7251d38e10d8dc97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6207fe2531b9ee037b2cbd7b8d6d89f3a682866b372ed041f04d4ea50ca74ae91a50c0447dff01543ec12f62aa1e1b561993f0290389c2c7cbd229da5b978f67301a5768032469c24e089ae3db0c1b5506f9298f2cbe2a499d412777973367242875a9d7771207b25cbe5a6cd8b0752330df2a121c72cbd0042e1441c0db9ab7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc889b98487f8a0d5a6d20955377434359312a95c9254a3268bb7a53d4b795f83131f17ce5bdff890a92c5e2b83e79a777cc9508930d46aa4de425d7852ff79861851fee1dd90828a9d9b14afd1e8b86a66e81ac8695cd4cc3ac9862dbe0456f3c465f5d7feb95868070cc0480e4eb84a9e0eaa5d12fdc69a695bcd2fe9a3e97e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68df27fe8de835dd6e8b9ddcbca3de8017d8122d93e2d72a8fe3f29b618e8f76a31e4a9d50eb998752e1ebf688e247aa575b8a809493215d9b153936e2cec1ef53d786f9111fc5733c6055812c3ab570869d22ec0b137dc384a7017bb0a3606f344ff740a53be2e721751aea43c10b09ff5fc17815dcfe22635fab549e241a19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90c2f4eb8ef5fb1df959923307b11e6595f553cdca5ae69d746f59bf64eee3f9e692803a47b86b77c3dcc98bedff61d2cafab48e89a21e32ff7fca28246414d1e1514bc93a1cbf2a891a026943246dc2d65bd4766c28ff0b9b2fb9677af158a38e31561d9c0c75dbc3f67227a8dba4f5cd1a8842954f537b547f4c0079481653;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7030a63ec4fc077b6b20381d9ff21cdf77d10bc8c1f3a6163da61466baa94155866c3e3fde34e5f9afa7fd4ab366f5aaa2990089023574a462c5503fbedf1d46a2c9a0c8fed33f6c75d9fa395da574470d706a66deb941d7bd5954e086805c1908019a5f995c127d536a0278e41c1fadbd7d2520dd19934389e45771467b5f1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bbe9b9a4b0194d0a9e3dc43a9404bd796afe52297db966097c43ec30abc78906accdfcc755c078377772204c8a98258d2823ba2486774de796696ef41275cb8fa5664821f8c9f304e3f6c26889756eeaa3e3293300ac5df2f447c764e8cd3c4dc88e02845f5d5b3a26b8a04ba900e596d6f34b1a9b57108151d9786515d9986;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3c64c254b76934b4b6250b5f4d39f873c05306706bae8c46183813a3669c883874dce86fab78c7c30d4a1d0380f441266de11c33b615a0c33c782b7ec5d79718ae33301a071177a5bb6e8d846f3fdc52d724296244b2533a3365cc85c6e0095a31b6143a21d3f6efc14ef80d15d402573c8b76709e708d3d7e5f8c8bed3f8e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h426c9f654390612da0bec9403f6b00f2d142fa0fc1a8434b4f3847fc8a405a083af3bfc2e27703ddf7a839189c026c50bd62577087c938d2623fc0cb8255d635ce06f0ca244efca46ad59c0b70f92ca43bb04ca5431db9244917e12a54278070181eef9705dbf7746eceb72af5266ac43d73c524bfd9045a0129671207f3360d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4e0c234c65aeb6c16c41bc349a94d713bc5f87fbd08ceb7dae19f8b96e761ded92030f33f8f064da87a83311a737440c7662393672a6851007d18ff96c0c3ae94007cf16af8d2c83e4fd9c7d47bb6c9e444ee487a5fee5b580df598b9f7412c9292120bc0bc62e96ca6085c946c16b9d1788b397d8e8be87d2418843e0fbc6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69bcbc13875fe209905e4c78dbb1f8f30595fd733e757c9332b785e584f89f365f10c6491f281da741d832560cea0d24e57fe91d8063556830388458a7420b9eefd85678715f35915c657aa0fa418c8c702755a7654b6722858bd77caed7bd3ea6e917116b9c2628fcdc8e8b364013449a8f1afd54474c45fc017edac8585db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h891516c30025bd1ad410f04f487088a1838ab215d8cf146a3c2b140a15b71376deeca9d240ecbdd50cfa49b6d978e244731d97a00dbfb3100235c1059030575d6e0ccfae8b15b20711c3995da5abd25c589c16897db8ff80a856b0ad2d24da935b1f6b9d7bac068483e004ed3de27b20a0e7a3f769ed2c38f7405eb14e5910e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25fb04d9155ccdc2b77cbd2e8501b462109ace82edb2fb8246ff2d665acb2d3f0647319b3a6189bf07db157da4c202d87f480876c661d47d89722430d41bcae5596640ae086ff9cf37031108d14a1b8b12cd09a968973dced04bd6c9b4f61bc3bf10744b67558dfe2e1749b7225d57898831d9b2e8e2709736168d60d68b583a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f01167ad0548d49c74048461056ae6fcb8d39cdce709d3e830bc587f3df93c78730bcc4462e6456723824fbcbf4751321610abd92586bec65abfe0915c08b10a075ede22044562cfca9b7e02601af51450c0ab5549b54fd3350080de47af19351562e0187dada201443f36d83c6125dd46925652da23ab6c583be28e1cf8162;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a762e3e50e4e54ba3f4966ea8904d8abde9cb6199b78183cdb2f98ddec2d3dfbbad9c4e51388dabe41d9b18cbe803ce0e1aa36fa40a8343bf4baab56b1511907cffdc42cdb738a5c9e9981898d8ac049f2f216e15e8a01fc67230ba057078dbbdc69cedae2f3248da844feb83beb954e4e117e7e6b41721830e020bab84c71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha15da3142afbf86888c2f14fda4d180e07e6fb2915a7724b090089b01c11b20265560fc18d3d63b3a71b4e23c21cc5c91ac660f491440040fe0ad170efebee51c116b3d05bd3fe5588ef1a06059d204cbf11229bf10084a7c46083ebfcac0d192c4c4ce67f619986a7fe72daa335d861bf58a35c22f1ae6b225a2f6cff643a4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c4239228d84628551d9314b15aea1dc0c5e7a6fdf462bb017d945ca989dde65b295d1cf25b0fcba3b347e4f4cb20ef3f7f75c74d2ab89f74d8ea9fdfa8b29a2dee082a876a103e48bafefc1908cffb85465a59b7aa3f66a8b5d6ebdb94244dff781ddb917003185d10d3c5d60368b844c1ed9d301d1460eba1f8d1c64708b3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0da91766b1174b821ef9afdfbd70c69bd9a769d3ec4a372826ce692b5b7f72b7a9c15a42631d3ead581dcc3b431fd2627cac6a84d1d72b3e19a8230587c6edbb3f2618b3dc5e8abe649e3c33edeec8d2b24f343f97e4b7f76c5bc428289899220166eb229e4df579d6478c56fd68d134d75ca3cd2b0b6a3e75d13415111576d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4888734cc31512028c8756d56fad7d943111b19d83b047422857417a967841dd4da5f4c562e3c75a0e4fe24e06ec67dde237ed00aaaa0ea8c3ef75f5976beb527dbe3110d664f15a7e8fcc5081e0a8f041d095aa6e166b2a708342eddb9939a9369f3db92267a7638a180ffc9b474e38e5d4301db551e176e131a860f0c3950;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c145bdfd769e9bae554b0d674c45719cab11835748c6644223dbd69217d8074284dddd891d42f701c97e72f7a76356e3739ef0fe36179aabbdd3e135ecbd3d9af66c6041a076268b6782d226887406f28a6b250724b13e944f20236988eb3126fda97ad9f7cac7fa26297cdaa1718d6d973317350b5bc9a836c3a4a23f8d27a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d556a8f5c682e7008cab1f013568ed525b6c6a7c37de4ea481847ac1de075fa24920464863728228764ff19012fa089f047952fd9831638bfc9165ce56e52b572376fa4b5a07c2afa1fd15cdaf7d6d8ac42f0781980cc12e48c91edeb6bbcb269841f75f874d7835bef031d02c860a604d858e55f69f70302816876ca245f0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h723798ad43ee5358e41b314e609fed074fd3f457b24cdf3df7e8fef0294505e13ceea0bfe3c3e2179631197f4cc37720ccf541e2972e30a3c8bef769db1b76fa7f00a0aa9f88aa89dcd32ff3c1bf6f5bcec4a272de291fb854612197b17839769df6b737d30e49d9aaa960c01e445772ccc107e656de402611cbe1fd313d18e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84c4cfe74eadd8ea51a615a334ecf0f8b08bb7bfb40ff562863ea9554a8f71b1146f0becc6ec652819acdf2c8bd98b6038179c0f8b7d3244ee9e8a8c28858dc8fce42a6c7af2b173f44847e55fbadae111cfcf59e9826fb14fc48827aa6225d54923b57787c2e7bcf022b680efc09a08e51206cd610141a5f8baf058125541d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha87eeac1895e22f9450633c635a0685d0a8bc64de66c3700290229630483741c2f9efba73bd25a3692f5676ef5d457ea9f1ed8bd3b15970361e28201debe13955391f4704318fd9a8b1e47534121bfb1697922f0ee0803a0c8e0097d6878b6182d2f4c194b052d0e2676579d55591fbca83804d75845a632d494c55dd95e002c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h456515e4e2a8467eb5407e4ec0fc419ba5d0b235ce4ef28d800e4e1ab34f0c44a367eeac1fa692611fe5573561673d6b9f40437f7de1ba7a817a847ea3ca17ed442b99b77d2f420a7c129572b88285f10d6da0c0acf4de11629b06028e8b849d29116c50fb2cd8bae478535c4e484b31671fab8ae82d0bef9d5c072e7cfdf80d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcefb361311d2918e7c4935f46126e684f323c98759d9518c4657ef81e1f69a25533aefefb9a915323058fc9be82c60f186c85c394ee69d0875c109bfebf01d0c85c396b7c0978b50d386fd05b148603b552fcbdf713ef8effafa3f15ce3502c674ad2ec0d111a574473834adee3800445b50a0cef0cc0454e774e7932953a228;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff627f94ca95d2dd5b8a3d1007f62166c42c243cd2564b4c1028ce4e84fef844422f7110f944766b2a146ae2fe34635bf082a921cb2e47f32df021f7feb4b5a7640dd5544421907dec573c8e9834da1cdd3059eaefb651dc89834bd5ca2d752697a1010343b88f15ec5159213c8deef4b4d154fd8511e8d5e774f85a6f6363c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdf965002a5b3db31bba42ce82e270b9de193318be9d05b7e8e3eee405a7ae52e914fb343e37ae1cc5083210dd8ef2eeecafe79f9c949ab7579cb31659a15da5042239a7158f7427a667f41969b4bdf173c3574c9c57f9d36d59e1bb2e5a22f6f691d29f614e15ef6e685e11a5113d257a697caa1aabd6301321c9de11be2866;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2010b8acab065a4244ce129efa75b73c67f042db01b80610117a65cdd1e4cc65c2bf8e94c722ba70e5e707e7538f630967ea540a1972e6b77dbf1e208baaaa986c360132e1116c73b72088e35b4338f0af6dc60edad16594a3f1414f29b677f9f7183cf32cd9b6bdfb0411e0d0aff170f7426745c512e9ca1bdd002ea45140a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd92137a2b2ae6d19455b10f9b2bfaa6b4ac1b7d386b3071352c2a4eff9afa291f7d5dafcc93152e1130ad26861da166e72359733c272f7182f4cc0a554788b36eadbd347f98e6f7807a74ecebf2379230d7a8ebdfd00ed140d7c121e6261c76e1b979ff85e3945ab1d96602a55e45c0c433f893002e055d59a477d03e3c2a3c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2513b30210530ffa9adb2a8d1930321b78315b64d2eb90f7bb3f2c5c5eff7224fb3d3c9d36cdb5306dd3462cd46ef5a1837bc2acb7237dac8d33c902d7e45c87b54e214d2463f80ce6f03329477f02ebdb01fe0a64a1e07cce11427b36ee38d863ab43f80097c6e46c961777d8a77ff9806643783a5a556bea5fabd1cf6b324e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h367b94fe25d9a94f363a58a9e42ae1b06dddf959d0e9e75c23c6a80d292501d624ea25547cc6c9a41fe73f8d2d6b1c9c4e9b6e8bcbad82fbfdc29542a135adb9474487ff2251a6d7d41418a46db3f5f3d525a67f59aacc3df95b79fddca386d9b4a0844eacc20c87154dc6b43e1417cda8f0b525b31891abf8bd3f81201070f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h564677fc0b9406f22eb91ff08a1a0c68496ccead10773caa4c4fe20637a2d168c3f52f4691a95f1f8854977b9b2c4c51c28e5f9d75b152eab0d1c7565965ea9914e41f05e84e4b6d7001fcb7e67696179667990e1ef1f051969bdd636ebc895c095329b449974fbcf06970c63ed0b52fe558e58eaa09d882922f3cc3a97794d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82495f493f049e02a4c4cf164c86ea6efab537209d7d878b60c7afaf571cb9884703181cd64b385c5b03586150210b113e6427ebcfee236dfb59af620832d7920859bf0700fcf9b066c0fa67e527064adcb67ba530610cda9c3b4b9d8b62eefc1f9c040c9db0b6d7341590eb82a4429d7f2009bcc79d704b182b14b2e024e2fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hddd4f805d2c8ef64fb64704d645b9159df0dde9b8adcd0c3b6284af390120a3b6ebb35593734f2d6131c2078248e86dc1b22e9243bee3e77249d4821585d1499a1f7c164c429c489bc5106bd9b989bcc84dc842031da1430d523d0e6836b6e15d43d50832c458139479a6387a7b0be60701542070aede41127523b217b965b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7712ffa3d505bfcbd6cab83ea8b223753a987192df87a5b77979008da0f19e2284e165f2ad904e954fcc8615ab5c70bf07f85538fb4ac93f994eaf62ea15f2d833bce8d090ee0a645d4ff32a346ad35f00ebd215f73ae73ec13366bd1008612bffa930a35efa3e213f355ed7649bf24e558fb09cff68db6150833e57ab60b250;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56e63c63cb30803a5155798de4bfa5929cd8dafd323d29c68eb0eda3eeef6239e884bd4d29519ef0511c8e0ae1667d59b591ff2873ce26be252c610283032eb743e00c294b0e08f832d94fa4626ba51a227a11672c12c2a9a12f75e5d571b0fb13d5bfa723c367a1ff0c6c4d993acaea6f302c91a3064d71e5cc900f5337c8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h807a7ce6c514f98776d5b4f23659e4bbc18a832103e59469d4304a56cead1b4467df75cab41b4636b8f08417e707535b553ab34a3f4ee777c06232368cd3c68699b1e82ca50460b9abca7102d2a7434196473e3084ea50b8f4223f450c0acd8918211ecd60647d9089b629298e0fecab24877171e382da325d83bfc1b021e997;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5903819c77a4cc714dcaaf6a6da3f22286534e0374490fd09796703d9fbc6fbfd4b9cdc291437c220d4794a26cce170ac5013519d8942f9daf401ebe00ea3d1509375c13e26948f678670cae3b7e04cc3796b93600f25c48a565ca034c4d2623c1843103cb0effcca2d944dbdd816f5fa89aa650a497db1e4dcd5d19baafe7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0c0a55dfc7fe3754fce17001a806f3e4448185831c79edacfc9e4adf9123a7a8c7e4ce410247335a1c788ed0804d3f85dd7a25112d1436b5b68f965635aa9728c847f5e5f48cdf4c0f71cd6f5562f0e723997302dc31828e6ed2ca0682b3b0e6b1aceade77a53cf7c4f2e22120a0eb94c07457d6766345b1c64e17438d4d947;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hccb81752f85a5ddbff6e27c81f94ec9ca67300b4d67ee58bc3d055cef95236762a7e9e981aebe090d22b2f6c14856856d254fd16c146184034bd433fd19b3d2f71efcd015bffd4031e4885804ff198e3c74d294a357e46758803b5cc693baa102a2a063c1626c0877cd632261572002f0833796ea186ad5a7e16930d44027c72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heae63c2f53bf025ec5234c73708029102f9551620d43fe4fbc8cde33244d66da85cb91a8ef0643fd8f6b279146db923abfde61a45665e8121413864ba5ef9d71ce84cec74e940366f3db49604af541fbc368e424de92dd1a33585847d5aebbe03cf76c3062bf4fb2e06dafae2d253860f1070dae3e67a143a095166b9ea8f604;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc19ab55724e486db22a01ac1c2c27f3359019486a27c8151fbbfa31ab7740942bf82691328ecda0d33a0c407ac86815ce8fd4f061513d17b4e26bf137db78e11527e1e25c4ee6d2426eedee53efc7679e1bd25cb22a180022218de60783d6dc71be64195a40f704f98395396974495f4279a659530b2ee2dcae7c92583f61a8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h435a570b71df068560909bdeb7dd49c430b29fb44028a20f54864f211eeebb7293a24cc9de03548be558d03051231a50dfbe7a31d80e14e0751b000c70bec2e77ce562c938213144537559f73fc772154ab6f98f984bbc0645b95a15ff772781d41fc6e61b488df02c024a3301c6582ccdf8a16b020fdf042638c08544e13561;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c7a9f179d3f4f3062a2f15fa6f26583adf294c995ae773867f11644aa6441cfa23aaebb0703ba1675dad83b4df7985ed250731ef455af04ce7e872a271fd9ab6c407ab99591e70e3cfeb8b7d62d01a7c3fd4352afa3191869ead1fd5637226269a7217099dc40848c97518418c193129cf63b3ce66605a493232ef9cd844839;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d6c0e6e010207a4d0827e2a811c9c43a7c78f6b32c8295e8db2dff16622cb9e4c4136663b045aee6a4bf2e2c088416ef52eab982c9c7b4004db65822229e1f3ad19b30a0006ff79e526af080b520ce645c6e66ed4292057e540576b2f4a57da12fdbbdb6c5f3dcedbebb4a5ca1ab877a5b42c168ee675e83859b6f0b7dd884f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73751e36fa586a7bb5dd4c0b5b0dd0f0d02172c0999e54f75c753417d79b477c96fc4be78b2b2fc52e98fe24ee2d2945ac7ca6a5a327d52df623fe1f5f377a5b9d199821d1f7efc4d32392af4218ff495280804f754192ba58f2a45303a4d0260b82d57d57b6ea6544ddd9bf5e2744158f42c70bf50935ee0eb6432b7b8ca132;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he378974d4c9d15aab6767bf4894863ac918b101a0f97b68fe52bdbdda35fe8d38874eb53033e22b1a0db9b110a383badd8f686c6a2a1b40b0d5375a49f9c1df482be7572c0707d6343928214ede8328218ba7c421b820c73da25c3086a4f5e70c16ce6ae0acb358df78ec1104488439e2aa9cba78637c1fa13fd7b1cabf96a71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha256f6e5d8c7ac7e2c1254d04491ee9b5c3d0904b4099f09077cb6557ff0aa048a74589360dd85983b99592fc941ecd70c874d94451e6bb4b8a5322afa8d84942c56b9c76c3e8e6930041ef4a47e3482c78dc8dbb37c0fd980f926bfe4424224e54646422b447299e04f3987583a87a9101f90b813b5013325c12c2fb87fda97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1d2c45d566637db71d2d2a207b2ef2d5b9642e74e2aff3f94a1977c1dd3218b9bcd3721876d649f1ae4a2ddc81730c75f49e12568a2888449cf09aa19c4572c00846606c552bf61b5962958cfe29c5516e8acf3df57a42cc48748b738629fca1a5f9b29d888d064bbff5cc4c8ee6a751c997e2c9fc83822aa21ddfe561b3668;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd430a5330040718963072d95276d37b78a69de07a3a953135612cad8b553a6876dd700ce949368fd5203cb5c3527a45170404983066106fe17a769ed9e5e34ea99da9806062a78b14d7cbba3871aed1d04b181e9094d15770ecc86bf289f3e0e63b4d2ee233f125284876e1e7c0ef285d98dcdafa0e069c49fc0d3b30d1e13e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76dab502e2b29fa652746ed9acda4c71cf9d9a1a7eec094e47c357d1db428532821a1a0a32f3614b23d0fe9f81f17e4a1700e68a94b2ae337a5535ec72114c4ff5536e26bcf568afa96fa213687e44d43cd498ab35af94f052c1d07ae241c71488a653175e2d89d7d7f8673cee6e56cee78943a3a84eeedb1d0a96577df3823e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h677c7eb3c9b78df68a7423fad32770315f93e20104efdf196503dcd8915f907013560f851bfc16f062cb69a912bfe3f7c12d3182e3c7a3b620983fc2a47ae9a0151b0f7c39f1dda08b67d1877d6c84dab9e29867cf00bc0ecec03565137dc39dcab7ac27f6db00354abd5937fba024c5dce17b89af236330348fb6f3bc1a4ef1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he21b5258153259f3b8ad9598d6bc1f166610b5bb3e9d59c688983130905b2d7a7f26bb248cefa3779ea48d69294d1be9cfdc920063b33a0c74bc0136a6b85f71a3050ef7e2a854987edfe4914e014038928061b4312a4261763ec29771d3462d590e0a513539c77334d78140e47f20e166153d9765bc67540406464e62d5afa5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7aba10b1f44b19386b35f106c0a623dd2f184b46325f66599e331ce2464a2ca79e291c1a45040f172eb71f1743d902b4336b03c4a056c65d3ac490d596278ef71d06e172282e05e786199318ad55d2327f580b2232c1e1e6584a10c0d272f5622360214865d0fd45a0b8db0d5853855845adc534fa6a8369a5925f5f1959390c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7965e260bad59cfbf753169a10ca18f50c0891df0bcd44190207b0bd68a4d6ae8aaa432c3506a769e0a5a5bd54792fed80340e43aa507129835436a0f4b269b5b49a730389136f2c3bf0093e3e1555cc48de23b7cc7d5d287308282fa5b079004c6208ecdf5ef445a9c34315be744b84d8d72f1cc2d46544537012d148781415;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c4bbc899d02963275141eeac006bd09401511415c9ad5318ed491342825139a7d34229bbcf3412d2997f717d735f80f539258e4fb50fab01a15c4efc1c6b698b74112041f3b75339fda78f8c03fd65d1f26e74d2e31ccaf7b575b729b43aeaac131ed533a5884087dc5c4d5439284c60980a256b7d23fb0ba1d8c9654841191;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e6aaffcb419e2f4384c8da3f1db5ab79e44f47ffbc9159fd098ddfe0df6458785a3a43f4e502aac7954e3206268aab32bdc4039354f2abcdea1547d3fa31aaa0fd65cde61198f0bbf00f2e25ad18f31b9779eaa481f98ce69fff722cd92af4a01612f061dab20f766f79cbd3a6dea87d896ed92abe1dd13ceaec8d538c237b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcc61eabeab42eefb264510710429cf23cbe5dc53fd6e5842b3ea9ebe98886600795cd7d7322ae0768920385305ac1a9035562ab5cf0599b63e210c46f8e26991f0113b2fd83f1d3308a5f683e4cbac3392d7e42d352406cd280395f771a0352919c1b1559fbd750cbcb91663d84aa1695129d0a1fb0593395144dd440fefa5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb684ad8a82d3e9e60fdfb0c0d838d9106ac56cc2cad5fec779437ea74463d0834ef808edbfc6b8190c79f626407a1af07f3bf6bd085b1e0a0662479e73250758072a2b5023af6144b595244d6eacf97d99f88eec36ad06f14fdea3dd8c03c478d065342b4bbb717285548a82b2948bfc44df807176ec7a2be90aa89066869d30;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6ec0894406ba9407ba3b17afda50f118b40651559eea7a5c741dddeaac7f454ab07b067e10332a51a32125a11cb359f26d6f796c9adba1d6025a0213df8521d8f6bc1fc124203e678a0ed84a364baaf96f97a7971c3266f166c606493bb356233dba1ae77ab2e3334d4f3aa5a15aa89e3bb14bd4358f30187801874f01975cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h689ac5c6cb7c8e0f7fccc75d04cc7239a763a8f1e1276624117adf6b685fbae2d0c23f84c32e6302b004b81247b4d3b75f205c8382ff2783a73a342cee5b1d7a107dd3e0fb4ace1fe401b51061bb00ab707791405296698de2a9c0d0499a02d8f841af73bc8ef55a250eb6729441e00b1a91856cdc2a4ffbd0f1fee39a59d6c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d745310a9573fa9945feb4790e6c74d27ed1a7c5c5dc0765cc6c040290471f556f61a353fc6ad2990dec326ec2f23101076bf523a0c849d5a9d7ce842f28da2c388968f73d956334e56000b8f643931f9d0d3e9118f6240c5e58a549ee871ef6b5d41ddbbec63057d2121799d8c40e9054991bd8809ec988863015a4055026c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17fe2c949e06d13f1d27135a8ed458110766011db02a138e9558d231d6d716fed1ba39c23004864adb421a2c74c5011c63ea489f1d8794e69331b49474a0f39b8507104091ad444efb225282a3041dff9be592f8f73abbb16401a43b501fe64466a5d6b13ef20b3339e0409782fb8be300b3dfdec3089b00b917aba157c3969f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2576f41155c8958b3a2c99621e144d9bc7a5f0d36befc7f0e75ea1aef1a159b16c0efd89c5ee5d58643f858b732b5c22a72a71335df257f6b5747b7ce86275ba10dedb537a481d1d8826433da9e90b066f07f0e3266d3e5b11adcb2fca6b78ee8f943273218906a85d9118e790347007869597966e6a70782db90045b706f83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c330ee3b8270427d5cf51bbc91abdb0c822e5aa501caf1d03bd632e77a19cf9ecec24e9947a18b1f6e34934343bf61b4e3e97ef0dfd2babcbe3b3b0709b1b3242411cde86b4a17a2f9542883e65c4e0b8fad1b949fe61a8661194e2a45f0876a6562407bfbc866a7268c6759817e7a24251beccf2cd4cd5cd02ac71ca54f9b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cea7762549bccd44a5b9e7550c6f7bced0e8160d88534e1eb2a8a97138167a41353a37f9209d05bab92d20b67b53a4b23194d0ec5dbe07d30d5fd6a36c320d31e7bc627346f83ae8a08ab003b65d1ba5e5e8736a44ac1a098072654211a46c5de4cc478d1139b46472efbf1166131dca1302639dd6296e9bfd3efec6fb44cd9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d25e23ec00f195912d196c2b719f6f0a0e71b99691b3772f30ec54d40bfd2d2c0b8c863e3f84d04bb5e3c111dad2648e0b32c36dc2bcc957592db060a9a34cdd44b5820e3318bf3959208e7deaf31706f83fbc84277440168c2f07ad14210bb549913692fec9178687692e32f3bce55a284f4e253d3e1a24b20fb8aed55b1b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h400992bce41c16d0ad371e252344c932b4a6e7c406825b5f4af88fd3138bfa9a448fbd01c12068013af157270426f7b91a9413e618b16824bbb9b563d188779c84ff4a150ba5c009b5fdc6dac084eaf27b74018d10e10d51a341ce885999e1adb558d1627964db8c9cc47193dc20fcfa7671f538a9506c55dea4a7d0e01d6da8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72044c528124999bc35d468faf28c127742d5424d55bd13c07218410e4327d010134a3765b9ee070563bceeeac3980a08e1d0d59f10b5cabcdb68c9eede4b8ad57d30fe1bd6d9de945ad291c1f47a51c02372fd96182bb2283bb88f53c75e12cba5e46d9b4eb454120e9fe979008582a04be175c2eb3cf7ca2ec8ae7af4703f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd79baf84c14fd2dba66ace91a708f6884f8d02728ce7d6f469942ac026cb093171304ddb338914c3a46bec4ea04b73b47d5f25bc9e519bfcd0d5e37b1ba708d30b712c20a9d9cff6fe777cb11556287562ad360870ca2b93602103a76c07265f7ee176b2a08457446c1497b4178bb6a3ce94084ffaf39d21a2a9ca1ffbc4c2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b8e7d838329de08740df0dbdc93c502ff326a2c049ad66a9691e8c079cae39df1bd67bd460b3c9614d74b566328aabff13241c5584c363ceb8ee07ccd10437d4f91be868b2de610b97c893da0f7a6d85bdc41dd3282e936dbe3d41d512f19eed953ab4f322f19d771e0e32786ad4c7566e06ac699a09047f56d7358b52db554;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa8895f82908b3c0539d1a57a5274be04789db143a10a8a36ba70f9b83589c9222949eee5ac78da03c1adaedfe3d1ccf6402061ad295b2f686e280f3fd29b81d1123585b220f1263b1aca470333385064dfe0d8311a1909efaaa91c03d74091ff2bca3eab5c8ee8c6252b790e319ff865c9429921d42459c07157ad7773e1cc4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha72b64a9137f9f74bb48063033b10331f1da2e4d5c28ab76642f0f5f47e2cb0779e94acf69c525ef6cd972a2846e8ffb21ceae9fd78f9864d46f613053b058168fd9ce0c27fd80ca21e57feb87ee3a6ddddd01ef9daba95db779f4277f5087c39c44a89eb9939c270830cbb26f4dfb33752282aa0066a65b6edf5f937456dedb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d00c595b05241cf4cfb523b28d36683ed7e730f529681827f26b605943fdfa98a376006ebf8583fd0e4d0661ba92548a3d4e859107ff1676e177f6bf2ac0f27e1b2ac0c576255720d96bc14fd6e91226c5e52231815f528ab844c31f9e45850e99ab2313c2d5089d4978e06b2748af8280274eb85c21653df853048cac335a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5c1f3ba3885577153bacc21ba711d5b1fe366e62a6ebd87484a7dae07c9c9af417493a5b96d3553707f30db5eb99bc0d722c03ae6d543b6740fc82646923b1b1b8d215a64124d0849488d2015d8b3c5b6f21779d73aa4bed5bd4ffbac74e94dfe7a56b7db176a31bd1787dab290c9f1d2111e9fed65eece56879e49ed77ff90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c44482970b953c7c2a8e98a7905377662399762c035f7583c026ba9761e13327cce5160d0a0fc401458f3d9df4b9708225abd45ed34f15c09b82d8efa0c0c8418d2c26d1755a03c157f2f9cc3e48f6e63de6513bd0b0353cd5350b4535ebbc14143c3aa1799068d5b286ea0d6ab4aae4e5f02fb65eaf9edf9c9c6a37d4faa5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3ede0db44a2a46489f73d8502600a971bd87f59707fe19a10104b1c2a36923880c0d92563060f4f3e742d473e2addc12cf3170bba07b7e3f9fa988b16cd9f1e5b93ade32e2afe5d4afeae67d7e9ed246d573c6fd47e3e0b1d9c890e463a3d6d302294453510e06948fd3c8bc2b5fcbd4292087cede333364e9b301043411fff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc77cd980bcfbcf12fc5dd7dff0efbf64afd4f2de96caac1bc815eb26912da5ef1c9c1a945cc977f6b3235743fa207def75d393440962ca938850a395e6ae435aeb65ddfe9de5f61862d3988e949971f56c937964fb889c5a99e06bea1213670bd1accd77b1149955d463d7e01036a679607c19cb6fc838a9ba95e1dc6ff32d7d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a27f43fad4331dfa55e718e8a93cb8f54c6ee7248ace8927ae09d097cbe9ee04221f1a761b768bc1ef64cceb7d3e1271a0d4fd095625bfd39e2022ae8a19b9b7b5971527ea2889df95703748b9a985c4a1f7bf22327445aef7b383d2bed08622dea19e694e8ffaa438744547470d010fa01c5cdc51d8c264f95ab17b1229354;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34b6f56dcf410e1b5b61c95c802e63ce15b7e30e0849732bce9f910d57699f62d0b69864bbaca60b8a512e8d5ece09e193054f2ddb77535ede4f7baeb4fe1d06015357491be8d4cd9a8d25f69f7d398a1b6c5c6173f0bd29efc10579206dabc76ff936d8431b80979c9ead7ec4fffd7e208e44adb93b2f0e4ced9cfbde11318c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h507c526c6593d8c207057318e35a6e85014e6deab72aff66804db128b207ecffe486e3f520443d3980cee0268454d6d79e93f5ca597b9ab03cf569442d7407c1d035b589174b4d1b16896a26b0cf4c332b7c6140d925f8ed4f7386dfb47410b29668bcc52a6dff8541a686eebc0ac193387a249316565e97fef83f47311d5336;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e7057b010a6f8d89238a4b1adee35255d3d4a9cc4a2585547b4770593c1901488987f3812ffb2ad75d3b261430ed6152f22c9e8c8da8e21d8196cb5b01b4246bc3c4f90de33a78e26a11445eb9d6da7d51dec7d5871c11c593d3404e2fd498cd57a26e17894a63f8ac76b5a4aa3a5e85865ba83df103585db30223871824e85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b9eddb73fc9295b563717a106c00a5e130328e4a29f292d64996dfa580decd2793420d521a7d6ca548861b187eee461751b1fa358eee25afb8c00cf86d0fe463b5dfb7f43d657d6a8ce466b5c8844391804dbd550557352c7255251fa3e94bf0abbbf239be2a59f8ce1c7cd1d086276fa9c2d63a2b2a4829014b8de8f435c31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb904505489abe92bf70d6d914d251dee96afd0eaa6d593811aef2e2ba64a803f56228d970ef90388070462d494f05af92980525cff1d9598371e9e961b9574dd8523b939166592cf6e59a85aa912242b45b262fc845946be5813902bec75717674ab1cd27ac3b1d296d1466e656bc7147a198780782b17bf0075c55706847577;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d951998dcf4d5abfc6de5e2ab93855dec4d6393ca65e389c9a91abb2c28083e038e7d7655afb7d163a9f195229db864843641ef3b43754675c8c04c1aaeca831ce8162a8f6dd744ab2826e2b12a8fdccbde8df47faba4eebf63210c93aaf17a09c7d7691f48c46abdc495700164d10b7c5285365bb83d8e351c406a5b597335;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h870afad809891e9e6c188f3021a343c466b24ebb1442350c598e19272ce03d97552d9a76ce5822ccbf2c33ddea2cd103f00e2196e2ecf4de7ab1def10296920282ff726ec529954ec500f344b0335ae4c2ae1353a7fa0deb0af907cd999247db400b546836c351b2ba2ba8a85dfbc8035f629d23cf06e7fa08557e8c5a83d824;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2f3505c4e3e469661bc2c342ac0cfc0c3616c3ca78494eec26a13ca55d084283e704b0743cb419c97264367e0c6b92ce471dce7ae9216b1ee58250fb704c17da62595d5883489f8b06612d47cf8c6251ad3cf6443155e05bb9e1abb5f2eae6489cc0e9bbf9f240aab3467e39cacaa04b12374b61ace4baf810b52f1e3f59bbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe44111685967fe73e2ffd93dba9946babe3ad6c9d360bfedc49b6608035ff160be144c0a7452c1d08a106653b1531e42a6f116ad46bebd0ca00acfad3349fa7ee9797b1119758bbe3ffbbd6d845ce65bdc4f0af82f490f975e430f29e1ceb32ad9940f19ac94d5586a1b0782381799e83702ad7cae6d8207a3dd5e29326f6b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2f79187069ab44afe0b22fe5b93bcb4ac30a5958e2aadd15f165232264919db537ef8c1b0847b9e716158b4290f6e10248803890576f9b5ff837e2bec0edc628618a353a735952ecb20c2cb14fc925ee8d958e0611b1afe43bc3381f071ba13cfe9b12cb72e76ff104068b4d5d13b92660a91bb7552a1d2f97cdd6a1ea80bd9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6da454df35aaa6adfddc6a685f3b4cc2478cdfde71e7921abae13f19aca72f71da32ae372c9b9b12ddca06ee916f1556fe9ccadd8eda0bcbae677e51f46e73826bee48dfc15d9dea0c76710ad844fc1e5631f02d43e252f656f0d9ddd5b24f7ae6f786c8d6bc91ddbb899dcaec31d188fdf8bbb371f3b834d31dfedf4f74401;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63cb68b555e651f0213d3d840b505ad6387534ce2633c2814f0fb8ef64940245fdbad0c2ecaf86e0ecae62271439ebc14f17c719f0affabe56b13c7034b83d41ff3822e7dffdaae4d6eeeb1df1d63e8266f07411faaec29cb3299bd5dccc6f85a7ed591ccd08bf5bee547624ba45b280dbeb86ff8e3ed8a189477790a08859c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc23a1a191becad368c47808faf43702aa0afe779c28d6bd3678aee15e792f4b5cd0916f2015bd7d6d6ad782acf693ef59ae0d757b19790f7ba4f5cd6a58039c2b1001b48834759259b444fa50f8d28e5d27d096ed49992e4cb6c14a4fd916361fc53612a1554751877558fc263929e10401c291ac620afb9fc1e96b205705dcd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heca6c5fe667e0d5e69b4ec6ce940ae7f865f4f264c2d10573b0743394f9ddd8d2418924caa5bba6a54f84925216c4188b64569d5996fdb8aabc4006bd45d90a557a136e8e61c4fef344abcefc89867d3af9136beb0d5818cb6f2ca7b77de47a0d1819abb2f32c0383408265a5ebc4cb2d1114e0607e0648e63bc72b0508ddc2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59cb211cc8997c1ad522695ddb1b653ae937dda1e3a813b2417342b84c87de0cdedef601c4f5aa945a2fcf2757e186bd6cf1c67bfbc6e2941eb473bf5c27ad868d980403311e5aebf6741faf1061bdfa67b70cc78ceb9a6bd6b484b9d8d349e353c4772acd2419f64f1b48d761e8e140217ccf1ecb2a0f1f9588cd9b144d8185;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h156394d4189711f571e886e4e804b53c8d32cac6bdf7e1503ad384c0272ed6768afc145570b0bb96aea2b4aa44e768962c758277cd037fd6f5623cbd4ea696cdca782e93f82804e02150d770d6f1b995bcfabbd74b39039286aa93ae71beabdae82dc704290e6257b0027e84801233819e37471934ab4c8b672ffed31881e286;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89fb8ec963d5b1cbe50971ee4e0149a852f02eedd90b6896bd60350e97974cc1340981c4ba82c93804fc3874d2128f42157688cb63360b3fee0070d04ad3e60f735f3c6ec6d0aa7f1a309c3e1f2482f7e108693361d36f4bcc1ac94c68e483914e70d1692db2fdaecdec53c909a4d5ce38b3c1d8f25f595fb40962337eb117ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc4f5b630e3a01dd184bf720f3f4a3f81d94255cdec63133285ec4497bb03e0055977da6ac2b7cb81a2aa4cddc6e9c9ac63b84e817cf9e94b0d4f39d7dced2217318e458bd2d8fbf4f6ec3fd2cf8f02d01176ac0d1c15f82141b090de6e6819da4c7799d642fff09c805bb79ecc1da46d30a6aa509f54dfb3566a2e978675971;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21db90e9dca2143a131e3a13ab48151bbce28ad64d729c1821a905cf2e83747ec0531c9eb494113ed021e91122c70e3cd6c35d3edef0833eef15a84027b265f1cbbe0ddfa3b1aef7dac6172702d0fe583b0b33a5ac9680beafd2942f2a15827463e14003dd750d84edb8d3871d1d9d4eaeca7e5477c1dffb6c5e8a113191782e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5c761a8d1bd4060fdad3b49ccb8dcb376b58e9d0dffde394a7c149283d5632879995a1a43dfc7f4879df2c89bc341a773d0471a4ebeb8cbf04c15ca860fd53fcef874a285901861d3b55ef6c8d5b736e306e0ee6612f638b309a034f8c1a458104ee338c94b5b09743ee1f67c2135fcc011a1aedb5a2fe7d5ac11d39da4b986;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11c600ed4c1f66a6ae8bd48f3632ce9cea8a1b4f8cb862d3948184392cc789cdda5b77b00b42e658abac317ffdfb791e64a5a2ca3f666796adf194ff66717d09116808a577a6cb208f4dd135284868e10eeb229cb43ae04df33bb728fe746745be85f5ad24272c334124f758eb55fb5156e85323b53bebc20ec0310047750dd8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9b2e12e279a5a0d7eb32d55d052e7935bb819b3e00ee2bf2e3f9c3f11591e19ef38fdc666be3743c96ebf906985c210717ed4ba8aaa5e6f724ea0af6f723bf29477f48059ab7de055d0f058267d20df0bce578f5e8aa3facbc8c60fffd6799dcec4a7476226f52f4c87286630004249f615d41034afac0d80e82d23b255eeab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57fbd05a2a7b9e77698bac9461f59e9de3660473a99675e4481c5c5cdef179f56c71b70816e82883ff1e5aaa1da3d6285449ea5bc4b5b0aa236daae629cee215e9cf6f390a90806bfc39847bf7eb17f828567e867b9f96d41f5710efae629d560509d4d83c750037cd85811c45a56a0661d12e6a3c254c186470b3b5d2a888b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94fb0ce3b8fcab6d2b1ca6e5303455bbb041ab947202788dd08149fa97991c3b6d6f969ada37fcb5a8d0692e3e54341b9d3b4cc1eb3fdf3ccb6d7419a4c476711baa2de7c067b4b40038a608de6a47b5622a0b4c45735605c718fb790f8d37e99af51edc7c5e74f5ab559d3d907c88e2b49a5cf89beed15330284b2272104ea6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h577469cbf66fc59902cd233757559d55e958503d2156ea9ace623a477d14e500ec63580a0a51c9705283ee1526850f85d1400d79aa82ab6b3da48caf4e5610b0093f51b5dff31afee2fd75512a76d14bfbfd17dea9c401b2e7d8048fc1f2e91fa00ec7460c5c208c70878c45fd395cd12fb219f500c429a8650360cbafa112f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d29df2510200f5951171f924ceeba325022855383842db345a38a50ea73b8a9da8352d12aeb3983818f7ae0c12075b94be6b3f8423e9fe52b0d502cb5829b7a9ea62709c46b94868df3592fc95ad2d45754745001b70a7db31a8834214a79dde9ea1734c7fea3974a426a9bcae6a7d5e2281f3377b3ca38e7ff4d6edaf8e7cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37f207ba3623a229f7c61f865042cd4444ebd400156986185953d8534e4ad08e2ae11021aa4d73133ec74063230acbe6abcf7059bad5a2da3ece6453291b5effa6417859b37461b3ed23f37fe1953867937e051723874ee0549eeca6434c5c222e45ac2807aabd8dbb7fc92fbc5761efaa56b9442bf101eb732a8aab8baa371f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c7871699357399cc0fcd9bf6e24e110160797c62c8f9af1fbd746deeae0033c633391dbeca832315897def2612187e2cc3b450f843151d27cdc9c4906526ac9d5986d3f3b9d6d6b0c8a10c3d97ec235051649d21b26b2dd517c74222f475e46fb4db0954b8995a6bb1a41ab3996afcc28c7ea6e22b6680dff050fd794f62882;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86dc6c6d14b142eb8935b5a82a20684a559615034486816e457513e4f22dbe5f3158569c8e5958e61b0c6ea3169e59064e56941066c5bf4848ed449f30d3e76a92f72f8ac0a84b64fbcb14ad95e138861a47085f430b86bed18ce6ac64f13274214ebe785914e85eacbc12ea87a11864f9ff497ab4d62b79a75a7760d266e4c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ed04a7a47c3f345de43962fc29d9f5e98e8b005f8fc74043e712db715ed3f1a29d836eafc118fa760a4bf0f53b207cdad9e6eca028f3fe5ba75b20356945e02b5972081d11e7b1caf6e899d25bee876dc7acd93e5719ec5c10746b0921b2313e73b256cb017f1c0122f395e4032e9a49eec093e8248538a6bc039fd8c25c73a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f1e6ef015b2cc88d58303d9f1045a6686ef338cd7f77690f0b28bdaa53b12cf74f54a486038ad8826420678209c3d078e952ca1d7dde0168550d34bda57139eb2c34d2848543562f8ed3074fbb8418433a83e5b12e2fa5824c7bf53bf6f8104a8f8445a2160ce5ac8cb728f01e598fc59d93c3d1f1b430f0f050a4077d60c91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he962d5b776678756838c55f87411150f174a883edbdab2a0365b694027a9832e54fe7b59cbad395338286e8ae52f2814666c676fa0fae3a0952454b2bffb9c37dac0b6b370c1ccde0e5d2408467859175804070df6bf430692cc568b7289e7d7b309e5e48402434b1d14dfd4c0b094267aff398aa50730adc68842161c1d84bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he11770f4931da05c9d5af82ca997d49ade4bcc89dfbab0846e15a7ad05d880965a91810b39fbf230039595556073027a1324ec82e43f07c8a97270aa0bb8f1a535898358eabe36b5985094a72f422ccc8a3df0d0e58f63d60a799d1c2ea2d683d3c04396096ce665a61c641edb254d228c37563c5f94c4c349dde5bfeec20b4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h419629850f72dfc93b5b3260dfab9bafb61e49ba16459823dd0371e9cbfbc185519c7a17573c2b50cb1345ffba4ce67a39e9b3160050a43989b1dc531546acae16fd21e677e957679ea7aa0cabeff4817860b1776cc89b7b9176a3386647c499eb44c01d898eb413953445216661880aac5eb9352972a7020774e87b172965b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2ccdd1b68cf4d7330e2adc7074d81653e8cc852d0efb6261bf884429c75e49851ed0bdf5267d9c934e19fbb90d6e61604a2ed224a337e001cfb08aa0f5d416a0bd5e741f33a6aa3dd74758c9b494a4d8f5641cd34799d0d6e9605aa5dd4e7adc4f5834481705b895aa0d53ee41a5b25f3b6e5368d74086a16ade03f4c18c59;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h764002dac8aaddc37011e998687418f79b2daf9da1542b9329e2b42c9ed0a715de8248f3fd6e86589cd0960d9fbb344a7c2b32a9097d4013b1350de107049c910d70d8768d8a2c5b431ed1bcb80f2d87b2b10a1fe034a0d9910d24d6b9a8e3d975303ef049efb0b7d21b2c405e2a38a2e8d48e4a3722d86954bcc7ec5739ab0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83a4c6cd046750e8d7b252a9070907a861482cfd267e9ae332239b70c6213e81438871871245344dff93e0e4169f09a06212fefd0b07ab849bb366d4aaefa40de3d757251967464b1cf04b28efca201102fff885e80fc84ac75e796be1a730412e55246b41ef39e51c3e6bb29d89f90a641243dd35abeacaa3549c8542c5dcaa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h945041a1a28bced053e345812786d030272555dbc911fc06376cfe5aa801ed552155881a11f9c77c3dc8a0d079d76e528fc73d526660fc5f1c8f94b3814f12a7efb6833adcb923573820cc475e8942f56706ba161c577438bb2655a11ec8a02fa5329bf79f532b68363b7bc5153ae25d1271392f4d42909d4827d06822773dc2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11076e70bfa911de4c30db161d18ed1461846421e9ca6e26a4cb6ac5df6021c72c15525329b2c539cd48d711ea7e605b3552074d679fa3de9700e613cdbd577fd2aa213b029893f68a90b5c389d5f87f57f5398bfeddc7b0eb7ad4c9ea9badd8916c77347d837355b3b8849eedfa963782eca7124478c37a1e07bb693a72c95d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7175a401983c56a2bcc30ca1e31bcc861258734b36fdcfc4b7d7c9698a3bcd64ee1ad18e8a1169de5d7108b8fb407ec655a06ab9766b59dc87d15244edbe70dd23469dbffb01a4e273d87b0175340a540cd999a4a72e0974316cd029d504018ee5315b3b06cc3dff1d6ceadd87d97983820c7fe00107d52508522fb22d28242;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd386911ed2abdd925ac3f453905d2cb18b0074d1adf0d967017462ddf520f03849873fec642ec23b1df94a18cb70bab4cbfd9b560fb454e4dfd42c7120fd490b21fd3617a71c0c727ef862dd92f74ba86bb5150b9cfd467d9ea4857c4916a3bd37493e79c6503b792c191d6ba3d827ea605f159927b81dea1b546644dcdbd51c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d50e4c2e3edfb27051b7e6cbbf80e47447fc738af4eb394e5732a6ef118271842a337cf9bce5b45500e06f54dc130efd7548ac2e56e889c9313fba86a231df721cbc75780475b42c195eab7f16efdedc59f96ab1c1a60b592a4c30eac244f49a4643f279a013801571b04fb64b76011a3e6b2cf06b50ae211a2e869bb67012a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h460f5bfd7e2b6dab74a03dbabe773c23330dc13a6ca6f088dfb6a595a89ccf801d4b3a21d2841090c61c484beb334eb8cf83f430745a4e9778c7171d5e65db46f796ed3abdaa9399c5071086288fa55b72d6c0c3a82368aa351aa4f65d5ec56e446f79a3ca76334c71a9eddb5bc0bea6c2324c8051c2e9a3335c187df3f3131f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he261f7fa9f267b47a5334585aa2ad327398a657351bc1c9330953417150fe0ccd42ad4b0eaa65ee035b6d6e280260687b7528e6b2febe2ddc54ae558399fd257801436429d97e785ff1642a695b82bbc620c35ee068ed89826582d27868279313deb6f2a6bc096fcb0d82a05c7096fcf32854927d43d4583107d732c9a620a12;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87b8177768b29791df978ca545d483ce9d24ffe78f690c6f7898cff8bdde1027305c16026bc5f3dfc5c350ad9bdcd37795868afbb8281a9d95b01b9be282247b1305e98d53d718162e15d5b32ed696ad07c0214ced12c935820bdd31404cfcc1ca5934d6141a11174055c8c8eead8c06446795c87604bdbae4be9887d1af0b0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f3459d17373124ee4acfa40264e08815de1d3838dab9e4bae92451baf61f1dcf7a35e8e0f5f8453cf809f5fea6604a6b75b653e6ebb5874d97729dc74b51c816d84742e6930fe73e934172c36f6427eb3fc32886c978f097b7c19f59238c20794ec3b4943d5394a8249cb3da851787c96aa97c90eddbc0f9e1c37b2e74037e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6eb98b14f4fc1f68cd11b935f917bd7da303b8876576bf2e4ea935e49468e542a2ec07c8e8674286f1c34e6822f0706a0aa5a87ad27cb9de00eaef6987dd32e20a3aaa691fd38bbc9976dec8e8a429f8a2de1be5bdc4844d5ae2a2ef44992a7f2330ba38ae838bf1fffb9e45879f862604d9c8f109a66e034026abd9ba01fa50;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3bb553aa19a85f7b441fd1f72c2b847e3e876ffc8aaf8ae330fa9b443f115f1fa2e337cb6377b3adfe602b80a925d2fb1238ea7b746464614a38102a38405fbb25506a4cbd091affc201a9206c836efefcf8c6e60e4f043eba950ae1ce1c84c32bf9e7cf1a6e6e59ac7ae9e69ca326aa687e2ad3c93e74f4bfc2ba9e05298ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58a7e979cf7b38186ab21f93c078911f6f3ac704eb0358c49dea48c680165f5f2077af738c042e5c24a1343f696466aab887c5d3fbd6a39388eaa9ffaef64fee16872daa85d6e38892fc62c9a79891474a86630f4e087c5455f34ee40540966a878e05748fb0014b5495586b18b229390304531ce193526234178b74624b6d3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78a266689371dd3b1fb0d9af0c8bb8243d002dbbae649c69e6fb88e87964ac33ab939b8646825ba3586d1cfc180ac1d98aa0df93a641180efe1abc33ce347c56796819589bd98f6fd26c59d599112331a7d391a750ef75660cb93030b5f6a9116325c2da5f01faddcecf2db99c1bc04e0e2a6ea7d144e9ae53a5fd38d702dc21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fbf7698d51290406869e866c8d4c69163997f429c76bcfedb04f4d1e71dbca6a96baf7369a00ece8306a19f1e4d512b197027bf3071f8170deb4a354744af0e008d28c316f10f0d938edf43a20fd1c077e3a3bd5dacc37abcc1c5fa1f923b3304a53361ae3fd67e5b576ec813c8a69f70b98c64dfd6f67d163d381e8d541ab6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc515309fdcbd5dbe816183dfbad3db0891d6b9aec06ba756c2ab34c0de75fe83a5e9e9964fc065490626118b7908cfa82ef55314f8eb2a4c48b1193eb6196539acff0e53548ef887e137c17d912a5dd25bc96a07772a2b78e41b30ca774c7d928352ff4b121e680a9d2f0096e9ca8b91b51029658942066d973deca56ae2c353;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde7350f42c2f519ae30bc0ce252308d17d06bfdf8e428c07d6cb12ccb0e274c1464c67961bf56a0f76b1213ef9ef1480275648aad8b7fffa620b880b1a33dfba295110024436debc071de11b70933e5c025ec1ba96076ea671d5cbeb91dbb54df290ae47064ecc7a8abbcfee071650a34289654a9377dec96e26bd4ad1b1224e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h529208a81e8f68b51d076c9383514e8f37bf926a1d8048e2083fb4868bddd955081048427eeae404573b22c0ed5914ff81130df8d459b9589664a8b2dd6213bac65907d119311580f3a46a31ca29194c8dce0ca0b778fe0c3bdf655a71cf08216977d77c6a7d84cb42b5e0d06c11d1e8696bacf2c3888c855c79d19a627cfdd0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf70056903fef34fd16d8e9a9ebacce7a3eed1a0d0873bfe285031e83f14d630ab507604fc83a6d27c784d58b047b88676e7f9dcd984387021e4040913b0e6e22bd7a90c49643a8c7b1f2625f3a51b2e08e7e59322e5535fcc1069c2c10675f99904feffb7c8922e7eda230ae1bf5c7cd602b8f0caf09473e9a078c13e69c9f44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b3bce4273332b14f864eec853630e9c9f5f993cd0cd516569ddca9dbfca3a913095c036338aa2d06e305a363e2b7593dea73e51148ca4b7c1b9d9225b7d20bb620e897cb86a7276d573818240f76fd35d3bdd882f5aeb4b2a76b5dc42805ad18fd430f64583278f078cc37ecf24aec9a7a48717b7dd067c571f1dc31e453834;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3111ff8a63965a7bfd6cf05f791aad8139b90657807faff2202eafc53c0ad8ac9a633e8ce847787245908f809295d382fe938e1ec916809388dcf247a9e13e695d537c87285dc8877407fcab67b9dcf8570108800a4f19d89ad4af366ec32d4cd7efdc33a91a05f47f7d7d19285d989e716b5a4fef2356eb44650abc8c47fdac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2b7e76573d60ead3e0c5be61e9a14e730b2b98411e48d2576caf588ec949796ba3147eeea88facc6d082ded0d3804417674505ce025f43e29579d365f3dd4aa207c1a2a7750b83af8a46d2fbafc7b68cc602db0089ca6a2d436272a5fc208aff628483b28dd963817d032238cff6405f591eff1a09bab8c09b08ecc17e5b109;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a43c6e7c7921008b5d619f1c0e6da27926d60a776977516e11fce1ca73f26c8981db11252aa0a5e20ce6a0c74d70cfa65d9c440180d6e657af2762b3160c5d3d8af43d17dff59cc85a2fb35b02c2abbbba717f381a75ad06d8427d43aa181f0dee09b0aada0dcc9992d816d4060548041616ffc64dbbca3a96b95e81c28e33e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h16485bf8a7cf0658053bfc5635b637f7c7a4e8f1dc182435d7d21c5dcb4ca50bfab8acefb78a274dcdc0613d4655a593e92a48691a4e112e21da2189c4a39793b32431d1fd1f7d7a5abd29c32f8ed14d48471b146b299082c157fd8109892024850773e78c97db2617fad55446dab22b36c6af81eae13d76ed22b0813b6b107a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcde612b353663097ac339f479c05ce901d5b28daab358f1e0fc319bac32afb3f13561a88dde22b4a43495a1d62a7561e42bbc26980ec0f55aae934f017892edc03b0e32657b48c4d30e27884d0820c2b69f879372c9260009f0b357bc0b455df74afd643853c102a88657ae23bffbf199392348b473766cc41d1f949cfed607;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0fb9a464abd6934c90e7458653aba6781a73cdab5fe2ca5359a687427f949ed57c8afc1f31da0aa887caf2d48b5d127db34f57b34be3bdbc66e121b123284dfe233e835377d1b2dfffea8b2bdd0a6be7008a247b90e02b59be1602e9b11ff721abd232c0bf93d7a248b0ba9bb7bef63f27ac00b21c3e38e496b698ad0221b44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5e632ad11f7dcce83c27c81253e7a4287de495ada476c4e27f245461d336e64cacf7911e717d244728fce721f83745323281dbb1a16d2c02e8d84ccfceab81debfb7e6a01624015e7fb70c3111b19d1540e801c1ed881978b6d45749e199f45a212644786fa8f1252bbbb0c7b81aeb3fe0f2fb5315ddd0d15de098be3a1a25;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb80d1c339aeb9c6bcd8c6bf35e907d0077f89a9a067f242ce4081dc15659a9e104d67f6ac505e9af7a443840376ec53783148dcfb6f1564b1230198fbaeed34dd6db4be1b3505f6af2eed166a1114c79a724e2e75dd8a744b4ef1a2724947fa047c9b5cbeac72f23e93e3b31a3dfc3421ef4a72b1d0fe62aa572056ebdc1bd33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4cabf742e446d98c086057235be6dc3c9f905f12523562a4cb96569442dc584da4edb6f4304815a62229205811cd46f67922e2ea6c6c6702a939fbdac5305f3bb0eb406d69633478ae5632eeb73d2e64f595e35390227fbe0f83e4c911d5508f1bcf5e275103d651d5aeeadf9bdc943a4bb4173f745f99f78e73fd6465fd0c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1e9aa6745945363d5bb876f55d496bc07d093155dd31a7fa3064a29bfffa77c232d8701f23fe0471ee3fc1e44cc7e861db5469cee8f6b9c112dca19b2a75deda3dfb1abd6b4709bd812ca2ad59a54ab49af802c5076d33825ea531ca56ae0eca479f2db60ddf6131b8d0008121ea3ff61817be4b8afda239dac6d727497f9b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h132d09fd6c2f23f4d35af946077bc4266c191697d0ad9f42f09c506d6b0cb473732852a40aeb73b1626c09aa04a0f1dfd91b2841682d2f128935d1cbe9e81451faad058e5c42d811b1137202ca8dc133d675c425917feb0f53632774629a6bf6ab277e335863bddebba7e32c6e55185b47bb405ecdf57ec30f9e2cc33cb2496;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b36c70e2a88ba5665a8563c2dd105fd999d452a8f119b831039dadbf905ffdf5f57872a0dc8cf2ac5b18a5f1d13c9f418607e639d3baa2da39449430c0c367e7b799117ae689d1457b71d032fbd341bc6095a51795e7b12bdceaa28992fecd3bbe9f04f520c775eaf2e778c266266345c3ee2cf151a8e7729696f4cbcbe33ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30de928b407d3e00175b5fab616dcd312625466f2f73f56544e998793a50fdd2326ce42d90f944e53bfa76b2ceb35d6cf689c9eb86ddcf054049f76baad1496f4e26f163c8451ad4f3a3c331da4563d011fb8e1605203eaec66c95dba42fb2d7872dbec86584ba11f390a0d16883957338c07a659a15fb317e7a8366a10a8976;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha898ab6f6adf11821a9771efb9b1ef014444f67768cf02a98b81f1fce75aa4440ab277b0cdcd45d56a4a88c2dd0af64538c12aff3517738bbbc7f384a69e0062ed53722c819764e31a9918a1c103413fd9a97e1d375140332bdb28edf8a4adc7d74056401836ee95d5857cf880a417bf974f1d06ed2fd136b38f28eab69a8c5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46526928dcf8658b9c8ba10c09d8f88b2ca41e1f57f40e36db02517661ca6daaaf8fb1801b67b2c56ded49cbd2025c138209129574284d624e77ade7bec105bc311a7caa3bc64fbde3244701afa6347c8e0ce8d4d0e049911997acfe8c20d3aec05572ca739da0cff919e5dc6afe2219bfa25f9cbad4d8d2c293caef6e620c36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0770d92bd1d5922b250ed046a1ae917420f4bab3e4dc7c25284b7e09206ccbcdb6dc9edf7fe9d7d6f6fd175c87c988d9971b52651d83868952702a8f0389c7fea3a94102e3d203938344786a829d32810d771213e36d566eb3a2a26059b2a15e2962b5fbed812cd8379c153d0adafd5d803726795bdbb79a75735cae54c1119;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ee31dd85d137643d98470afdad40304387c8dfd75970236a1b9f879fe67822253ce5999a20564e7b83c39e9bfd0ba3264e17a1abf780b10a4454e8b9c86eff5c467f63b22141795e2ed5b70d1d00716955ee290a252d21a6bc7e4e8885c28b306e25c7177b4e6ba99562ee19e5bcdc5439bf3ca1b63465dca4e9e12244cf282;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a772b157ca58fbfad9b7d9fbabe1e477e60b4b87c171890bb94ffdfafaf99925c68ce67b58529cf532b30e74aea34b790da51ca0cc8432dc96a855547bd4b08d298b4352b450acacbfc6e668d8a0ea7c245b51e43ebb0f1c44fdea5ed901cbea4523317c223ae26811908b9c2772d5505f04efa296e411347cc904b06d1eb71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had28a6e1340de9a6a852124727bc4cf379113df9a088d452a448623bedd069394bc7877590e76b115b7d229b0e9d982d477f11c62126f5059c6e808c5b01e8958b240b0ac568a216251b06438900e7f775b931e34c8991550adf5ec48183a31f788f0ec07568167c864dea41bed3ec0f0af86a8f2cb2ecd7666f531930d74503;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebe4e4a78c58edeea8acce66f1cbac3eac2323804e864547aaaac733966712e57778c28f9ae9dde7bb3851b28b330e70f1a97439036b7e3c63429364d425e501fa9f516508c57eb9bf582ed75efa5e6d047a362ef43a79a37259f7c3e555a1d1c3666867b5a4fd50f61c19dcde7ec0fe4db1bc34828de3cad6d74f8d7f0e8b81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84c75febe2b29a174bdd2a125dc52708aa006e9e2dde9836c90fa884c1ea1b23c249944756cefeb182df97fde37da30083f4f9328df347df59a9bd9f4df63a990089294981fbcb82471e29c000a7a61d3d96470b8714bcb16c5db8d7639cc16e9b3c9cb7d74a6310dd4cb01054dcabbca098d517e8f805ad20a23d50d566299;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c7aa9002084e0813e9a56a7cfb979397fd745e1c801ab8f1fa0dc7fb3fb9b98be048ba7d5e728b1c7e13d17875214628a519fd6d4691b34502b1db114d426246cec9ab3e742a930b0a42f5fc8f90b728521b2926b136e6403a507a20d48a9409773e6955d69f70dd8cfa8ebfcb47493c5d07c601f33aa540f51f720afd92bae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96a7a546c0e12bdabd74ca988dbaa59f775505f54aeccbd8b03e81d444a21a1f8a888f546b037f3fdc9b31ed1a5261e48f7155f7e719a2d8ecf7a52717f6a189b9f4cbd46b0925181869dc0e79126b80ecb9a96bdb2ded96628919086cbaf2fbcaf2956bbb70e404b619fb1c86ede1e35c76fb2c12f1402b37af1757f3faadd8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29804ad39fe3faf5052e889319e50713c0e1cac6772ae394e9953c6bbb04a0fff4b1a78fb9ba5bab8f171aae57e6d07d15ac86f66584e4f4d892c88f9bf5f3f480e4e873ba31f5699f7b9b9ca74a3fe84bc2ab2ba041127a9878138d734a22cc22ebfee4ec78c8de1c0500e97f7c632ad87873a2e6cc4d1c30b320893a769e6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ec89419372b9fdfefb42adbc9c292e6c88b5b6b4baebb959519843c9592d254555ac3adc3a9951009338efd13a9cefc8a9e7164797694e422565acf6dc0b0ac215a5f28a4d45943e0423c58c8aed24761dbeb08acccd2999c8858c618d89505942dcf0f83d1022afcd0430888dd025da082dfdfe642e41108e34539c1c9747a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c6d1fb8c18b96bbefea1cf3732be58733bb801e7157af05113b3bb88a31b40bb631f221593b2e923c094fc8aae04204f862cc7e3fb6706c5f4aa8c96877024f62b4bd2dd72448cf1441029c3812b26b2191ddf1f409d535dda11d23fe30258331de1b5b9d8dbbd908fe8dc4efe482ad4bfb3ff20bb0c9a2ccf2979423573001;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8338cfa538fa372ffd195d49d1fefab865ae13b65c1305dc61790278c69c9dd450f91ff4ed9d12b8fdaea62c966fe17e2077482b4833ef8dd9c8f13d5413e19d7cf4f086e96c6873055125c25fa2024e54b589b3ae0e5002dc4ac318d155dd5510b697cd5f629e8fad991b89f1ab09d3e3dfe210c1ca09ca4f30fd14a2c829a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e6fbea7816287004d3bc23104a66af91b636cd1245a10e5b53ebed91f4a2d3b4ac80fbd0c91c78ee4536991f4bac4a4e33969193a661916a03ba1b95b3ac6b83f9fdb27b5653343a4f6e33b17b7b2facd5f66e0eca70f26e21c7415511ab2c9fa40bd21fb513ce02a370902798630e993bb8641d51ad64c86053614b9a7854d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7284cab79ce226f0f24b3057ef8c958a63792ab06627d96dab78aba164e62f1536fe298a524aa25cfe3d4f9e2369eb819f7f8ec31097ae6a10df01139b0426a84c42a5957ec0f6a32cd4cb74b4ae522abf2907da52f87cabe31e82f9ed2cfdce485fccda951664fc1adcf80855276968c36b66afcfdff8bd7d519092ec140c17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5d598bfe34629d0edf946fe411acfd3ef909da1af07aa478e753b952c4006933bb57eb866f1ec8257d3723f3fab1786b406f5acd05e5eef571f4873274da6bf3e0544f994e132eaf5a9e202e36eaf36b2f25b555645b8cc3ca8356e865d385bc2ca93edd639f5559d502c52ffc7c88dc50d5fa0d9a62148c2c19c4e2e984db4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61d14060282cb0866e47270278613e57722e72ebd67d69d5365b2149a76d25859ece91245bbfb86d7d8f1468a2a31a270cbab5e3277822e0e27b367046ae4564d012c19f63d1f594f95674a0a79533f974f05894946ff6ee15e829be776285d4133f1337fe09223fd5223e6ac2b9ff175def047b34a6430e2bc84d5dedac6db7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf96159d39897e91e6858b2415f452defce019f39fa5fb16a4eab8940305fae11e5daaf5cb61a2ad8ac2c4db1e3c71d2ad8f3dca8c386db88ed21fcae3a4f5696beed164ebc56d6e07a7ee628e326d0a4d7ef441f5b17b4dbc56091d9a62d26a33b07a400ad5468564182fffde302c64e009c0a7c237fd8739f192add9db058bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5940def1f527293eaf8df87f565f86bc381d0712695aecbe283950bf4957452df67907657530fb80565e0f904a9965fb1759fac17a0119cf6f89d5e9b97c25a530df6737b7ca6d5771cb6966f50793b2c0e7e42006e4bd311fbdc271fac3c1f7e3839805fb9de232118ed659481e3f96723ab88952286118148f0df8e7611b4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b921073ab07c2851d33716e2b2cc0d1330d1943aad24d91142fb1df82070652f7e89542788a9ee83393f86a31510958b1727e46ad986ee60b624ad75f056c9ec62fbd22de81ea7ae088ce5a47cd0eecfb0fc10021b873c177d50eb2822aba4375d8182e2a16a5b5c705784b83e96d1e4657b3305a1597f06ba793babb99752b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94f9fec14f68d164f0b7b454a285a55cb2c16c121afce4d2453be9de8c8f68de4ab4dc1ede7f1f069f72fc62699fc4ec178266ae3bb16d3f89aa29e8c8fb9206c5567a0fe41c3fa5ad9a1c6b0240c05fbe15f13b6cccf80a5f6890ec8c47c7060b990a93ad94dba1969733bf52e63f40fa2efe82c4d98fbd7a83f8f3d54925a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23d0f702e1290d1e5a14ca5b1c62a1c11ae389b8f9db986df59a3e736d926de795fc393a92a434f67142cd0bb6db33d7f224ccffb6604011aebd45786fc756f7a867654dda83c277da38343dd9c52b721ed4b4808ed7330974ec3794672debc4fd89671ec0fab09298645b3600eca13ab6a9f49c38f31fea9751080fda7ab00b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a6ab4e8f6ca51df9b848047852bd33b00f29e340def9ae5ff335b03d3b078eac1c799cf62ab805d7d90682dd1b64eb29cbb3e2660731215e4428f3bca107cccddc33300a580f28ae7239526da4df639d2b9895ff41acb1551a7c969aee6d6c0c25d224edc8ec4bf43bb6b6f7c9921772bf005643e69dd8a490d41c9878e3686;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c6cb634a6c666ecb3cb1a15eb75213b4040ac65ab955965d12e77d501e14c2503b38c73e2cbf4dc0c94f556344eb7bb1dbf1bd93cde2a17dfc9141b42a4c95d10cfc2ab0e13bdc2f443a461d0b45d2a2cb77b1d6ec21dc895b2795e2eb57fd6cb063c82bc2852e74bb1573499d37cd4db290d0df54753cf0959f15f8c4b5eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6086485ba64fde562f2579a57dc19fc8d9dcdf93dcffaee9583b887d26aef23758f4d827561ad3872ae4516347f3699491d2c33c882787c3043737e6df61927fc1734150aaa3ab3e7ddd65f5eae1465039f607a8d4b85aa7ae47cba513a3fdfd5d7fc799dba904416326bde090d92d0033bd8954f00f4e6431b54f9b61ab8036;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1671e7b5340324b2d045d91f179df8641d8c614bd1b219950d0eb15dcfc641bb8e351fa2ac2d05a508e04bd231066377e9537a6e7ad363378fb90fdfd685e22c6e767b30ab52f8ac1e44197474ff3af2b3efb3fd44312a18fc4a5dc0a97dcffb6665e2446ed4ca500ab8f2c4efbb5ed211dd3ac91c8f98d9f8839fe9aa79f39;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25f42327efb028b533acaedea1644fcdddfad3215eedd4d02e560e35716569f742e73d70512765d6500b11f353228e457cbaa37a396cdfdde707c44118a479d019e12864075b9648560ea3832ebcb0c8e50c062218d312fb6bf27bd01d177fa2eba1e0d12c7a87b1dca7ae4f15d678cf5c85b520b86d88d55a1aabf45f690087;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7336f12b510aeeea4b805b3fdf098e4e5de2c0a175cb59ec997d16a024c0f84a222510c7255110be7e07d59b82f1a7d05f4e960f63260da328567bfcf072d979d62110879dbe76b402115e34aeef824bdd06e475f7e7b0708a3c74247725605fc101152b92d4918c8de8deda45ebf65015c7fe7028f84b31b253e08c4bdd3de6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee2bdf08c9abaf9b18e39e25cedfe0c2291832a706b6845c347d1d5b80f09e1ae880cfb812613a6776af86d6b5e7caa1a02fb3db22c3cc2f996f60dc1a85b29009dea0be28780754e3a498bf9366457adf57804b6ca34c3c31869fd8fd057923addb395ee917ad57623be03c50e0adec3c0b348792ac621c343b15c18bcc7541;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d05cb05962cd3110d20f357753e644e549905f545533a685808d748e5961f0c5a697a2d422f5a00ad0b3f7ea42ab0a039746061b5ba6a0c4ec35d58d164a75b33477cbb91c5ec50531e0e4ab2cfa45055d3437ff2111429156c1d8e5ab39fbe758634f8dace87c1516a0343bfd289851377d5e446b0b93d572434d4fe6f4a37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d5436f97580e576552646e7e9ba38d514bddab1db43f607b94ccd735b227da5c3f0024ae1864ed69382559d86accba90a0cbc18bca31c23239fa0a262f1754f4a4f97a49213ce36f3a8a3f062ae5b3567180280ceaafdd30fe9aebcfcc8014b439ad68fe9d71963a27bb7651932700d48671c659aaa0be2e0e56f66d0b87cba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h640e11c811d4ec9773460c08c6ae0556a2f88d850cda44f830e73bbee279fbda3bc37915d909cfb50a1db16486ec6d571b2b9f44046c3b1641f015ac225412abf067be047cffabadb2be19fdd908601ec124d9f156fa0d8182e66f186a00b3f6399aee09f2d5e1219178cc2ef747ac06bc4e755e134a5a47d4cbe549adb239d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h710faabf65735ddc80afb07a8e6a9023fcb80e3c0f24b448e3092c438f527d94a2ed96e4788e381dcd485c63c90609afe4d19c17c1d4a50c5ae5ce478bc3020081a3b8c009bdd850d13b6714b9aa2c2d51038487f5cdb073625fe8014f0bed61bc876a327f3f2640d1d147a06bc92bbfe01cc2453931f6bafb3a0e3702d6ca18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23f16556e39737d9987f8c6b136acc9a1ef9c489139292906816c89f7ab61144aeaec465c84c73e518b2e260acc3c1e7b90733153c00dd69ec5235a191c3ca1c91ecd590db18ae0edc21ad5f3844f0f795eb20ef1d250e8874542b5e8c8a7a2bb39e825d47efdbafe7af3040a3dfdd84e73f02eaf061057be75ac8e27134d704;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41728b37496a53e150186c94dd34b492f1ea7a69cd8f19451277de658f1e92d6f2f33f7f702f1c230b32f7d2918952fdaacf477e2e3d72c4ce3878eb2885b83de83317430a84cb403247dee0c56b9291ef53c705d3f67f3c66256dacc68d5e880fa03be1eee02956573d30384c22949a6283591832f43a26c851892e40c6660f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7abe790356c3b45061300ef634b333deb227a6277437069feff224bb3e3f470074124ba432bb0a6014dc09fc11048c0fcf25fd52d9a2853c977be09262533f55f52a71b4aaabc6cdb12e210aba78e0f68f4668384ac1d526d9871a9ed957d00d182845477d53f629753251e5ef6dafbd1cae2d93039fb321fbef905713f2e1ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d1d7e5e0bf48b64e6c792838bb696f1706d003e4e9fc46ad06fa9ad05e2c48cd524b5e1dc6a0fbbd7769886a3bd1d5c9e61fc6b67f1dac82526f9585c76eaac6ddddd953e728ca18f4032c366490cc78b44e2c59827a94f8986601f98e9b9bf3d11305878713cf9c4f56bbf6b21d42e70b8433ef43424f32135f639cd6c1fcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba62763ceea44b4d8ecce0b5dd3fe5f1addf6cb61c5a82aef9151cb7d577a1dd2ed1542a49bc5c857f62fd67b072ddc818ed526e143e3435cfba50bc4c0cdd81acaa0c605e05bed9ab066e4934863f05720098976f479a00de9274bc69e9382db8caa062809961b8f4c512503ca20361cc641866e5fb225af88658466c82812b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25056191fffe696f86daf49c90809209e99728cd4562a110a21df26421d64da3894f487b119580573222b71acd60dc99c99feb04eba11ef687572b324225fee6046912aa6c52913960ab5c4168a09984625dd0c54e534ed734b44e892a7e5c0cc88ec4a63ad4f44f470d9d27d5750935667be701c1641311bdad86145055209d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha213fd832daf6c6580042831ccbee0774748bd693ca48735ebb47bcc62417a6caf5afe439de349adc331d1ef61c7dc27c1b1ac1b90dbaa092c03192685de0f12ba8fb3133dbbdb3a71557de778adefedb6c1ea03943af768d36b6014a75701bbf11c24fbf6cce70416104578f6d8db2487aeee7fa8d70f39de5998c432ea7487;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94458dec632ae9430baa82bf4fb5eb5ee655c47079ef5ac4caaabf86d8f4dae1d518dea90f59d03a81fa9541e28db0a684e78231728b94ec88a7652512dd5eed2bc067e20036dfec682df0d949e9b0bff5be7a5f15f499c073ef3e4ca35353250c7f98167aba5d3fad9e508db73e8d9f08f255d7f790635bf8f986fdd89b2a2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3300e837b66886f4a01a3c2d4fd85b00be535a0fe7aa0a169548aaf94489851000bffe5901d3d17f9aab2aaade78e983a09be7e4e23bd42f6d84311af501cc40d371b2a0788abd9636a2bdabade9200f10639f873c9c0a55c4140fa6983ccf541261cfa422e004a049099492f02742cb90d600a97a019078cd5bc98e93d18aca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91b98556717328072c7bb115fb1ed283ed22e5f9d98fd707000789bd918029849844989b486960a471df1180940843efc7140a48f23fb91a9c4176b0a95de8fbe416fd39f96e1aee01a7bb02f52c83b1e43d608e43eb8e63431ff0d5b500784ecd5d784f1ba6849941221375decc51673227bb6c0facc66b571d915583459f1a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99859832df1668399b9f065e6d0f3a89b86110ba8b89a50fe6dcef0fa095d267420bd37b756d7ede26206a5883dd95b2a73ca614f856e7788828abaedc1d947a13fce27cf17563ebc61cd1c8bfbc67f52e1722a957567bd6d95c46bf4d00950e7ee2da4b50d07bc262cabc265cb5dab250402d3569c49466bc99b9bf853cb15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65cecde72b3af6efe3b0f3e35eaacd317f2c38a92ed352cd16d9777742124bce68950b17f302913678173803fe87a3b3152638bfb362989a00f6a3a79dfb2f955abc83633ef78b59563c346c39c342c39fb25101048011325e208bba58e7cbc889a718ed82d13a423454715437db446245fd0fd9de2b28ac6f229b7fa17e8ef5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4aa05436e7b6dce632d1f95318e0f6fa08cbbbd4cf58a0e123d7414fee7448c96cf4bbd3609de2bc2bb193af9832accef94d248dab8105e65af68eb0aecc473a58ac00712d90ae79ae8e9b56fc8041016c6f06c78191a43a5003cd9413b2125a50c2eaa0c835490f145202f7a9ccde8aa9097ca37a97df423dd2e8707d02a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ea134e21d1d4cbe5edc44d1c0f9fa1ae232ba03f2afc0b91893114f0262b04d602c8c2040684ff2830f77c0e2ec34cc954568fea1a1afe4a8ca1637c2c8bb7723a253e2c6333815c5acd7d824129bbda60fd454a081bc3d17557f0c49ba6f99d6ccfc14f26d6b7afe029fa0f941a4be4c9102f358781f83b706fc4c4b4cc696;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc64297270477ed25ecae240ad78685ac8ea046cb65ce987252f986d43b3af2df2a0cd9251f0ef646f7077b7373a65e4ebaede1798c05e2c99fc75fe5648568dc91b7c7989ecd025587e232a30fcd24af85a27a8b994f9b89e59dc720f110ae537d5908d402c395ca74b6fdc5486432e3a47f122b1569c031361f8dd1fe9e8678;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13e29c8b3ed451664ce08bfc03afe58339142ca531398945f85a58db5613de3f820714491d1a38581e7723bd4cc1324480ad7351369e5ee9b0b80cf746f207b4bf021d281885e8d817471141465222601bff1678952756d91429f3838666412a5ff331bd5c55fa7f2bfdf599c93c276bf5d0ef63da06eee95ff73f64b207b94a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88563bfc35680ec4ca135039651c4aeaadb58890da59aa0221c4f5ee2165377f9f6a75191d951e9e075e7dd3f7bd331e54d6d226e140771873d7f0736ca385da2623e92d6450f18e280706dc2903b5e0450b6c34f9c38c98b358ad673e9807d1e42870c8d30981456150ff2c60f80cbd8cc1a63159a8656f9198aa63c8df43f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h686e9edc12c5296ad47a78fc672687a3f71d2ac17f2d452ac3cb3aead722d2de381d42a97d94fdcfd6694dd24657e24f82e3c9f8509d129c1ab88b91939bae4535c0592e6c439f7e01bf48d4d428c69733db52c5846ffc35a41b1f5dd3bc4f78a1180ed88ed2fb602f36591222c1ccd2ef54d4602ede274f002cc09ae3809e69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69fc425de86df0090abc3547617e2c5fbc3b6ec25be41b7e997bfaed8f625731771487edad95b11ae596ed51303cf5136a69084dadbf66d068710c685afa1ec830fa72218549ad435427cefa10ac6cda93a3edf09bf294f9245d99ddeb1ac3bb68a5ca2bb1fc2c105697285ef0703702448a74f3fa64daac0738e3499369e6ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha99be7496dfd4f2e5b9fca9f9eac18fabe8fec219fdb420dab9e3d7931ae82996581a1aef6faa939109ca3de09b1757e5a3de250e2931c7a53549f05c6b1567dc9dc9e89ac0caa4d39402f7f5a11edfff3d3f553de05a7538f0b7116349d9f4dc1a897f17fb20134ca6c06a4dc38ca2a3dcc6f9cf2a3a8b3b94ec8c0ef0a1c75;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cb69754db2ca4eb1950ad0512a38042f45d535001b91cc5282994cae164082eb8ac0267f588fe70bc58d688f7f77050380ee67efda4313d90049a85a05744b329f4f18953dbf1d50a5b77fb22b147bf13be29713f40c4a2afd327ae11efb4e6d9e9fcaff4594e16df584b0dfa262ba25a11ba196a2c7c02806ddfec4a4ac635;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he26fb7ca19e371855b750773f48d12b8518362321e3f082623599df7e708a6ddf5f7b5c4e2a6158acf22c142c34dc96cf1555964be9cbe19771e328aa039b9f86b514aa6e7585dc70443c46b6c1b3d746c29f0d8d81f370e8739809b3a7f9c8c2dfdfe0648c9fee3b7a76e8043e818e08d27c21594779296675fdc8e5e098ce0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h242d3ab78375f1daf181717366b280c595d18345fe1df382046e20e8611f2fdde9a2b4e788cb6b5d2303f4937d660d0d3ea5a6cf1d7837b89c7179a444a4f505ae0f335b2b1a3909787847b881c6d79b4d9cbd6b590694ed70fe4c261166da3da57661964a5e825a063471ba7804427bffb945760b38e8f7b9088f24cfd62c16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49e13eb35d4f551c67c1aace77ea01921fb840c343e15f14e7338710a103a587c050846102f0a80999ded637fd42e8a902afdb9acf2fe2095c5c7086bd1f10e8e8b89e7c5ec0928a8c519a40e9109dfd4ae091e69bb38458f9b1aad476a15da8cbae417e586bf04a0cab553eaa13df6b7babb4a922f43ee06aee45dd678c072c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cb5d4a0f0ee093be08256af86c5bcc971ec3d1cdcf0e11ffe992ccae865d4568dedb660455a92a30527f39f9be2efe77bf0c230f7ab6fe758cfadd1447e19d1d5a3c3652f2c29092ff295a8404fc998c488e6cc2d9ca5bed0b2fd6522de95dd434b6f89a871121d54667ee8f929fe3e6afc76453239d1c8cdbb6bb7e22632ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7f425153748463d27eb12391570bbc80c88b7144299591af774151a9a107082d5dc4066038766de8ca0faf094594a9eb6511784c2b3419084448fd0d2738cbe2c8a7c4bcd5a89f5960de21360cc7038dff2f6af1078a6e0dd3b465b2ddecf391894740c9c96ee58b0d932d85606a9ce04619eebdf877be9c1fe0a20351c3ea7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26b3b373d0b52f9ac15ca91791ef21bdda48624f1fa292ac703069343ac38f59c29a3b1a3d5db54c8a258341ecd3408c2896ac7d283e4d34c04134a5a80c1caf16750e65db20a722c3fd0f12fe246731f2de3500137b70e9d58959912b82baa0b04186f85a5709223ee4b882b0d5fb3ede75f5e093fdb5339463c248dbb90244;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19d2032d1e87fafceee793ac9f907ed13eb6b1e1309105881218c7d1425f23482e08ca9cbf6d43094b1f0b250648704b1bb2d38c41589d6fd5add2dcb9192b70f1c45b6e846c78cebbe8f06fd50fc103afdf50d80f3d646fd9174431ea09b698b2c3ee869e27fa69efd90a394bef67943d5555937203692f8f619185b4842d26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he855a91f12b8ca9bdcd77d0e44f8b68aba0c7a34f3f13fa3a6c06e2f5ffc242b994a32d56bc806c26e3d5a3302e4a88565927f7e0c488eae87221d8eb502152f0907900e416506f84a4d0b40c9404765f4da4cd7dbc5299aeafd401dcf0657317ec8efa3296591d4349e0b328e446bd67e4d9c2cf0c0f6a9317970e7cd4771a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha86bb8d8a617106e1bcd9132c7f4c6853fabaec6b5352bbae949b58abf72b4e04df99db0dcd2fbca990597fd7996da65729041a3dad3cb10d7e94ba0831358c4aa5e28832227aa9204d3dc3052a87c56d0c8a3cf148c31a9043f012634865b13d7da6371199c9d33098cbb89681d6aa4f591c4c31d0bdd6b8fa244a4089bc2df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30fb4699ecc487572db031352d88394ea34001af119bc6caac6df2910e9389c49e546cfbefb4b513a8309bbb6afc66bd8b51c40bd1be5a6e48c701004df8b59531ff6e150e7e5350e2cdc067ae18e8b26433d6092d36f9c9e7cd6e7910ef6f450888403e90f53bdc63c865abedd6890997d563798ba767fb5611cbf80bc5594a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h372f76717021a4ed3a62218c0bd8e19840154e403c9e561eec14b6e22a7aaf5bc59cff2c3c53b5ef97490658bedd55abb4de9805ec3a2b063ed36d8ad2c9ae478156375f7cf1a21e9e51456646f08605a7f4ab897d9546d53ac8f30daea14e494ee072cf04d693ea61e96a4a413fe4896dd1ddb47c19dc75d9a456fa76cfca4c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6802bc9b53467e38b18152593f9e7ea10ff87ef53026ebc4a7543250724d43027186478f81c0dd171752d040c87341168ecef80f58efc3040fcfee122282c85187e006884d9607e4bb644251e26190815edd81fb20c13b4fd5016c7e520c3d7f6507c384d34f90d0597f721ac88291dcad0e61cf310c7dbabedd04e791cf912f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12fd59b54ad895bf94f7e4ad481ac5ac6da625c53ec86298029a9b58544bb4970f5becbade2623dd1098c7dd6109ba368b2ea726f203e6aeb88a52e5819a5a48d13305a6e6bd465dd636f939c9deb397fa15640b3185ad33742c83666cd26ae196f8ac5f6eff0080992884c6bc98c59bd8d2e3c94287c320a4637ac39e450877;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc00e85c4dc57df6ce18a8f134cee154c2cc9e209c5c4fc72aa7f3b85f90bfd31cae9175c39fd0e4e34f1ed85d71b681b348ed3450daac7a840c85fe9cdbf002a3ab6979feb18e972acd9158b0ce7fe955b0b1789c178f858f8442ad18255bcc51c488bd956e101d44d91a6b36f0bcd59ae70c16dc5642ccc3945e9cadcedd830;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d851600bd923040f7d0b4eb26259a891297cb63f53a614799a76f80bf9d9f1c97a072a2e22e46310d45258202b5191ad095b4ffb4911b49ef9d04f7f24fc085b2fc769cf2798ff6de54a43f3fe63011ab76d9105b331c6e501d873c4b46b25b5ee59de62f01f1d7872bb0e529818481b4ee04e46f27049ac9852df4c87dab71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h649a15e6ddcb50a096c99044d395324fe1c223db6bf78e7427d6dad9e98544a85c7602cb101529c6699aec83eac5ee01ad8b3a62f0bc4b9912d25434cbb0e5e22d295251fa931716d4c6d9413f80e467d51ce3fa6ccbe1c4f9eb6667694c876dcdc8292e044d4a19cc86de7304e487f1b33f745aff86b663c1a532ebc8c1631;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha30e01f2834f6c5b80a2899950cd5c5f4ee3567771c67c09ad44774c46343a48afcb62233472e2cd0e84424f93c95f21120d70c207c1cd3af236f82011d395448a959694621c5d997248808f3bb16b34b9ac254e1055518768d2821a287b8b3f35166894171359b512757a4df7f297bb6d1bab7ba8585a3f51d9259881276032;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ce1ff004a59ed0c3313215e4ab31ad6a568c9da65e417212da1cc9ed97c57aaa4e37f68b6cdef01ff8a10ae128bb4c741906480aa1fda8b014d46176bc661465e96d83c1ae4724f8637b53056cb80ed8cc9a8521701962c7f8e23cb509d22b154882518379ae8c86805f42702d987a5db6e434e377f3a2bf4b7887756ff2bcf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7daa7b10b31b4cf6c2425a18b81df96e90532a1c95ee09e0618a07d47031e0da7c221f1ded4d1947703587d0356700547f604fd9726fbc2d31ebf81b636980ae6dbbbf44be25a7aa931148372bb22ab6fb07bf50996c13ba3540f11d470b739cdd312e1e8579d7d052d543b27c5a1a22a59607f5eb40db033d605bed08a726e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5805131cce0ed5fa65d034a5b4332b2c72775f07541820760c6456fd9a6f010fc7060782533ca9384bd0735f26cb2a4dd9eb62c338531908cda7a5aa210c3ec3c00fbe6b312f28fa134ff8118528a838aa9d2da116fccd78011e9836c3fc3670d265086ddda3c1388f3fe8dbc1b3272c83b625c67439cb35691611248afde865;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53efb6dab6a2a9a315adf22595d965f66db25642902df3f4d0e956897f62a3b1c4f6d620824798cbe454442cbb3caa99525f3feebe2b57e092831ea64791253f661181746129a40f95c6468e093b125ef4c12e79e4255b49cfc3e15c7bc8d2561606087eea74458b2fb035cfea08d3eb96559b721800217d0883967d040eb1ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heed7e2b1f1efb986c35210be8f0c1b1da1e2476de71709d35d7aaab305f53dcad4b8a0facd51ac9b5e132dae163412b325e0071da5780162ad35a825ad0315153580a4981668da7f4820d17f4be6808b85d68414751045790e303ea60e102decde135f1ff6314e4e05989b898cba9abc727e4c34276b96965562599be92998e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6024e3636bf181a2ce1f938a3152d2ac1189a5676050ee267f935ef3d91e75e12a7fd893c5da718c63403c52e2182308ebfea0d2f90e43c818c4caf4094a20871986c4917d8e00b3f414ee0c02fa739f93c389e4bc0311ad7c6e13cbbe1f267c573ab16fe45635ef17fa9d331dae4aac57bde16553c0d0c526f7e120c796a623;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72cb9407f21d9a8b0243cd83e5df0b90637e45432637a2d8e3706f5e71097dd8662605f2a147c5fd106be05a6c3bcd624459a4a8f28b754e324dbc168c8a5ef526325faef7d2930582eb45032d05c31ff60a2fef98ec17e8b3043ccb2294151b0cd8b56e6bbaed2875cd24852574e8e2c117643e077f18449830ef1e7c2a917b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3f5f33d78974a962fd1e831b4130434ce0c0200309af6232d6cc951b7cca6f84cfab391e9ee83739eb68ce7f959016dc30c3f4e6005527f88befa811dbef31b242b9577e26e3a62ff8df09060ea2859bdb282453d30e00f144d28c7bba06e1e8e217f46e57876698f491e6fcd0cf293bec4c3eca0c21063a4b844ce2a1703ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb4573cb94ad805abb4a5fd840ad166a1e24c3ff1f26a6d570cdb709d656dbcd029e1da0b54118f6989fda23ad001564d4f47a57fd8dfe22794974c29572c289fdc6d2c0bb2946d53b7eaf24764570c858f4e7c2a7b5fe45883818b4f4ca939b8f8f910dee30cdece8d3c8d6dc922d10d4fbf5825fbfe9b19831a5a564bed453;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88b57aaa9eb28e5b3b961b2d1724227a5d28f3f8bcc4be350e899f1f3da7352f2ad982a7ff5eb17b46a281f2de72f634ee8488325adb804398bb495edd992f6f648c42ae0148ec84a10fd6ee4a322905677fc0ad637f9d85d81781edb9e801456a114aebf9f68d063f693c362e1b28e323269b6b6214b4d8e253aac6a0f3c8a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e8f33be7a16d24999c31d7eff6916ba7295ca903c01ff1bd1e9deb92f430b7482ef399ab6b128003488537c202bdde1c05b82ba5e6a10f6d0aeb8188e92c559a13462d7b798f4b8336340524012eaf14cd750d1407ee9a5d8af9219a518696ee0bd0b3d45f7381041a9d75f7b4eb3c3a331537af8e4f9da6eb273762ce72ca8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6f18aa046d853d30c4975546233b93276789e45a20e4ca40f531567a99419b9dc98c3e3322b458a3a2306223dbac7e2962bc89963df76e9b883c16b6c671e0cb8286ecaaebaeeba3d75228c43ae844a2252f42bbae9c2b691ab9f8ee4aad8039aa0bbdf8e3810464a7833cea871a58e811aebe03b5128655ce56cbdb430b6e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd9af4c929be2aa8cb026264e2c47f694818c18a7c88dee4843f1bcda291568cfa34deb7ab13456a83697f37ffc029b9f2e8111140b5686567edaaf8fad8b31beca83a4796708cc871c7735f693b5c8d93dd4bd9a932b93720233e29de52ad3d60047088cd16d2178f2c9a42f49803a97cab2eeb02dfa7069bca9094391c36c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1f2643d73524352ca6183694f630f10072fc7a2d33812a07292bf8b3d43e87b4b8fa599fc8d97fc451215b0a81644b371521007d81870c938d6df76fc8b4b7ce868e4d33cb5871c72838f85a50bf808492cddb7a3a082229b7ab84a2976c596cb0db5d97aed354af3da0cc0d343da05142abc59c7841a84e8f2f0d42fefdf3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54be9416bab3aa6968436e5cf8715863f767e83d53a690883ede1fae7602ab1bd5367b8512eaba9db95aa71ed28f7bf5b0b157175be9aa507272a174f8bd81c03aaa3c3bee7e6c984f5ae7c7b4f0d35f08ad1cfc531c9f383f17ccfacb03098a4d08454b5436744b98efaf197eac09be1282236360064593c7c59157a5092c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd29c5d4cd401bf8a56b5616269eb795fec6a95590997783d98ad9d3264ddf3a16295fb4c33a6eb5948c7c116b4aee1f20a6265c87ed9d7f944789ff5bb2ee0300762bb454117eb03b838f36e7a4887ab87369975085b311f97aff51dbde440fe826a92ffc06de234d22c234aebb16eb0309905ce64e9de7e86c6ef79be223f65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d3551c0429b63419e1d6b3bce412c75d492f630e8f59ad15c08be5a0e06df02f9bd54be247d79783c6face207feb133b122bcea274a3a5820f04e1907b28ce30dddf8e097604fd11210a287aa9d24e00c60e0e565b209b6dfd24e39934e9ef24add52acbcbfbebb662efa1bdeddd285a7585022466f36e0d6c06165e060b6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c97edd1ec3f9d0f40f0fab2128faf871fc63c6ab4d90e806ae81dccb8fbfb8927df0bc5a6220edf4a1f0bfc741ef3bcc27cb69429a268eb06b2544315f705b152e3eec88569bf693542e6e687659ac0a95f08951e25f220dc365c77df3115e0d8e29566690de3b55785fc2487dd3b356b6817b09cfbed00162ad0cc7b1dde85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h491dbd555ed0ab227ae9a98ab29f3ac487d9886a2aae90cd7287310775b5702c5f5f24a7dd87e88b10f340d24aea201fe0be314338c6bea5e82d627b278f2a0ab639091f42db752b6e058dfd5851c24cb361061f5def44fa84066b08682db6fffc488a1a21d61f265dc84460dda1b61232cda7ac737f72fe211bd4a984f2207d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a90655301c9f10b117b7791e07a7c77a6d33f944207a44400d6f65ce125163070eb2625d5b91937c1c87c5426f0cb95556fef966ec4da2ad7badcc38c6e5e9b51c15443d0b870943530a47faad9e3f5d3f7d39e60aa98030aa2115df8573c81f8fb9e5659f6f0ecbf97bdf450871f6b273b42341ccfc17ceef1174f4e6f2d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ee1badbb35c7a508c48e1ea939bf0493665e1e7bb8a617ec46c7897fe47f0fccede0c69a6e480238c9a4be658c73bcfb35cf5670d907f98cf92921b6a8dffcd15a13526c6f61e4515f899d146a9439af99031d9954ef56dbaa7b8b3847df097114726694a7e737d10ab2428b9ff6b4fa78e6956901eaf68b765058d3f5a7e04;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8558cb56c868a0810d8f306199d2e0fff70a9e7580bf3b08ba0acbf536d5118b33555993e0357a4c651144aa79c31faeb79bcbc9745d2e2717413ac66bdbd1a8ad057b69e899fc6c5fc0992b1036838541770c4a64b968460eb5450f56ab665c2b0046d4a7363d30df3f39b035ca51353d06636e2a6014b983c3207b79757009;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b0684624fc54b9875957243f9e20d406c70190aba3789dfc7b84c1835852ac5d45fa2f844298cf4059c25d63d8980ccddc368decdaf5ce87d41c7fd737bdda611d17f69e46d9f01be913032d896b4eada3d33b4f8f9bcd9b15ae9415c3cf8b3255b5786c8e8c4f0f62fbda23f6cf3e93994c59f2aa6e00be8ad6322f54947b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d2500d6d4b9bb2570298d5e7eb05632ed946d295deeaa4e255e6a7cb9d96ff9b84b5a0144344f41e46ab95d86702e80fa317161e2ed3906af7499852e1a0247b5a07a11f511f4bd26abe89bbee003c7d3ebbcd43ec46b86bd35472662347f7453dcc0275c1da4b266183596478ef8037fef4bbeb0a91f5059cb8cad05194bf2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hccb24ae6a7b5ab4bbbc55193520229e97f73ac09799b5f33a40e2449d35f21469b84e9f277ccb86d503161c783c9e03c026ed68ce35ffef15acb268a62b92e0712cf2daba90a8771422e9a13c2f2f5ae0eeca922c0036a7f21b4219828b95bdbd51e09c3b78efd443f520a1446f34b920482b04ff5ff1357707b7988739c2cda;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd46eff5bff198691fe01ea8117ab01c12545044bbf49585c6370e4f7d17a86f7b731566e9147604a17cf29b37b36396aab4fdeb80a0d576ed638a18e7eae844ad344749f8159dc9808baebda38c75150388afda9807dea3425c0f8c9463c500349b80e5285a2f0596db130031ed72b197a220bdd0b6be92845012feec9da3e86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc314b9c7278c3d41a172c6e88026df099be6fdb4854f52b58eda9224fc9033e8732124d3554cafdea95ae47be0eff8faab8080926ded2319a8473783626d0d29ec89bd003b14e6a97c61e7a834472b793147ed2e7458ae4cdc515b6c7b38b4fef8988b2d5b685012c35254c356402d87fe68fb229c54d1e3c617f3ecf60082ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8aa1eb20296c4b6b4c44affed7c6f891ab2565a5df8f4ded5ea8cdf397076c5bc090335e975c8c2c75dc92b55cd2c02f1cb625e02f56c8454ae54f79a77cbc25bc35a1de2896ec26ca90c0bc531baab018ac2702d286c8650ffcb29f4fd25d17e19a623885ff8b57e924ea5ecdea9f6a457b6d2cb6a0e464600a4677dad2960f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1cbee8a170590b150882045946c73d4d9f0893c26fe282c110e0843b00d9ee4e00d290299c5b5acb2070a98595f2761fb5d6b1f46ca11804d2ce87c2c22d9c013fcff0ab3b879d260df563ce3b41323d1d6d42f6a6d15f02d1cb11efedb965a72799197c1311ad39b6d89fa77134d7a31b8e611889ce42849f183ec3366eadf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedda632d7fc6414996c014e59ec1540cde3d9be2e89a15e785ff19ed7e816151dc5d76530849100d0fcdeeade0f4b4df9a22b926ae627c49e1472873d72c354926fc3bbd4ae4ff83164bb373f8a0588c42a33fdb440a8fa35ebc482cfa3dde0a8ba1546d9182fa1684f337b964daac656f7918017cce2a06ddc7707da4935b5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bf0e6b99197b59a6a64c8a7abd03bc116f3599fddfb701a4d6c28c8769a9ec65879bf0ae780d537bc3804f74606332b307639814b308a2693c1ddf2431072175109150a4c63ad2141e1d70806772b13b20e9b11cd5c7fe3c4b420e0d85bdf77732187b69ba15f8be218efed1c17e8d229e467048c3929b2a1c0e91bcf51d0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha807e5757cbb7502ebef3e62b750fd7616186004c66d4bf8c5582103eb103f858d388d526e607fa45b0b6a307ec8e235febfd228e2ddfff0a2c7f13a91cd988e6cafa6454bfcbac6a9e8a7e4a7ac9856bd2914cbc680ea702ece381c724e16b11114f4dbb99d1cda9ec5a3336aa7a0926f06835ac77dfedc8f94ffaeec39dbe8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6878c619b97844846cd7382cf99987f9706def770f88273e0ffbb734c10b697d10faaf40c3a4cb26bc886a9bb4ca758c7f54db375b8b8dbea403e14104a01b3ab9cbdd621392d5d07658c39ba2423dc515aa10dc02b9979b1bcdaf536c52963dd938fe412f01c47017e4417ce14d36ec6956f0038a449e0966dadb2f3a733ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71dd07bd92320ba6ed5c052af280b87747d6e4fb5c546303520f60223fec65d69b319eb071ebef2ca4d933767407fcecc7e13c0b688538854dba3db09b70d82e732eea86e903b7978cf52126beb4f02d8c80a41728be464ba99eb987d0c21cde60a5ecdea1c8c743759295728e392b1cd89b4bab14c120e7124b70ef849b7dd7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed3cc5c35f8b34694e6088d3abbc2266f63845b7d9e45d69f2f68f65639c6068b95c997aa199c8c10e49c21af1388a81183c20cd44d0c8af3926567f19b3071beb3cf0c2b8cadd2ceed1bd6cb9828182d7d46b99e7ab084732fb8140f90f4468731a350a205a82d397c59802b7bfa24cc1de88c62070f4b9bb78961d658e5965;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf229aa68a9a170b58530eda66d5326385a95746c12ce353bc112731b0c0b76765b787fda3b3d5f2ce850d8e4d8f901479441778ac633d05cc56f79bbdeaa22f336151f006f69b99ccbadaa3cf79b83a1ab95fd2d6fbca022676f8460461acd676f4e132ad0129bda15c7cb2c3d2c3dbc145b013e7b4587dcfbb2b263863095c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3adbe085795ba39375eeb164c60d8da5a382e4f9e4a2645756ce51c92246bd99a3e616cb8ac80bcb6e044ab5bb7e977653655e7efd4079a5954916a901e125f9f52f6837196b77f683d908dac3b52a62614c5e42c14f09a7e51f32d4ec8b67336048611442b1a87c9825767734f6876b9095148ef2c4ac34bf79a3ffa7dcb506;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b8a259dbd1815104492c3a0d93e48d911ec4702e5a743f90c68acb3efdd1ed3b39589aa4f58432f744210dfc3636b0c56127e6ef3ac6f3c89038909d597f05c9b284797bf9c2a1a916f1e0722cb1580d4d31594549fef53339e9849810898e5b8c722f17de179f78cf137141c25c9a9654b495c77c9104591ab0fb801285644;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83e35f742a8346224e7fe00c5ff1dd6a3f4b3663cf2a6794ea089159a50f724a96864d44a3cebe4e17ee13af9ceecb8af54048a1b3e5ffa14d3a0a8d9a3024765b25d884602b817b6c2e5dd6464610965b7542e42afedca3c60a3d6834e67a2796b2ba6d1f92e4ca7838fd8a926da44980f48d0060be1a9ccb30a8a3449285a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hccc0581bff942bee8b53c51809f19f4404aecc6cf07c03795fd6b980e28590cef8c4d5908d4a935207fba390b907cae86665c40485314bc8015c5985a77f11c84243fdd63388db5c9ce314b396119fd130bc4f2060fcd60e0e92b170ffa93b4c27bfecdbfc56c5364e4278051dbf75176d523afe3bb738d61f1147a495ca5a32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf28c6f0a910b5a8f5eb192a5029e81189afbf2b0e7347aa376ae9682d3973d88d0b6863b62d89ec199789b4952996c360a2988d46d9a869e030c4d3fc1d2704db582e123a27758508591cf00d8d879d402ba3860583b8190297857a1c0f4b84069acdbb3095f21cac19d5368bfd443ebe94be97f9c7538c39646a879904c296;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50b09075a24160c3d2bd19be8e04e374860f6bc20951d57a9aef115f424eb03df6f13a2ae5e52b8f63b9dd8b909ae0e965df9dc236f3c72313eca7314e484a923ed49c4d251cead07a1d4b09a67329bd8b2dbd7efb563584647e67f598035dc014012651549c4533e520702145f3f6e63e93d6d72977a527e7ae9300d845617;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d7c7fe23429f5c383f36e347238f5bf60b5e468794009290f61a65aa6dfe96a08d7509616a5434b1db0c99092aeb60ed9bc52e0321195fe9f5fcf83da67a832d9e25d5982ebe13956c796096e3a3d39022c5afffd83cd0bf186d22abed1c7e851e8dd98788e620a3620705a54320172ad4aa5a828851f16ec6a94f61940bd46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0ec26d4e19a1019f812fb505420b0ede6d6191e2c1b8a8b5ecd4da35a67a40880cd095d265aa2a0cf45dcf15a7ac2dae0d4084c13f989fc25cca270e8d55d8577351935ce25a7f326742217249f6243bcfd44ea135a887188bcaae6efedc1c3ba7af94ebcbf2a6fadbe16c9534ac8af9e551b47b2427b5564966d3668f3976e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6105630fa574a175b99ff1755ea908e24596e76aa164158e71f8789e67f78a5dad2900482ba040873f45afb33ac95f440dfc53e092efcd96f69a988553f2db2a68a4e2a1f7f26004d483862dbf93cdfaa84b26acc7ae2db3381e86bb9f9468eb1a5f50f1bc9199ff61322fca787a4f77b2f2a976ecd7babff536951c80dd7d90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f3e3b618189fb792d81fa764ee56a995184a5127d78c239a3746b074a987c622a9ab3fe9ae8aa800798c50cc054e8c49c437547ee59a3cc64f9ee4f9f88aa0d9bbeb7d175c455f3d10d579bf014e600a1e3f9e077b2b86b5c994a503accd8a8386b5bb12bda6730f7ce7c8378d8bd50af0e5adf8c5785da13bd5b24dc4fc23a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fd212a5b50ee160438cf21170b8241908b1551ea4825728258f2febb418d1b516b629704500399630b47dcb05da0c6f3bb8a436f958ebe3f355394a8247c82cabb7fd933d40fecffeb75e91b49c5b382d53b6131b4077abec6d8e8dfcc878c62d9ad74e10d64d190a79d220b2e86fa01bac05e0c8be76115ea2aff19450c583;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c26cf5cdfb9162aa0b194df1ac34b404566619b20a91d99f3b48d29efa6acc17505ae34178da5dec0c8e7f07d3229ef129c699ee4db46960e93e33520ea8a4944c51d84ec7581e9e7e106a6bd822835d63e1bd81d51890af8c311e11adf200e71a08e308a834115076bbae698be326243f9705481183befb96ef136d523786d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce4f3ca94a117f2428080daa5044fc6e0334869dada2a830ea62a4669326c6b86b9508e31155041ae7b3e0dc14e623efd0d26a1cf84cb1cb10a11fc04e6dfef60c463bd112bd9749ac9161f211eb55e226140add7df559921709bfc0bfcd1d313b9584da7a1f75b2bbea36289e7c965542761d50acc1596b217fcbd71a0b7d39;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3637f1072b5d3f8a992706ba9474b1b8fe6bf404b49a9b53dba5db1a005d8d51c16cc18a3f42668cb30a9b53ec277ad52d3011982b8b42b9a299fb414a071efe4b347d5797c2df874b8c9e84b8e5e43223ab73e3f347914e52e99a91bf68263b69ae205002972dc5df9a32b967a7fac83635d2bbdfa37b925a3e9d0d09cc7ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14e5fdcfe5fe5b280468b08003a3f05d3bc536fa53d7f165feded41a2ae89278ffc320302f0ab154de3c8478b17b5c6a522f173493c567339bc4a268972a7df0d48030082f2fc12ecce0fb893a2998e78025c37c4df6ff4008e99366a586a5ad1d90f3816671edfd642c94def759cc82e2096912dfb13d2f40692a37c55eafb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb85cbb5455d419a14da824f16fb3123abddf46e742ed886aae6a31e047c6e45dc1048b86d8f0174c81590ad03d2459b4077e0c2dc94d7f34004980ec39f074ace5eea0cf722b3ecdf97a4b12c19a884b70e71a17d7fd7e70dfae717960a5163f2802f202691e0f882f8661addebe715ebd2559a0774d33c3be917fc24981f16b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2ca7905001e2e8cd938634976eaf6f08751b915b9d93b1ab19195796ccabca93a1af0e088493828ba5ce126d072f4726517561235f25a41f6f20844184435b2a588162e8f3070e4d2c4e335cf9e51c4025f353a56e5dec08a128d9695ee851425841de314f6750bdc1b8b5fa7296f72bb853a86aef5cadb67f3afc221286b38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7664e5892e1c16147bb229099731ab2cb29f6f4ca82ee94c105340308badbc76758620058427c5c40cb5ed4a5bda75cec18cd630c2d0f1af04988f12afe2695c12343306484347d281ac27a13c0f7b22112aec18e416bd089e1d392958c76f4b1d7856b147e453dd52c94d9b4de465abbb4177a2a33e7803cade079a297b9706;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h615596e7774d900076c5b0604106565f2850ecf0a660167f7e05c237010439f61259ca0d6c043c1032feb47cb300519a168299a92717c72928c627fcb4b90c4b9d2c0995981c0c4af6a0c2a90e1e003a10282f12a7569e8b92363725e744f2acb67c255594c95ce482771b70f5fbd8900cb1b459df234e684ca6c44b02443396;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a54523700f30ce6437a58cf47d1253ea30c5738752ccb7d0f23813efa2435ddc20d617e4c02cdbb38a544208d993732ec6f459ed5f4cbaac7b4bb86da20150fc0b318172637d7c18fe2626af2fe4b97985e49731b46cfc0af3317e4d25bb948cbd6b942d02e6c1ed734d04102637988c13a2fd009b4cf5a014ff9bca6e9dda8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf73a3472f58740caa66b6f0ca3c800e5e2d1ecd6c932507c68de6cda8e65ea53d7ce4d52f86362e9dccfcb6455fcb32c510de0bc90ed77e32b1f6664b1b2dfa4dcf609790a189a4bae02ae901f8b72db94918937aea992d25bcbb821cde4b6981c78cd6207e93b9c0f0e493d31140828ce761f744b83cf9f3a36827607e28ade;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0203f6c1940483f1d6d56611037eb489c44ecb0e17b002da552c27f5ae1fddd07e2aa3fe6e2131bba797cc7b2e8759cd1ac17e312292c5ade7e0c200fee5adcb72f3df3df8cb22a078c2a25eceeb2e6de61fa3632ceb2c502dd819ce8523d10bb4710246875431eee4b99f39b1c61ea388e6aa35bc5923fbd8f7533c13bd88e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d412d2712377467ffb1c111ad304ce6bebdbc100ad1d0be5cd9e1ba1003ac7ca9b202bfc859f18cca5217d4188c9546f08ee55d98f14960c6550e4d441723bac49c68b6be5337e6b3d6536aa2a25190fabdefbdaaa791df16c5d4c849afa98f2558339ec15296bb974211300cc5270e936b47b257a695267fa017c4a90d7b36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1895c6f95bfc9311c5b186c4c8c4a57c8eae06df1a1f2d68f79dcf9439098530099ca5d6a5bcdf1b21474651c7572bf0a1008a56822df9ee6408d5197a052c6d399a7df186b2050be78ab7b67f1a2a1631071dbf05f87ae52f8a10a197c000ab0280677b0965708dbf45f52edbadd0521cd904bd695aadd17e88efe48e901e34;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ddeb6d40d63b7b9d80997ce61ef535bbebe3cbe76faf2ffa469634bed2c263066ac8fd5657a0a5439fe443de1fde996ee6a43f52fb655165369d971788d7477e75adbf645b809b4f4f315c9bd93f70f128e4c92275814416680121abeee54d2381291cff507ab15421303ef82cac29c1c7037387b077d0533cfa9673bf72b09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17e0c1deb93f1500ed1684b5fcecbd4f5c03c08a5cbe8f347ed6e20c6ffacc6d2506de94b1f83713a71cc2852d5abe5483fd0ca6d392995c8afbc8553aa2e7cb06bbc87a9de8c80750ce715c0de1224b4b230b2a15c4375a94c22f345820885d8a5bafdcf92830efbaf7782b7f4b1e19a5653edb4fa664983f94af4e08470191;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h562ee55da3480b0c93a5f5664f562556a68232762e7a411a34056076df7b2d81e0639a353714a37e27a6de547c585ddb292e8b252eb059c4e02a6e681c573e600e5eec00e2abc11b6b07b23bae3a877d7a6f4437ba1f823574ea5ee4c4549ff791c1b06d630528a0031bc90a630268a2f59e60a05f658caa1ec563333c1a30c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7cee20ee803c990a8587abf98a78a35e6be55d36375e3e8b255538ae86ba1a25c5637822235c38b1f196d6661d767275607f64a4e8f5790ac5fdf745520fad61fe1221cb37016e538a131d182162c1055f7a6dfb5e703ebd5f1905a45c9050044ffb809552968161fd68ab043cc2b83f4418e889967da96905891eabc6d67e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9da0c624379a977634664e9dc7d796aed2e21fd69c1e06d179d7203565b909cb01d8e4e393128fd446011b856a2366027b041be3f8c8d229cf8ec25d1b6e7ae157d29aa9b270daec9d69dfb9dd4c71d0208d2d5f71d567b4caa3eb028b9fd0317af18f6f7db047befd82d275538600334037656f7370d377ea1f0c715cf190;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2766e507fc20806655038177474618b3b67bc4b9cd302beeb549d8e28cc0ab8db1ea632e9c7640973f73bc50185606bf5f54940a52179fce051fdecce015fd977380733196254d1ca77ba81ed0bc2db3d57de019117732f2f6dcdea0e20d9d4770cc75f92d1615079d6b21623fdc417cba9e7bb58f6dbcf098a932e916858e4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86494e22ea1a008e4c7757f337d17f677f03decffd9c8be43cce2c96b4a7f6617b9172e99519c5e0ff7c87b117311d81563b7dd2b8ae6fab8f04c57d30fed62f745a05d8b91fd752b6610ee02d96ecc7a74bcd0144b3971fdeb601d66b20123fba278fb30ab3fd217f3354c635dfba3e5a05de0c5ff0d4121eca660aaf585a91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8efed4eb96942060b57cf0af9df9e3559f21faeb201a477eca95f658be35799e01ff0a722d8675eace0e97e85b1b3268f5e0254275de0373dd693448161a34f3eaacc572700542a02ea38012a7ff3280b1f05176ed6e36a8b5cc67414f9b7f5674a77a3ead1d1224f6de75283e6aaf69caece34dd9928fa0d5bd09da3537fd8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6febef0a1301f65d82e38116455d9c677fdd328ddb494820d2b4593949f7576675d4b65af8afa83b9c79034c0e397609a12ef03cb10ae40231bb2b03ec7472c19ecad111e702a8b5ab42a070cbbd8f3f3784c7eced0d34d1f799344dbf1fafaea2174b893d3f7f7f18bd5a860634441cc170fa3e7b1c128d19f6f57e44c597a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacc9fd92cb6ae406dcbd5d8369ae3817b9d6084734608fe8d6563fcaa576a4885cf3374158e30e83749dad514b22e3a3a961e812199a5b8cdab18e2e1c39c09faaec9b5b4b1c34378fce356699ef1490b82c099114e1da3cc7b226e68e89a7453e5d6989b49e7cecf83cf6f211013a2c3f6378c27930c38e4141d2ad5afb30a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h127a7cc92d7434b390c5a44f077c71a30e401893a7af2fd2f37515675b512ee052a74498a24aa1bd8c0ca2ef2a821103fd622335353bdd8be2e335449a232e0c5545e2615540139e68b380fb39665dc5d1f2a67fdd8602f48b421e8378f468ebee4f045f7badac209ab8445abccae622ee1137f118f4f304aed298de5ded3f73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36f0397e0c9f82c7ffd177c2e87fcfe39d7b7c2605221dd0344ae132293946894808467d16c4adbb991c91e70a5d27fcf9e4dbc7d75304ec06f1c16435e32044d9483815dbad447996d3b3cd3ab2d3bf622f559784ff0415d273413f38e2a9389b0ed3a133244e3d8d2eeaf5ba708606429417c16e65fe949eb7d5b21ddca253;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ac9aef13a9c70ef4a5243e2b72fa89fc22d06b30ba0db394a5a238fb7a78024c0b7437da1264227e9bc3104081c5e0ff67f4fc9865b5ee3ddf16cf7ff8d948902f5c9cd603e286e36d2c41626de2f4c7c7926b7be7578f2b1474493f9a7e71cd8393af756e16c2e483951deeddc9e99b4a25f54ed6116718425b11b5843a295;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h350bd803a545fff59bc43dffda030d6b4a1918fccb07b91159b863e4c010eb7744221d05dc321743d4b35fdfa246aed3289c39de54f6baad80517d9b5ae4f50d630153b022c0f68e95cd83e3f078a7a0031a20587436821cd015ae27a5b3217e3e759262040498e7a2806d0d80f9818893fb2dc8c014addd5ae83c294bac15fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96a7a28c7ae63772edf5ae009de8e97598a00c4d932bd1b7a19f241eddb580fdfed0c95dd5e03abbbae96e4955e7d611ad7039dd68a7e586a6b61e2af6d2b57f9fc83eddca2e1fdef1a90fd970609273a1f9489917a3be36d0e88549f9df1270c2f0db32026a8b9abc00d9d44c176874f6717cd101bfd442184995e37b63a48c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5445bab75b28b625e3f41c4e9c302c1ac91c5d5cd90dff4822692651a1d2aca06015299d04d16fb11d5bb179d3e5665a3c50a6ad499ef4c382c3721e0590b60461acc8d71ca79d27f29687ab7fa767af5247c98eef25931119e2e50a20f12d128a2f641a7435b9bd9411e48407410605fdcb917d9734e7f391636e4b056c280;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c307f3f1eb25de9536526aac8cfae64f46d07488f8f6a4e470bc203d174a961ad8c2415e6ac7fb2fd1b5ebd724738bba9c3e9496a9ebe37f1c9ce650bd69af8f8f9afe79633813d73e95735af2a6ffe5109f2abfd8dd43bc678bf12f92e2d401bc9780e5cc5088b816ba74daa8a4150eef952c1a27101a73cf2f6ced0273777;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52a118a5a3e6c8420deba96e6be7253320d444b8423ae4cc00331153b6991b261b794b1561a154dd631995a5511da3579fa27951c949736ba0fcc6f84f91dfbd723ebd2c5330c01963d823847c10bd4ecd993bf6142f2eaa07e2e4429c9ae6604bf67f09b04eb9b940f94bc1d1598206e9750a2610128197b8a714f9df445fbb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41da25af7355310847fa5105ff09b7013d2c0a35eeeea231ea94b6c046186a4883f195bceb4f13f019364ea18eb7e335a799498f9eebd3f7cb24f01ec2c3fc941ea387dcbbf1d69f7dfbf16535c6489f42b14bad960c997bca53e848b3a79bcd3b0c92d4b53a4fae9f7f34a25261ee6eb891eacb72c96228a801c24b894ebe0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5128af859a0d0763eaafc67b9bdb2ca2697d0380264d8376938902b08c78f8f9a530a60969fbe3f13e1d555078c46b514a5d282e4e3186f2de77d28458570cd87ba889237194ba731474858b44173d856f083e53b5cc5653bc320c229d881812a3556a93b117fe3436891309087432f68c4416aeb2dae2b47931c7d56280d25f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf64ed7425323ac7764a2d4edf4ed0f02235a40f352f674bb097c3393d4bbd7be4311dc04bcda8d3455bf0701c22ed08790fa444afbec60f3132e0ce725b96bfebbd498fe939414d3ff70968d7db82272d38709d12698189d785fa48a03ad962fbcd3b646c0a9ac624af3a404baf058481302ca32440cf43e8b2616924526fe1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2670753c15184cf0090f4b0c2d0f09c485737904cf83075a9ee187a11e673bbac533a02c9f6abcef5c10a6fc3abb48016bc536b8dce390f5f7a04ce799cf190bc8e808267ecb411d2423690ed92fd97a7184ee690e484b14ea208d78e3b112f81e2e857e8cf1710bdd2fff817c3d95488d17ed8231586039f6bd2eee2643b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8791bb975641b60766e6f15effd72e3fc1bec6e6496d61e8a48ff58ecd53b7a98694ee0bfcc2dbc2a4ff40fcba2c46effc1d273901d8a9c8e615b4d260590db204ce45b6bcc48d093d26315f68c3719ca8c58ab533dc0ea5c72e0493054610435c44ee14fb472cab0e42924928a266bf16e0fa6907851b24d2e18bb2e07d9196;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf537a41c59b63a5ad0a836c4f509112477a22775b25e5d1d9c362ce09c01fb08ba585989c538d1e29fc3bfb19335698683de89ada6e151dbc2c50a3c04d2248e76c1d547be131bf1cd7e062e1bdbfa3eada28d9993f8311cfbe2deae96b21f56ca0d9598024ea18a7283d8a8e586d9934eafb9b7e278cbca48bb1593d1ae4f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0047f703e887078b6195bf2cb28eac8aed8e9a19fbacafc3e42b78cf83887001c001eec6252471e5dcaa19237b915d905bd49e3d30be4c1770c9f3b504f6cef30689742c4636fb398d8fb81b33388216eafb8d867b3ba17a6c9489cdd54e0e24ae5c43f51cb17f3943c62d1e15523a29757f73f08904511e068f43cdcb93449;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ec24d370677779c70ce3462a49636d0a3a9353cadedf93c16aa3613e1f942fe99fef23169e6a72042f8ae731d911e52f0afb7b9540bd35f2d86ab2d3b94be5471ead4924e1d32ca97d5a6b87aa8f69a6847be32f6e3c3ccb10cffc21c5feea2e6f457d9a75a6e2663c6d903e9f3177f4b362dbd204d651fd7a12f797c3134d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f6c0701085efdec086b63b91371ce433da92038ac80284e030e67d5100eb6aad54bc4de44d1cc8d0bba6cce57d6598bbd9ed0a0dc41137e7e436ff4a30bebb21c392aa8953c370961b756a1fc291171467001891a9d207130834e460eb6485f824c2fea2643c9e8c6a38780337339ba276b3a6a8f32744e719dcc028c98dd58;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba24192c88b1bfe9fb7d60d2403407eb55e4f0914ed0f4062e29549349df90330af5d846cfca12f6fbd65824e402d77c167b7c4d7b58ad0599682669c4f035a5121ac0f126c7c351cea7e4fd17fa44ff83eed460bd44ee833d96e46a341ecc17d6dfe9c988d288099b2637e85de564e1bfe817f18dd8348caed8214cb8278366;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h134f74a80cc1740f3faf0f72fafa6d41c1a83b01168f959fcd5a81b1c95680111b0246f3401b514bf27d3b2c5c09d18ceddd55fd44f36b64d3e1d0180150d5bb09f6b59b36aa122ae1e9719b37d17d9b1fa5c11baa47df0566c9076935df32744b30872a6b0a553793ea3f1b64f5123d14b6660fb36d02269e81cfd6f802d9a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h546886c94b8c91a39bf79dff6c165105d864d8d2ca1092f808ac964ed056b3d9ca3d0e4815fd3eff23a9d05af4b88b59315ee04ec7e4adfa54301e3f83ef797efe7bd751f72d192758f780c2a378b06152c6cb625560893343c0a26f2943fd11cc4691028db0972e484ea10b21435fb130b3b5b8b5628754289749d8a3208eac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8b24a97adf3616f231c48aa70bc4f06b72608057c6dade739e24268037de9c52c774de2f364155d941ba3597eb7b8269d5e8d48c6f7fa46468245a8f20a02fe5e07171e6323e21fca294d3733bffd218d538caf7a8735c01465eeb8ae1eb17dc298326cec1ec0f21b852291139ce4a6ef55dad455143be2ae887a1bbfd62106;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0f90113a1944bb6e00357037473d3fb589bc2085a37007414bc27f1e83f94ef33bd8f1af978e2161e81e3e0ab3da72f14162102de769b974c1e1e978fff1757089c1feef17dcde3ba2de2e344936a6bf54d4dd3a4763c712a69b0b1c71052eff6928192779b1172b5c2c35bbb81e2e8d74ae82e4e7a10b544562bc13f61a282;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae801303a02d4b334526946b81194782f2a05544c52f96103ddc6f42b69712a1dc7df1560dbf8bf12ed1029a61ab7a0a9ae8e60f4c4949c39e9e2fcfcae21d0c6106c63af150968f9a6203699c8cc8677c1044cb2745d287b4d4c058013699cb1d9997903cd9047ae0e200242e5867220a48559bac863e4e181b3ffc708e9ee8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31662d77f96caabcf6e1e674c587201fdf6cdf4b7fd1126a319ba78d8ae8d71bded39f2c0312ce93857114c2d0ca499931d9ec3cc3d90bc4ae2e709949db3f5ba0589b3da3962ea06ab93e850e1b84bce5e93809010a394e96971c12941e24b80f0c19415d9a5266bff00496d3d5b9dde01650aff8efb865bbd360d092868ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e3df1c8081c50e025b6141b5e2e50bc4ebb799f61e131ab4304ceec26edc9452e5a688eda038e821cc6acc8334636be065136606e4417c47e11e4cb3982d377e22b10162d3e89fec07614ac9121d8b9cc7167d50226a26bc08cab78f1f993fa1da4f76202a3cf97d7fcccd5ae8596af7b017d899e9081ff767690187c8eae5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb5a4b2992d9632310473cacc05307c7c7e7ccd4972452e880c5b854afa956929aee5c7f58d5abacdc85e25b4ef02bed7f67309483fc23ac1d87f4539827e7714f03e42d4e7cca2af5d13618ceec9deb0145bf896736e82b86b8bbeaa3faa8afd83de4896fddaa328223b9d146e9c0dff81550c007df64376508b424e26cda66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b798e207cb1f19151146d3d3c2348830108a02d170ab3a20436b74d9bdeaafad15bd425985c7ab5007c9b874e41ff68fc6459cc36ff36ecc076c8ddc65de98b1d0d8fcc1aafe76d4e139bcc91b504415474d9a572e5e682ad0b54a621051eb3124ff9bee74cfd4148946b0247e26672bf396de62b1a57dcac532dbb455dd4ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6117561ebf1533d5e03e9c73448c76febf5d0bc6957a88634850ece73ca489e86a2330cca0a367e3927b5df12abe17194a6a302e963d86a3af20db8e27cbe6a21bbae78120a30edfe0d80e21339bd79ef34d852989378c9e09c3f9fa480611e87317826bcd5dbf980743fc7b5e1c3e5cf3a30853386a3b6f9f8209d7d4da9a3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9882d47d0e887299af3fd085e3daee1d0e7de57056bb16bf841588b5764fddf2b170a3a0381ff7c03dea083e1533237d1e37c894252a1100d89a332fbad696e1c406c9896eda11293112338557f365501b27838834d636910b6d6c294e403e147657b732fcbe2775906bf42cb5e3ef6be7ae3e79f17c33fc4da85c6c2f458e83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecfb8617f94899f17444fa923337a08774d20713c2f273fb56af95dc0620b6f6f3d3316005cc659eb2fc54a9e25fca8f65b8209c4258801d8c1c48a6f7f8b423e9c78a80e55b8e8b315f9e41ccce03a60fcdcec83c06f38f9857015280d29d5a19cc69930a7303c212be1632c3f8149aa473acde8613a41ab7e01c17780b85f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h513a18dbbd037f058fb2433c25a0a0623775f2a1ad38de9e37c4c1368bc71c936db2ea9cfb04954a54f2317da9c6308e68af17b5a6ab0fd4a8dcd21788f1fb831702dd1c2ac6cfdd5aefec4eca28dd8a2995979284fd81638122fabd0a220562898483fdf7d8d26902161912f7a5188be0aa084b1836a05f4a1c50565d8a7e21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fa6bbc0819e0f87ef7be1aa8d5645a7c93aed020a8170372076cc6f288e6f89acd5790b37ef13e3d002f63f2b0179f19fe0582685f26a23d29c1b04931d68abcb7cafb597edba9100fe235411b0a949f49db27827b5e206bff40ae52c6faaaeb44f5ea21091d7330605129ea10a3b9b1ed7f0539f9586a3fc94b4c6982e9814;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3a99371c4af1858e23c8dc6978021c541f84a2c9eb64f1646664d450b720fd18976c0892fa98592537fdf03666dc6b0cceab6ae9a6c9c0351dc2b1f133aa6a9952d9330c2e7a3cc1bc0a9fea43f27097f1868ecd49a20220ad1b5c7af5c929bee8724c1fcfa2b81a1e3fb7c29a4e64cd2c87bd25b9f952aeb55eab416a3eb3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79a4349f7b912a1125ffe23874675ab2d0645d5a5af54c46f9eab53ee9af47008d8da9cc79930d5a050638910535338248772f02d2ad22bea0cbe0302141553af850ec147d64d9904a50a0455fdda1491db91b566ceb1f8e933954224438cbaf1aca7cc99e60f43c62de92ba4cef4094ec466a63a3eea04ec164aca3bf3bc781;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0874689c3ab74e98deb36c295ae2b5d077c6d16415d4e386c7876b7d04bdd32a62cbf7e8faa8d8c1407183316c977df0d5abe1a5ce15808e997d5f085c3ca71852d5cc1d1b0638a8c921de12610b72edf306aec376b8a02ae72634673bf33ec1cbe350151b3a5b6e8b812d335f4c0f45f708d0654ed8eddef90f7f029653d0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e3c7022a9aac2c77338e6f08cedae2a9dfd4f7ca1f3a499b4fd3ca845391fa3e79a9001b0cb37513eabe88addea7904e31b774e064a5513884e0238b6a625765f817f16d354c54a7130f1c73079b0629e634ebf9c209fd61c3e0d6716f29656eabda894e107a237de031ce8460c428170de46bec5076b79b8b1628ee8a9421b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1e08e623cbd23119e2da2eba190962c1e0f988e258c27fbb31919c7472acf048d95c3313cef7b5ee61221341df60ce08833e534450d09235d8f46cd001afea8c3a130832dbc01b5a9e1d21b6126b1f54e79ca459096b6e2b9f20c907431dbf2925cc23b3efa1afd705245fcc37eb4de574858b396729dd39d82fe2e292eb8db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b91cc29300def24f66bdeee0138a1332230ae4e6643ecfdc4ca610dc73dbaa7dbd7f552b7e80509a01ded4a4fd4d41f9c1836fb458eaaa185366ee374218ba88fef70dfcbf5048a1f1c412d01c28a9eb6c58ea9f87852412e1ee77e0d5d5d6644359e8a601c9e7e0699d42d46d8bb2c6b8c63e213007fbc40e123e9cdfa7255;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57a15fbd6c145d85628f499b7ee66a0f844a737025cf24a8ea6ab3af8753b8073ba9579ece0574c9952b1fbbbb274a3d7f06036876764ddf5e6d50048fa5205692d24b0d3d44eae82d5b4006b1fb2fe2459a372170a6ac0304ea4d6ca949f8b6214be268f358446ca0ac39d23d044ccbf796d9a3e2d2cd9b5e1cbab757ab1f7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4882b5e8e925e64b0164ea405d5d04511fb46600f7b688a2ce8ab77ee47d6a2381ede70c8782f416dcb3dfb3080570f0c655915ab71572289b8c3d9db705b849ec2699fcfdf40e7e1b94ed2a5da2b79e67f54dbc5b132a01dae38c3e0c31f8c9e9be5933fe08cb41b5488fd02de4d0480ad509a3759fac530b97180a9e5bcb5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfdc079aaff9ab651ba304a3b30dc71cfea5165edda644162c97c17be7e3e11e5cb53e682b11cacb406f46a3c470bcf2879890d9badb78bff7733552785676d327b3f28e6632997a5c6e2f16b6497094810afc17a500bd2187d8e75ebec2e2f92c16a7ea3c5c8b30b94e44b3aa9ab5ecfa0c3ef8171fc7238b21cd35a3893987;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d17fde48a97a3fb83ad017d52b7539d78ea6dd0309a6e156a9181bc159a02e74fc08accd715f029badec650b1ba7f7655e7396931a35cf1fafe7c19b34e812864ad8b1a214e7a7d3074f43efdede0f1626e17fb3c7f39e7cea0efabb39a375eec71ffad703fd1cbc351829d79d9e2ccb1d57f612b124159f0c6d9689ac549e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cb3fbb3b624b81cafd471b8b2956e2ee2e14e90bae73c894a1c801c529aca6f3342a5210246d74e8fb028512c77693216b6a40c00099651eab085b3219353da0965c77379d0e6ac620b736df17a3b79841e791dbb4bcaf7551e0a8e82391d53f14ee378cbae495b82c79cdc63e67796c39fd203795ac418829c9789a9ff3a60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h210abadc726323a9da156601a56f242f941285e10e1e6aa02c1cd53c25f9b05553405e93cca8bccdea9a6f999e27928718f6db6b3070c7859079895e5f7116d8d70f3e19491ceedb651a1c54c0bd206e10d8a4b3bf88e936c5ffdf5bd7aeb9ab26b275d9b2bb51d4f9bc45159117325b8d2fe5033138135c4f86dc637320bf20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha592919f5bf0697bab6bcf5aedb993641808a1d5dcb085004271ed28fd2ffe16d1acd87df40414217caeb11b13ce9b08ecbf65b820a43bda1baff5a600c88c1aecb25ec7a15ba5cd5520065ac7b58e7a3253ddbf33cd1bff946e4fc31549790529d4d597b7ea245ffc44a136f19dc112f1dabcec4cd393a21c3a976be106a5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5536bb13fbd675866be6930eabcd47d65fc3876c2b01b70b40094d97ab464aea4480ab1207f948eb1763fb553b5c06bdb6dc8b519769485afb89d7245e1f8993a36dafb83f3c63538b015d92b5ff19bd155224f798c07ff72b44e23536d0d8c1f1c1b97e0a20be2227fb673082473685d11644e73ff8d697e99f0f3506d75be9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a0764610c315c4cdc6b8f046a7da1c8dadd3a116cf706b4f1717589b1c922b42648491b0ddc2fadb7d6e4e065e24ce548bf20657f79848eca57f9a29b6a285777c8877e2a89298e409167afed67fc25ae0e1f438cbc3b0c12487257adf2b9f5b4f8cbfe5b28167beb266e9b8c7156603a9370869c848e3c468a53705e2597c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6eb066f158e7f4b4930545dcd27fb196825af1b19a2dd2b89eae287dae8ee5c8c55fbfb75173c39c1178d5779cc9e5da2bd6474dfb06341ab0f0126012b22eb671b17fb921af3ac1809ad03ef5536bc1d7aafc83270c5a98d065916bc7611e45d7cf768ecc987b40e5e34284bf3249724698c672c030ad1b8db13e691e92955;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13be3a8118ccf34c1df7c3819a13f5fe15d527813fd6e6cd9fc693e9e1f96251a6706d813d17a44f540137a80b9e23e58d144df5d3ba48ad8b3623833c86e01c08480c19be0c09f2f1ada26d6cc6d62a22d878f0113d13069a21d232b9f5daf20a5355bb0f3b958f0a55df1a19035a72f8e9bbd2ade69397d1c61bb75162964a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h549a19cca3cb6ad554a33cbc2284244b14f145462ae661731d197217a395f9460348787b04324f5c4b09ca5026bcc78cd184c1bafd725bf64a8717ccdea063c9e5321d84707ce190f59b22b68bbb56329ce9c10631f7ae8beb91c1ad00cd39b22ba5197fe9495169a75cffab6510fa9eefb8c1223b3ed7e5f621194e013df75a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h530dc5a657d27a2d29d4ceb0d03eedf4071c196439a96586b7ae0f560b69bfec9d8f8e03fb2374bd7ec9faa9ce45ebcd061c3c8b8f691628b18c162dcf3859de7693b1694755ce3caada71ddd37cc6d4ffaf41aec3414f48953a6640112ae6208658d26a165f6b9b9fe216fbf522c01c66236341e39eefb23ccce0b548cbee35;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba8ed45c5a472d84b8d0f540e52c0cd79bf6f86cc72424056cb5458b2d6167ad83d5867f120895e786bcc351a82a88be5201c5668dcafa0b73c8279c32cd9e33133747f4cf382d66bd2fbb5dabad626737fa4ee522b0c526f53ef4eecd42fa5275b299bdace3e5fe4c8367ceb6cdd49d0464eebefbcde53dbac06d89479d0242;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc224207d23efad206cf0447a80a6f0bd1ee0267776178093deb0db7d7c45c39702de7a4b93cfe2f6b842a56458b641ec8959b3b53a16d45ee8564d09cc3e31e23dbaba19ebe79abf9cfcdf1238f0d60358085e08b7098cae8566db10a76bc366fac79aaf5189605acb6b800948a9808755aa50317e22b8166b83ce08727bca2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b037b113649cf22610188ed154ba707038498225e6f270562fa24ef36f15972c52b8d7cd8ea87dea34478857944a283cc92ba57b51034ba61b83544bf65196acc26889be1a993e2ff75369ba5c099e155d81d0ed2ec60f44ad854b7500c7501d1c49fd53ae91899ec0d97c5d3fdc59a6401863c54bbe209a7d8bce2083ed451;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7292b71ed286be154a3a156813d85c16298b33ebf2ff6d5a4ceb519d49cece16888c61feb556f174b1fefad2bc4bc68d05bddf44e4aa595482cb32f96ee92478b2600d997eae869499e90e8a171a43e2fa87e561858e0853a61e33bd9dda09c3b16affcdcd4a83ae5dd8fdfb96724bbe12c2c56f4c71081f066911643a3a07d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa887b2c39c94a0a738af3fad73c109e96d220c5a9e03775ea6f44926ed9bc162a5cb2ce4dfb8fe3fd35fe1be22b5f25a0d5e403279971229cba978c9ecfa148488e0a70510314936639c81f256fbe7e83da88816394bd2d172c4f9dae3ef146ddd5d07cad1920094c457ad39063b961fda2ec13571c8189b8b370af3c84ac95;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1c1eae3b914bee7420fb01bc84df9410b4951ab227f151b686c9d64491cfc61837eb77c38e846a5ebd5278ebf70223599a84048b78877fd7cab6fc2cdd00ac7b285c66ca3ecd00eccd68efbd3e3b2b3454ea307e0b97dc8af66f9c6787c3bba4f00d4904be65c505f72206f96a86fc1356c8af0fff7c64fbf9cef7d3a8b7903;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ffa3164f0db670bc2c25ec007ddae04ed63ffabac8e6f047d071d2b9b5b0f02b41f7cb66b3840c95fdaf543c09472a07cc31eece403e0cc667dfd5a2e7d63618b33d4d23e415c5d4836438b5ff7b8b832182b5ec4e157528cc1adc561eef0b12cd68d3602365e10ec56a54a11caf26cbeee5ada197fdde3c1e1c0da9770015a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedf3af1c73ee8cd229f25a32f68887d00ce0f90f9dfb69fefc3db6991231ac42edf04ef1c7325a3e9b5624476f9e53f456922d420486a446b26e82c9b9a88e0d12a5e7293f1115b33f37a7842c5a22e6a0e028db7718a500753c2a69fec725c10f0e86e365ff3013f3eee2c1e1494eaa66d2e45e67ab791c138cfb8b3dcca555;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23289babf8619c26cc44f6c0ebe30b1d6ff3c5ed82ea904c1ca86155c787b10effe60a680c14c77a413924135c344e71497ecedcb553b528fded8d517dd4353232ec82bde0abad3b5797ad3a0edb2d5abe3ca7c12d1fe5c16aa82de5575eb208965df4a99ad01cb46c2dfe43c440a4c7decdcb511d7cb2da348038de4946bb46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5280ecfd8ecd38b6103b6427878b359b28fa17b43bb5d0dbe2b00a41e1d46d39c32826bb37070de875b073e41c7cc8e9df552773e6e97d850d25e8ca04bb111e076632d20d70f24161f2efbe686a13d19943761bbc045a1b6c94814fe5c3c6cb3de9b40c21e9f3e32957a1b377286ac95d5f543911989efe8b725665ee6c21ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1a16064bba1bb09bbbb234c098eafc6034bd2d4c5e03a526230d6494291a6376d75245aa509a1cbb9cdb31f744086a4232d8c22bc21920a1f9a07cd45ce26357dc14f9fb4ffc248ad20697a6b13e4b41df28cc5776ed7f71ca2d04f8c80d88cf6ff0e6218f1a994790b534f3633bcbe48d9d456b625f798014388bbf732c368;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed894544aa32dc781a5fa50aa55671db6edddc5ae406237cd07d4f5e0207eebcabbf1ac04fcf9afb053912a2536811fb5cd2fdcbc138008c3015439d3089a344669a6611921a9fd7334ad041594a04c2d4be95cb6a4f3df88b0ff65473af74636aa7407aa44fca2fd01df655a432eb4f243be053708a6bbac33afa9d5b913123;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bfabff522499cfd872e82d9bbc52983cb18e51c653ed8dd3f286c70d4b5e1bc00800fe93e1d7387d9d24c153b541d21eb1c56afa80a76075731b7dc7221bcda5dec4137d2934aa1deff5c7b7dc1d176e7b9a587fe131d21d2af0c48ab055de8d1603274ce0ed38013e453b18a33ece6a474fcdd9e6cab9d5d0c8a4af5f15648;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5783f077dd63c388686f59016ea8710a7c9ccf0bac10cd6b4126bc879b5708197ecabe68a5826f7f6949e483cd2baaf14db9b6e77c3d96160cd9d616a4c3bb83c54f801f5b47a20fa0758c893d67061df5f688f77eca9aa99521bda15033edfcdd791f5c574bd42cb7d09c9a3bb328b35e864fea8ca1baa7e8849db5ea76f3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33997860b7b9a41aecb76ca4f83eac1ad3c14da73de0ceb2c9c24b59a184528c605d949230dd2625c80db2c43ea1ea209573dc8d1ece0359e794ddbc035f00cfdcf49fa9d5e14cd40673fba63f3e10f7c9c976414159f16cd200c06c8e4f89bfee8e3bdee45620362990af206baf3ba592828385f584f5fb73f82a96ca97b83c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h176871525b9dd11aa952a15060012ac53b4831d74b26edd3fcca7ae54fd0a72738eda719b942554d3d0226f78fc14cb17807acedda6781975835d94727b8e00dff01b833fee5eede392309c0091da8e1b37d427a60f6f2914ff7d4b194c759e5cb3412164156c55d7ff9c2ff4f17cc8153aa810272d108d0fb3b78ae062ba855;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he84b9459d7a4ab94b25e16d3f8b8e283c35b004f8a9bb4734582e4541aba352d0f69332431d21499fa594625bbdfebc18b0c7a86465b347846b795744940f97f805f85de7e40d3ce67a7c98663ca69c0de92f1dfb05d0a60c120ac2f67dfbe8654cad30995469f3a4e0462c0fe8b8ae6946bb0323735aec6b0b7956b34ad0abb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5f64b3a746b735e597b77a66c2eeabf28bd6d6a1f2366eb35bcc0a000400098af391f1744fedc374f1892dc974d40f29e2d150bf77e7e023baa3dcdfef0634c67d730d84ebc5b9274b26f805871fc19c8f40b8826b83a6a0963e20d0d7655f5e9934e344d2982f1bb5bc90f4113cf7e888505b6c8fe35614bae6e56b644b2e20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd53b860591a17c74057b54d321dad4c15c5b06184b27d5a5d25e34634703109799489921cc847f9ece91c5570eb0cd3052e559eea59d4305522e44b4b71cba6172a87d323ca44df635a1c27515a5196156f103eb1dd7a0e8b2e44950f6afa5149e8d6bd63c34a6cdba119eebdb70a99fb74e4f31266e8a73978e178d3be8f136;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61738a2ab63db417943924d8b61804e3b00bdddbf2215575201f16d5cfaa748d58675d767895165e824ec69dd3a9019e55cc3acc704f5272a55a8e31245ffffdb1bb705438a5ee27aec41b12a6c2c12266180b3bcbf9bc1670a5d828ea52f61993290b987ad888a3a3e433d5f4ee432d0c441abc1a58f998a782f0a41c6a1a62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h281617d81bf21c90bc3ddf6f50a5d72bc34ce9957e79e280671082d324d869c81e66a4c2611278766904725b01b97978911544bb5c22945b61d30fc73cabfa0ee6a59a60e48fc1a59cf61f0fcaddd0aa9ee2245c16defd3071c421c2a4a3c8542329fd30660e3f34c601559e8d301888b6950d529696e14a2a9b6f6809a174e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h845cd8a091c0e886eeb9ac19063ba153df69b000730eb281223b95673c31569cd8947810cc4c97a64f9c0bebc187e90d163fd24064319b82604657c5df6f5d42da95cedb3d47277232d854243019762d76c7a56d43ecb5192881804939c584a26c4efe923b3aab8f1475dc79da7180c30e0b93ae3373ea980dd9624f9a5f899a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56be27c07552f842f3acf3430dc2dc4ef15fc5e0bf5cb08be11b4409b3d19065ef0c99309453ca1196550e5ee9db2ffbf80da09cf0fbfbc239bb66ff8a1e2a3f1363682072be2c3a8800963da517ab6fb176c3d1762573d3d6650e50ab4704ccc45bc55097c1ae6ed304dac0548493d686009665df8fb3ab0a331c2515a4b578;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e0485b07dcd34ff2fa723f828ead7f74a49ce6ed2f614dfc0d2da6677258daf423bfd7595915cfc52eb8bf5a4c49f292a4a86ff7cbd86dd3d0938ef5f6e6522eae3bdaff7d049603e233bca8feb8455eb49c2eb54e1f5a9a303e9fea24c56d480b0bc487abef91366334bb270de0cacd064f37c02b627a097053d4f23f0b7cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habf9cc69bd00882c73fa8e431e79d0f55398a92e42875cea7cf9338035d1ca988a4add895b9aea57da9b6b01eb004e45e44f230a935a62d548f70f50f7d3cd604532ccef6c7008e68cfc4aaa48d3ac1504a543ff993e6885303f414809a0c9d6ec4a2db4abf1b42196bfa3dc971afa7c7f58620991d50c420842b24fdf84fe5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f16cb8bc9c49a37790d937e273c1dad2cef9ac4eb52fc6213f503c643be8ab46390ab75d3c8c7224f4c4c2d5889cdfae736505b65332b8c38c6be62198f3f0750cb298534803617a8b0832dd85a57919c8e3181e3172f0de3a5654a4417c213d17aaf7b70885b4c56cca0050fe70c2f74f4b37abd622fd732b22222abbf4ee6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fc0c23eabb2689de0c1d374a9641322fec1fdd959c571c65ce34644edcd919dacdcc5ceaa18137d85cbc99281e42aa05f9db58615430be9cc522ba1333bf8e52761739a5f23e3408d82809e0e5a9c087f16138ae47a5af588a133dac8a7055460865b8448608693d9b8aae698df7ecc055868dd36afd634f75d32f9e7df3e06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf04edfa3a3d3590eb597719d909298e32863bf470ac7de8d7a12b6000c6fe7b35188f9e8f898d7dd2129c66bf5c5372525080b9b46cd710af44783a68f491acf640b14cae8bf3fe1995ed7b41b0da393ba714f1ada3c5e3a4e19883ccb98b6d116722eeb0a95f35f33e5d76821d927353fd187b5086c62c2bb8e672b521389dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha38dc322916050272ffac010c6f59104092246e0c8e1079a7e559750f091a88c36e4ad223bc2abd30cd31f7b41256dd49e9c715393485f853351d4f083a771bf61b418e52e1dcb7416f5ce5358b9007c63c4f58d1a7378e744f57b05111d85292858fd0d95bdd55fc4641b305c3fe27d6cec84be9ddf1c21595835a590e102d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3a8725525d5e76520b2a77fa5bfb392eeb147cd1adb23fe2544a1a0fc2300cea9592dfda94142845971285b63abfbc3908459f292aae4d59137b9ffbff8823ca7f27269e7f020db3ddc03a8e48baff5f6375d4236cfaa2228e427caa12f87cefa636567d1c261d3ad62c4397e6160a5ea6ffbb04c05180b8db06a5b70ddf39e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d00f12b3a53010df4b7e1730c8aa8512eaaace82c9cc604872cc148806d18af294abb49da860527aaf2a06daa6a1f7accc73e4e0134ae4615f1f37c0f31b8d58619ce7b5814ffa74e80f0ffcb3c130522d96eab27a578e28e8515e6df1c0743a8b559ab3f001bb42dab991227346771a64eb161b96574dcd359312101a974a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf8e135b71cd641b1f3461d25133c618be3ab26c8de21d4ea952ffdf6c5e41f71fbad9c942e7cdb8fe71539a9e06ad4def99232f33b2cbc1e0d7376c04bb49b9623fbcccad405d118f17ebe661731b6d498ee9a4cb04f2e6e575186d7d15db96cc3b81aabe8b0f8e5d74b9529ca80481b5cff5ac2268b8f13f5ea7e1748aaff1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9dd866ebf0e6786d800148df47375b3b09c3258bfa3b9d53726c9f322eb8a1c495ae7e528602514de1330a6e07776bdd62ed8a966d7ff1da693f0ce6ef678ef4b425be214b0e0851cadba4ed5164c4f46344e308ceffec2a757402cccd2ecf3386b20e9c8a03ab788e585a5a1b6ce047013d5f5429d9591f1c441182f30a005;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bf4235045c5bd4b0fb39fca228f3328e83e60af7d74fd8901237864c2748a062200df9113e0d2e6d35f4cae42f48ba76f004a1aebc68b738f61ce6cefc08b1879a6ec0df7d504a053490d298c38043f19ed9c9c67ccdd98ea1d0d6e44e25ef195fe23e2aafb66e502267c409fc66a516178e9fb3217df8f239dc415920b6932;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e7547f59a6df18bedea66d4bb2ca06dca220111c4b477d0d5373a8c72ef0ee75d0e7c6b7c458fdd3f8df6621fa3f3476ee37f1307bdf68953c9369714a82e497117cb1ce2758664b76ead189b06a8f096be2a900ccb92804359d189f6dffd6abf2e7cc0ed2b45fe8527c76902d636bee9b0a97d48f0a8f48dbbd8cb10e6a680;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18fc0311ffc369fdab2174ca6a19d5b5ce98dfe333d8bf23c2d957dea4cd3ae9a1b1080ae9d49434780564aa187d45c4a481961b0690abd9a31f1ba47346368ba16ab330a01dd6179a67f5a49fc9ab45850add7ab569899642bd369ed7844a0b2e8f445a43ed929f43600ff80dd3bc9571e3f10a9cdc52b7077e389c7a1ee29d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61057280843822c2d311fc37a4f5c3a7af1e8b7e7f2f3518af448e4622ae46252477bc7ae7e8d625a0b0942653f317dd6f20e4af58dddebecbb540eac787a2892922f3bdde729f695d03bd3e7935367d8da7760d18dc2043fa6b80e8e7c6572e67cdbf1a123f6e5091a5de5c190eb6418c942d9400ae0a31b826ad6af0e06e2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7008b24ead7029b9b4df6a76dd0c1dbfeb322e3b4b871f07c3b1b9bfa8ad703574b94327decfef550a8829c50ccaf8798496c91ef3881e06be4daf87a635fec14f5aafbf3c69959b2f04be42be255c208ac0b899e5a7ac9b61cf91d67d55c215e1149160f943cd04086858bbdb244505ddfae81689bd50c74ede8370362dccc0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h437a71f49578e4fb360b9b26ee7addc249552e9fb20f4888dee80f3ebbfca0401c7684c99674ec1bfe50674fcb56b1f0e77885f3481d516dbeaf4eeb0920887e7f697239e1c902eceeefd715972292bce94c6596ad5b1d0edec2d77d1755dde26fb5b6ed1a967eb22aa61c7038bb725086044f8ef31cef50fae02c350e5ffe8a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32498877351360e34526a2b67039fafab267653232dc91bf9e5c37249e1a8e3070e1c58a998ab846fef3ad215bcb0574da5aa0ec503de5255e768c54e9cc19e01d342db0996d5f2d23cde6e88bfe64b613a84541e597ba5a28211fe2298094fbb70d0dec00465b6b6a4d084da5410417e70055cdcd697cb7be232d64cede59df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfeb2b70addc83257b703c497a2732c35284610398fcd27c086b82063b514ce8a52b86b0ab727f54bd86d46ae316175cb4bde265400f9d5b0c29de603a4c904d417d439a1c8a96781d72ea2de7f8171a3b75f212f462845c6d3a5d7a99f2d90525d72698629b47aadd107332f4329e722988d9f8741d58eb2521a06ae42ed0680;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4334ce673388965773c8769f87da4fbb6a6eb6b528b2b28a2d57c4f8e0ba7f6269dc56b74ba77e1c7dd349f6e985156f18b2e43f8d721ed23566d2a691098bc06974690b79de7f44a17e53250ed9e7fc90a5d7761c75d76e8985051f59ce7f3900f0ea3d0e2361038a0120272e87e26210c78c9277a2d103c49b109fd2740bd0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc58672ad8dbddaba1116fa2b7def8f0dc50b6234ae8c4e321d4b52709a5e3ce1ad9221df6b316c5c030ec70bede675ff0448c415ef3aa9c10c3bec5619cef130f209c9c298f2bac94fcd5416b015d2f13711578f71692da4bf860f9e530f4e6f57cfb35c212fa2896bebf3e6a683073eedaeb3708c52c215e7f88ca94f8f3688;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4aa4a359f2af409b44ae407d86cce9ca915467e9b1129b2013ea08e705023a55a0b46fbff8823be254c53487e196534acc0123814a7d3d6c51056a2cf29b208cb770ad02c74d3b1385a15b0b23f02fbbde2b87b38aab7895e90c050e2f821dcaf42fc38009f657ecef10370b98c186ef6fa7c166f1f8068424881078d0e91af1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h185163fadf1bcc8638dffba2e4bb0d64ebfd9d5c1cc417760622f8d98ab18b9239572682293e3d6b09df6d2760b01330b45eb1e39b1ca8c311a4bfcda96f09d166acc650ad1a259c57b9a2364ef98e3817a351a56de97445fb4b0e35144fc21c89ed995439c1e880b5b02690469f981d02a1f5cb6114bc43bf689e7abbcd4726;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca9c22fe73f94bb8b58bbee3e7ef0145d3e5bdc5cc0473298b6d5a6c51e0727998d38f4a810ddc8f8fca8c000cc61df0f66fabda39bdd95cab6d296c3999286538c165079741201f314e9d3f23f1c70a401e0363ccbc6ebf64bcb268584e58c81618226a63f3927aceabd76007051f2f343d34496d0f3e6cb63fd4456d59690c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50af4d077029c88635e7a047625b40c4d403fbe7b2e395b3da2d3a18bf1739194a412a6fba22afce2e6a7897928aff49d9e8aa8f18a81807e1760cb58269dbde15576afc4f8069e055fe6a62ba6cfa1950d33719afb87016e9595cbdca536dcdd118d158c39ed3a77853d3c94b3a02611c95386d79b2cce69b5b3f1ff6cf6a60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44247dfe0c00180f15463dd12f28b474ddaeca931920855c6f977795b022d2ad99b62897c0e36b97b5ed7ab0c33363ddc41093629f02a8360a45ac90afee96ea1256ae4e1b9d36db35ce4a5932c8968008b9bdcbaec67478a525eb4439209be41b9936f2d7d0a053f34789c14e626953860f1b209e1d1f1f32c81ebe79380b15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcaf6dc8329fcff1d9253f39d5eae4ecb1b18eda153b337c4c7bcf3dda7986efa0d325bb4ed1d9b96545b94d221d4a632a5f1c5aff727973d69250f91c00ce49cd4ac85ac0080f6601bfc2827a253ce236b9d10987fa1046b4a6294d4a5cd4d34ccd96ef7f05142e5a62ae70e4cfc7d598cdc1fb3a94fb98ae6ee1ee24bc458fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45dfbd7f52c7aa85249a38b0fc43c4c5848be0bbf515e4da1ee77b1f716fd0a69c5f38b764f4fab91192ca3b57b6283f437ef43e3f2128253468a760faf7bc420efa154c7501d6b7910117a7fdf8b2e03ae97a972dfb4884155062c1e9fb506821614bd36f5f9a9b45dfed834f9e2762795efea17b893e953de5d3ec1daeff35;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd575d546ab59179ce42c15f2b089719a8ffb66de842e39803b0c5a3e9309df3eae765d84c3da833e252b4c4123eaed41ef9cd82abd8f6f213369d26f2a347ae601cd255b295a7d751b1f9940f677fc5b722f35ea395c598bfa7ec2b2a25cc5432f60592a6df29faad3bf0d5209d431e4aef6db2be620e64de5810c54ecf380cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h849ae7084cff6c0c5fc52f9e52f0a2bbd46a1d4303b616a71a46edbb76ba635b22e73dbeabc19ab6a4b50218934b3129c7f91816ce03e178c0d8f431b355a4b95a57db3015f2638a628fc765b00c307d1411b31225efd691b42536de88081200c77fe178d6faeed3d339920367080e103dfed4042060e56fae962f951acc0964;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7da46ce752b9c0e6f3347627b8facb86f96796907e530ac45102dfbefae9f66b7673c34756490c95b4aab7240f0d7c2681741eff512f5b0f58673ed4e27a8dbca4e1201cd6c0cb84af4a1180cf33e6d737c6b73b77cfcd897d96458f9bfb739a015fff542673646b6dac88743311ba4b2d1703e3c2deb91881c2bf897066d20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9bc4e567860f7b08c4d234c4abca82ead55ea8e0832d7ea8cf493c0d04590994122d4c5a1af5f2d269a24a6cbbcde351a284ff879ad312e1a06a88d3678c84517ee26c24e1cbf2d68b8a74f7777a518951f389ff22d156927b4c189977a2fa1546f0e0393f65c21cdbaf55bd869c380a1a1b54782327ce9c7951726b7954fdd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1cfe84b2c6d5e5380c985402466dc883a787f4bd86edb07c43bc596885d59613a0e27bc1b8c680fee7b1628a12f8d8086aa4819305c4225e01661441f0a95694447f43e72cd97f5e9ea37d2504c5521c919ff741374e3c3c058ac8eb692b1426378e656a0fb3e2179415b3ceddf3ec25da696d393bfb730ea9634deae831abc6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd04dbe58c1c607925ad2b8edc60341edf0bbd4b6a7dfc8a32b92d2b0d503c3a97110b96fbc50d16a6ede303c4b0ed6bfacebd5e8f420968d85d76ec4bf889571c37d4e7b6422e5dcc07fbfb0f3feb41deab62d7da6f69515966200ded526466af427d6962e64961c64c1edb6fb6912e2d4ff66fcdb7ae73a7a60e36328b172c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbd1211276390b9dda4cb501b17b7359fc62bc22564898d0bd3d2627480b2955cd8baaadb69805af3322e3fe42d40b1a9df7acd9a6d461067830650b8b096060a867252434a77c4db87b56245db0277a6f98ccc1bb21927b4935d9ea432850720af190a92a36a40d3084eebcee78b2a0c7962c311ecb506da89afdb6a240da32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h217752054f6b60338bf5615fbbd8b6d3b9a59d3b4157dad7eb84f6da789e7f96fcc2c9961ff9ff35c05b2e513c7cd35e87a5f3af4d36aca1190d05e38bf81e344f5fdbd74b8b179b316d3a3790a6e235316ea1376e948784a54cfc590cbb1ac282670b6988bc423c1ac9b1c71e1b074f2277571b59ccd62812ab21cf6b87c02f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b9e782a943e685d53c9227719d4ecc96bc4f1e4398630593996066f866e220d7327c04afa40079ea5a5ad4b5e47fdb3b1208e5fddf1d0c65907070fe1c4684667271cb9a5e678533efa2a019b74fed25c8d93d6c6b605d812b27183cd19b875ee53dc66b33db5ab30251a0ec10533effe17a4db84859cb2cda54e0abc69140;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c57a321f4573d1f8d30a55f61f4721dc04912b2fbd0af90b782a707d3de9f5b38d220310b3f989c9bbe45f0ea70fecc011b1c8d70b63f0834c395675f95a1cbb07e108b23f3e8f294072c4740d9826997bec1fcdb0a587d70ee14f2eb0b244a0cd6c51e777e9f68936cb14cd478daa7341d6ff2517f01688ab31bd711d095b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fd246502bb99a532d232c8c083369f99b07fdea53dfccc185eb7d9d4d198e9de19884853b2a5a44688624776580a2c95634930ef2e53d54a8e8d200126af4618820890a63c3e0e2b493b439f4ccaa2dee163b654ec231853fa82c9a9f4a86a7761d2650ddaad537813e69f71c9e913cc72db627d61aeced1e6be1d079211fb7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7353784098df6e76f91c1a7a373b5cd6a3f4c5095c95e7277b12cdf2aa30d23da06a786f089cff74b3a83616eb8fdd962184b0932c0da2f158000a06a6df1700aa6d086095d0c852453aeed8b1c7e42e6521c816265f0c8f3877f45193e3747e58cfbcd0fa65c8a31d8491e5ef467fbbac0ce2653f1408651472b3502287da5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h960c3bea80640b648a8eaa46f070beea7ea5015991310f7e0c681635c9ea9a68bc950d663dfec9b0f4d3d36cc4e78fb85a3eb0de7484f7febbcd5ab9d8c8cd631993eb6fb138fcda6238f7f32036a1be224b1c24823229a482cd3629688113f5b6ecc0e787339cc3e8e3767de39b0558c0993bbd5b2129c07cb8026393a1fc0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17775d35ff829b136e849267c8368a36f2c30c7fbb4d5b2a0bd331e808d9e0d0b9916813ce44e2b68d55d27bf8eba8f89260297da6e7cd983e1ee91a62a2c79dbafcc544db2489103b004ea38979c3a210ef63a9d59f3ee568e9b2353f780f3477036e27fd36e150fda6e70140f711508c963c0fb7fd8c53e4544c46ad7481b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9edfe2515053f7bff033ce197caa48ca0660045d5567b0b7e15307897d6b05d99e07c7d02226f5c7ae8f1109cd1077e50db8f7da39c4e2c291da57eb851276f7eefa9c086a3d7af7371bb62eecf8e4bd3aa85c9484fd11d05746a4120d782c6a504a99be370400d41a859010d1760cd4641296b0d385659f6a07ddbafee7b870;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49ed103ef81184de920e085e77394e9b4126bf8fd1e5d62cbb9733c5fd45cd70ff2b92e5a7733347c6361a357410c1fd6bd2c1968329aeb68da9deaed943142ab6b0f0dfab87d9a011b0c3f4174cf3b43c90929663d7b2399ff69914bff27f2fa7ed9ddb7ebf71af6ec0c4f0ed4fc908393c9c48f8308839d2211dd2bc281f90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53542863d12ef79b3f73cfeea7132554c4f4648c4a4f5c1a91afaac8fb3b44d0b13aec116672de3410047c4efeee4abda7bdfaf5271f7f794fa5e9d368826264002001b86345f34e4bf96f0b99e65ef87e11f55d2dda883f4df72ef675270962cb90022e5b0d2642bcaaf168bdb255f8104473c598d09a5ae912adc03240e6a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90a03a635d2bf4d4693b976e6e88757c655cc6d10269ca511bc4be2023733d41bedc178f05613632ce83b2d9e3b7681c8f5c12252929bf38bb269e1c4c1463e04ebb94758a738c54fb20e04dd85e4523b43d6a5c66be60005726cb7f6977860edd64b25f25b47542e94f883a1bb77c9a4f6e30382da3f836a192b6a9263c356c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h363f90dc1e77f44631406d1bece943c333c34f0dec00a49473c466d65c4cd5b9c5f024f4ad7c58fbc62edfd44b804e546c5eada6c43ad93a906002a7f42b264862c921f9cc4c33b51d171d2c42e4429ef6bede256222fd1fd8d6552020ac026f96ef7532aebf116c14ef6f9b1c074b2c6ac065493adb5f4f4ea1c2bd04f0b95d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc3a8605ab63ebf95a071856c152b53d41e939057fcedfa91e7c0e0b34d84569306c7b8985abd51e32941878fe9725ef1fbae2af322d22541ccfc3d9701984e8b9258cb0003da6ea0afaa339a238566ce983d884844d33e0c55b4653f5d1d69803aa4a42db969bf9e7a0fe5ba7d5a033f6a865c0f33e258ffc9f9469ec14c041;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc1be0574111ee634f349624198e953ab83d65eb67add59a72a64d6dbfbb37efb60bdc847eaaeeddf5f01eceb4a65e1253d45030da34b6919767134ab9c2633e4f27e090e9c778a29286de6a6ac6108bc46307433b40c1d9ccdb0588e51306885184c6cf59fce38e1b93bbb0fa4844017989a1eff6c8c44f2beb94cea29546ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he615fa04ec3dd0c6b7146278a28eb705e30b7115900c9ba6c30dc9a8b4a9565155249d90e9194391aa6fb6ba16482b8b143ca7814c844f9f9b94a57be687e1979fbf105b37c949bf2243bdb7181f61cf3d780196c0ea2e517e010fc74fb1df3db443fcc4faa3b47a98d8562ce18bf55dc140849273ee1648001da8936fdb6cac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2afb90b7b7c375765dca2e4e8380173ceae71b29abba2ed146b028d01a6bbe003d80a34ad6de1476c7728ffb1685029a2d75ef37274823287c87d41e4ac2c82765e0bfb8dbe914da44c5a546966f0c812ec069017c2a4166340c054a50a4b18d7ba711343bb920477c83259d08c1c426f45c6add5a792aa544919e4b11f1373e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6071e7903b65fc5946bf2018b8819b0b0dd280eb4d0fb1565bc4c1be676d76f1099af9ef24bcedb99d5a6ae00eed158da2f031a10ed4d8a56b2c8c99c02d82effe6f0ac20214011a9a70ba41cdcaea703ddfef1b5c2a5a6b415051a044b4179a5a3da21d6688799e1f98ae92d47c18d082518842bafa7b0f429990210b7b928d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46ae39f2bbf5385d511ff3456cff17e4185600d54170c8d93eb0ac431653f9beada44cad2fd0bda09a31556f6b8802a903bf0a963965849b5e7253640e0dc53814ee6f7502dd26bae47c22248526099cb531ec7cd6c1d22a118fd2f0a9681a77d13962e6b66f45616ccbb340b2eaec68ef5bee3c605cb81773d4b164bde63748;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heccc1ebbedd7c64bc9ec6bd9d3e48bb285546c5e7e26519448b76554f0abaa33e3816171bad81f7e12f0f7e0b2d5b1fe07d4719bf448a9156c91a6e5cecbdb36d2d7ec0651d3732b69d071592f1403eba12128dda181543f91d7dd665767fe474403afc41593ada911811573799a499082925f6782564af6804c4a031824836;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc83fd7455a75bcaf94d7e67d7d7d67603575699445fa1ea8271a0a7ba98e3a072a8ccfb20fc873312873b82c0511a57e35cd1226fc08993e7567d4bb68d89aae0e40c9045dcf7d9ebd7d48abedd73b779c5acc07654c166f4d9a8b85bbb9d7500a457d15b9ab34cc8b98ce227ecc7b9f161b0da710cdae7de196a5e09f485b27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9c8d453ef7061bedfde40a0f0c15b0469674be98736a4cde504ca6fc1d2b725d868a6388a12a41d28eee1e711450170ddc497eb2a8a5d8cb7ab6786552dcc8bae31b2e1d473d5526e095e9ee8dee798808d1d0d349d43b2469b83f8b254418ac9ffa19b5d05e6091685f0efe14cb00c6654abe72224d1f403e96b0891c3b486;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc561f8f1737c25c3f3e38068293770f1d33223b649489db540e05e1fc263b7b5359cc196fe5eb62464319013f9c375585e0c9290bab702cc8d23dd8baf4a83c2635346ade9c48a1737a8bf2c55149f0642dc00f08a82331427249eec23f8e07c8a97d5f9711d4cce582b71afa3b2a53d5bc2eb9654e5aa6a5d2851c2b39237c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb84a062fb22293271f85e86b27c7d428c80e51161ec3438165e88347b23452f78a8ec27760737cfa63ac2cfcce92280f5e57a6bf7ea4f3216bf3ae0aab6e284360ab1f5bd2f5996710fae0ac51282c66b6bd931f04e890473dc27686daabd5eb2db3444f09db0d36e043d3053a8ccf1c8505faadd875db2a45d25872679643b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b492eefa7b4f9458538fa49184f3f2ddbedf3b83cd77f97109ea7ed2c699bf4b992fa57ad59a24aba10098d515bf63c057a3e22aaa7d84d08da4d5c12ab924e2313784c62048cf57f202252a6dc49ccb81654996df751043743411192ea73eea2cac9cb9e72c32680fc3d7844da66f4a73b555049fadff47ddab121238a7891;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff4df3e6ee84d194db96b6f9546fb0460e8fbd309f34d8d2ef12450718573bde47f96c240ed16d9c98a7fd9b52b9eb2df3a4405c498f71b8a2ecf781c1ebf6c152c25cd5ccb7f6c30b6c909d0c4905664921bcae85c219025ae5e789087807c7dcd7d9c77b671b882d7963274404488765f87809c261bba2d0de468d8814e583;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb43a91311a799244f95eff25f6efd8283d06c8a7fdf229fedb5759db41d39f1748f0d48c630abf8cd96823a4231c74b55a378d19cfa3919452dd6cd39ba6f38c667e8de54dfb0fd9f2f02012f0d753852ecd2650b0b97424a2b4374821c8c93072132774460d045bcf6f557930a747f5fad0b3ef14c76eacb0ad6d98c1ca42d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5143eda488600354f0d0258993ef9a4b8d3950f2f53c14ce96347e22870057ee4fcf3f4753920f27c89ce0f8f9abdaffb883ab82da5c16c95d510de1c6ba97f5b4f291b9acf38e49e9c920ed1580998596a577b10fea908cdd44b562b5dcc62dc3b587729ffb9118e0cc7683c0bfeaca94a02684613b477453cfe4f873c7502d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1aaefd3720cd0039dfb9041930a394898f00634978182d1171dcc31dd9ed2ae9d87b1bd743799924a3714ac26d05326996a3a859c3974fdf0b39af55b961019e3ec89e32eed8be1b4b6c78ed56bcc4d256baf5fb6140b6186fd05fff84127f0f94519f10aa604f5271cea32ddf0a172164009301f894bceb4dbedd2d846a2fc0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he77875c89c988f7f773d188e9cc74a8154f90c22c116b59596f81869d470906177b3b0f8cbca210e8e91bf6e9f52207a276acc59358ef3b8b598add43fee4ef606872458353160663a75cd6e94e62b1b794ad0b4bbf5e19b72fe2255b30503cb6e27b5ab79bb73311e38d03e48f68cb9da29a87bcd15caf783a5f963e0269e78;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bc646425bb1c71a11562d9f459ddf0f54f6e087625e160fafccedf5f25930829d89f1da221387d23ac4193a399f54722b16ebb26521b43dc11c54662362f291457c7d49b6d74bc334bce2260be2846732248201cdfe002ec31d1b9d631b06f656b46e57a259ddf8b9b923708cb91dc82accd07998dd491a9a173afa8337b978;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h557c53dfd548790033ed52ac61fc2b001e9ac863111523b26a126a09400e0da6e6e3b9f29cd24919ea56ee14c2b009f9a648c7b7bf061a80e9031c5a2a6daf6c33692a74065458b04b55c265872e2d38062d89159229b21c14e369ada65559c937f8b55e8061915eafb7d79b21419ecc9db1d5025422c359ac6907dc7c002e73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc0fcbed1e9d1fe802fe9e3ddb42cf991611f7a39ffa2a3c370cb735a441802f82344c028faf65f9accd53d253960ec6be0f583f300433487429cf6a3393e528534523e57dd99ea3a845be21a24c199503bc0e331d22e884d324d977c5be7c0ca5fe3b46e358e5dafe9f51c9917b77eb772de4d96b5d8ac362a99a792f848c35;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7718876b76c3a4302ad00b12b96e8ef42eb0619475654f951852d28dfb735df452e7ffa945c27d93c0de20dfe1c805dfdbbad6c666f6fa67643d6d7d1f148fb588938e0db0aac145499c96ead9cde4c2b09bea185690db87031322c12b5aecbb8ab2128c5b7520a3228af688dbf61f3a113264e80b5c8913d92f0312a7e6da0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5308ca9c1c1d1dc743e3832db7f47e5b30dd5fec2a0cd838d1aa15d8754bbec93016a158e794ae4bfc7e8da98dee49cf00fc0284f260f9043fbf5c77419fe6c7fb87037354634038be69d1b97e021d37ffcb62ddc78775c01b51b1dbb58cc139b5012030aee0b3835b0d4ffd9f408128e283343245de523eb0b7e352eeb4833c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7bec82b7ddce0e0e124b1d584af2e789073ad32f0deca50dd006a8fb8f5d339ebbd9f64ea3ecb22a2d388c9fb22406e697ca853e9a430a0476be3ae46eb4cd753aaee020856f9eef000f2078d5815b88f8427fda5d7b17f778b40207c888bf78d4d8445e83a8291b00c3cdf26ae92f698ed066ff15e408ecec4d34f974b03a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3402bec7cf95108350b9bd6e13bec944340689bf59a6f7b3c1b674c523e40fb809a66691c390786752b63adc94b28821fde2cb4c0cb0d0db2a4b9b231b51513196c823c9a2cd2e441435526292aa960ed0e6502bc2af93faebdc33907b73871e8758091b83bfee753bc24d2478d57bbd4a883c32995ae6c0c8a791365f9f7363;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8184833ebb7ce59c3980bbfc6ad004a1d3356a2b642221b5dd9b62b972a0adfb3256561994d0be9879acf9006a2f6c94d3400258640aa2411ab23dddf6d93022ba97242e5d13385ac87610b1ba746058b786520351c781d7ba0865c7e40ea48ae51a5ae0e0700a536f9d8c9c97076de4d030b5cfee1dbe2bc6c5212530f858c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23ab6875f68347b3dc837cf1b3695ad3ae381335eb2ccdab52eeb8511aefe034fee82729d4c3457d178e60c200039de0169b9ea6a7e3f3ea8e68c6fd3e74ea125e114baf5ed3de43e79c0caf5626230aeb06be9abdb1d1c9aa554b212ad248cf92b8df2e1cf14e077a13b6bc02c70f7a86826d72f39ba4201df8d7e4004fd31d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fe57470528e1b60f449994222dbe864212ee5b3eff529608a88e39dd4df8e840b3a2be6ddc17e783d172ca2530f05390a05ec45fa5783825a945122d0359199afd4d1230dc514b62d3ca23c76eb47173b22367782181fddd56cbd28f5ee80be8a392f633444f420baea1384fd874c198f69dc3e81b92d69d4d3f7925b01d06a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28edde273d6e7fb8a66f16ed2bb836cd9c36b179725559410d4e93790fd3fca4e2dc5b3f6d77a1d4f44ed655bd944e627f9c4bca9f42025d48e9b3076085f32a22a8a1f2e8a8f5884c8d6189f33acbe204dea8a9ea0c7ae2352ed22cae229944d19d38a4920c563ee437e970817efc931a70c586c6776bab32e669fb7c4b2c44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h876f5591a54c9d5773daa3b5735ce6b0b882c72994ae459d2ff49e2c7ab50cf79edb6d4f4d040c7aed01847eccfe8710316a29f5e697ddebb23fb6d6cea08d9b8fee2da356a4e4fffb48cde89ee3edf256d55d9bae1cb25352ef035f10d146314351c74048b24ab8c14bd85334422f9f2abaa06ad7aac396c2428dc3518933ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc16f09e40a8ab2e74e77d4bb55bf7a8207f3f94654e3ce4e239c06276666d5732f74a1411f6aebe473165403d04283b65ceec5b9e756d1bb276ca4e13c45cf585ee002e34cd76e36898941adef8ebe17b97ec18b2fbec5cbcb3de76bf9efd2719c3ee3fa3d655095f742e9c2910de9465babd64c6873a6605035b83947ca3ee1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62f5e4a41174acfd054773bd1a2f237305e19f667f30d6ede96f60c3bbab58435bab5880679233f2d09f7784a3fb8ac3ef06a2cc68702879cdf65b81d4809569a4fa4020b37c06ffc6fa63fa7e4dd8a54db503cbcdaaaa53e66c0b69ac9cd4ccfc826089d4a3dc196c3ba4b96df86f3fa2be1aa879d87ff1b3042ec72432ee70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ba85c029ceca44737c938b4917b3a12e1d4b5b7adaa6239f8aabffb7731f580f4c56945acda87951200c52683ea63f981db8b104b4698e283ce6ab56bbbc85e800930fd3950ea04758fcbe4262f28b447996a9dc9a7787b91167d3e8957eef317997076df0e447fbf7dac346455b2bc6c32b06adf981b44a6f287354bef67aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d5bdb66fcce73e1e6958f314c22cf65ce03e82cb77824ba4031e6ac5dc7ad456007d96c45fc145443422c11574b47cc256f604c3408e5279aebed5f6a3163b0cdefce006ca2f8a831d38ea85f70aff64ad3e6a5a29aee291581f4c27507db90f56c676ba4c8efffa43e84ac21f6fd9c0a40daf57723f0c8270dd5947efe524c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0813aaed1d5d70392defe9efae919aa9298f5c5c349f8c09152f69052a06a72f2a2bb3d9e5973d09dff51edc4992ebf55821cd8273831cb551e1cf4ceb473390d5a67366c0e9677a8102fb7650e26d780051b92d68e46771167134a7bd07ced5aa0fb1fd9dbd8c90c212c8da3d7d69995cd53fbea9436055458cabb4c21921f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38c00b0df44f82c688db3d2ca700a1ec69b573549cccfe7b150823182e37e14b06c25f2a08ef8159fc806b1e49c893993be9ed3204e53eab4766d5246a80f03ee248edd3a0f5eec158a6b1242971eb2222c6d0b51c5fc8a31cc29cbd48bc1310c28e704c571af69a63a01bf9a3754a303c796cf71e91e9cf0a8037bac7cc75a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58a3245d051ccb540efc22c7139bdf4f3c8b683d92baa0f1ab6e8f1bd744001ee374f5f1746bcf280302973b1e5e9c50fe167d910717719a43addff9aff6d5f22ff732a871672bb1eea442e802dd33600cf6427750de9be64276c19423158c220c5131b613e7f2a66e5c612b2460c05a3d790c28b57f796dcb4bed426160f0e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4a8ae3e14de8801a9668d9c36fb74b4a7650920d1956b86e6111a56a2dbe3b7055c78a573594ee97d5b93707b1dc74d27e81a2117276574fc395e64399f8a35672cef0affe895ae1f4771705d9816f8ad1e0483fdfe58e64b7434467d558500475cf67298678a2a9d8904525e35cc0dee97ac20cd485473c4568a65215a945ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb7d602f48b4905f75b34055377c1d3594cf5e803c8eedb12b350e1600abfb3262709c23551df5777cf2d3a23d5b736a0c868a2958d6f9116bacf967aa945c5f3a520e878817d1325aef58605a0821d16ae9a1310f3d46fbeeb968e23114785cd2bfa5f2edff957f92b31958bd86230bc5f647f7c235738b628bcca765496f62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd7dc3279780faf386c4e7be2fc12e0eb684adf1ed8df6e18fa02fca1fb82c47d0a59e0622fb579afa5ff28718f560272d8e51b1a2c09b61f8faa2e52d43fa1eacb0c3f978bb5fe32b7110d6178531cefde63147065faa9c721a76425e98ec7f096ec63c439ac0af5f6741f807e0341c70e1d7ce6564a2828ca2017ea20e0114;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha23b64429e9bc7aa93d2aa8976b28d799e601ae8bd2b4c405cfeb63116a7e5b52a14a7155a009e0ff2e8c57f01218693ece49ce932fa1b4ecebd4d45d01e539e6a26755ba73679e0ca6621bc3a1945a455555d0ff0db16ceffd7abdf6419518341ca25a2d6b59aa0f43cc9ff289e7cbca835aa72c0105e831f113a2a969ce685;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habcf9dd430b6be1b8926dfbc33ccadd7dbd8e0883276b85c5ee8f7d8f526f5dabd4cb155b0a85d6ca287c72c2682ec5c3948322a84c64770a754fb9025c52622408f747c779245ec772c6e056846799dffe41c8e1c1ea57abab422e1596105860db07d1b9a6dacb7f8c9f39a1c21acb44939dba2a028fafec4495eb70b774593;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e36925b2f794b07ccb71dfe28bec42e964368c30acae2ed735e342a37ae7ef084aacc317c4fd4422415d676c6b09f26eae945a07bfdc74de52633f1715c20f6cf38d590b35be1e5e0f13c71154a4af2ebc06032343c1c2263d4565d1fa3578ea68e16c81879ba991a8f94e4dfd37ae253d26b36b163450d05529dd5227ee452;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he760790f032e1bb3ac6e983bf04f443b4f8ba5f24e7ecfd12d6117b674e79c196e25471c71fccb0fba42e5f81f1fd5d0ba23901c0d910aeae743412395022ed22625b0c64eca580b1035421730fd0cbfb559954a3407d5de170befbdc2c8e96b4f6ff3fe536f589413e5d3d0e6a2750a2a1186c4fcc5e6b6d60bcf5a27d25d73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfab944fa10417be9a9b2b4bfe76ea4632ade88458a566f09f4d55c6904976adbe221fe1725ea27df1940ce2751481048865d580c6f6d98596f40ea49a35372c32f2a29e77f39543ef2a815fc399a9c239ff2ad2af564affdb411ca921fb2db12f467fbf6bb6ab64746a55d59c29530bddd515c5d62e1936e62f2a67b4722938f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85df935c9770bad76e0bfff0df93a80e79f66e5353c8e6d7acea403dd0b535331120892e7e68cf2dcfb7f1827cf20e52ac7bc829580b173bac117aab22d03e452794cc19e5ec6a6400fd1560ce71d45704b3e9f7352eb5c43b7e389f25f2fe768bcb26ccedfe30c17165928a52870d4674941dd348fa96f8073badbb02afffcc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7574e00f2de211ff69d4db3625eb14582f95cf54a22dcd8f2ec615977bc99811281409026a84bdf822a254a45924fa01dffc250729ee61c45ae9141c5d5fe85a4ccff9a36b4249df38307436bfe404f4fe1dd530971b1834ce7b3f2ba1b762b1ea1998a68052c030109fe6522ef9c2281fa6d3e42f76272921fb663b3631a2f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc470a5c46669e0d4fa944be0e05295003be348a797f3c1fa5ed757476a8b0e7dc4744fae34af5ceff23c83940eb1701acc377795058c6ab4b694c2bc77286d89f2b8f9cadbd967f8a0016960aea8a1960d71ed1ba48247046298b71cc5d1b7206c4166201e77d47be5430a565ab0e918d128d0cd3377b507c4bb018290bc1a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c8a2afb616f72b5214e236dace9fe3570d1597ee3d1979c9f0c980ebe8280a31d8b23fae048fdc1b0cb719ab0bda95665107458afa65fe107c25c2286bd3be3e90e35db76432838c3717c337f34961a4046fec61bc658a306aca311936e6624e4254889f3579a887b2d5d66271ed9d94e2076bd7ce85932ae1f6232d9a6205f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a6dcd0f088b84127787a9d1248af769a961e67f5744041faad7a9319776d780fff3af6572a17fedd0c3f1ce36a80394cf3dcc1f586257d3db3388c8259d87eb47d51ae46615aadb6c52431fd690b6c7631746367caebd82bfcad84dc6e87c291529e562515949a834dd05e0927292a56747e00246a87ca3faac5f8ecd38992a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcf0fe785f4e7bc49d294022f6d901cbaba32d0e67f4dcee42f24e06803e2930743dd1d78522a3d49dac75256173e411c1b1fcf99ab233b1f448952dc5b4278b76998a62071686b328e1b9259e2314e02a499b3b8cd5b7a7b2b532e41c35f959125e1dd6bb0c94f36c19e51bcce44198611e1ab274a5cc4700da02f5b8f9e47c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5b9e3c0675c484ffaf6d237e5a3349ba7116aa60fa0cd905874d75caabb6fea07c7bad61d3ed9a762b5081ea79854b57073e7c36e8703c6840a4bd40e0f6970874281daeaddc3d5d011a61a22ee1010b11ca30b48b1067ac3e85649cabede7a9f1378c922b447fe0196ffe753f24bf2b445e05ea7517d0c0a10f2b9c8dafcdc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1f209b5b3f29383d7f2deee553dac2d5094f1477f9906a67e6571a251e0652c90a21a2a7cd302eeb7fe26d4500cdde26b26f0d2a59406500e032f99dbca0c89a7be0121e2f031e84018bbe651d5fef8adac5c8fae47efc74b9f3e753874f81ae86639dfc9be4824b9af474d3222b6b1fedbab09f0d61a1871a3c322820142e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc961e6121a3524b82d2efc8c48b067c930ee86e76af6246aaa7459016140b44fb40c63c741b0b5e6aba569af2a3bb67b623e241301d2147b746925633a9872cb3bef568fee7c9472bbd3dec1396f27c1f4d476a3c1c316c30c1e83778c11c6f54bec6ed00e5a7e4db4bbf36a86d148eb59051a623c5a9bda0b8deef8a4b22c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b6dac35c903f537cc0bf6df9d4501ae8fb4838ba5132945a78775a5805e8b72a95e15a2d2aa326ad59a486c18184075b1c008dbe745058069f2e712a75311e29870d1956e0223b2fa1669fa4a4a3a8ecb068eb2f2b04c6571df29f0a7f153699eeb5655c6d2f76971673539e4634d3deb32fe2b9bd650fbd487498bae5a3e91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf75eff1c888f8df4a0180150707e3e131ce4fae5dc6d7c39f677a901b8ef909ccfe04f0b8583ec79eeff5f6f303d6126800ff8ac19667edfd129b10fa33fe52de2e9213389cc64e7783e9904f1e50bb0a5fcba17c60bb85068d3631f5cab79bf4a985b0b185b61152b7a97d9779588b4be58c263b782659db6c38de048bc4e9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d45cf4f1c428b71c3a10d7a855827c7897255abf146de079accff89a93518677ce474f9761d96da941305a91a4a259784d47cdcc8ad3fd0b3d3c0bd8d55bfa6ae5a8aa57e41823ace1d46ae216307a525319d8ec708ac5029c9f38e35a6fa21ef26f4dd83b2ec7f1dc8702385fe1756c2c700f8e7fa373d9e13acb926a7ddd9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h213822140134ce9e75c40e8e66505c535d10ea47d82174420bbfefc7a2f736a3de63c61869b4d56e28bbb0aa89a70f017f9b9aafdb88b4104b3cd13b3e47f6258bb8f43d45d7f8ce79fca5094b8a64033d9f70fef2be183da3c1de020629bf81ac15b20ce058540dc660b64ec3ab3845487df77e5c86a8a7fcd228ecc1d9d390;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b655b10d048dfbdd354bd20209f71676eb8cc99675c1c5a82d2d5c8c15798c3afa07d661e5780659176362a0a3977ef5468a4f89223295d064fa19b7e576ef61b7bd7efee784c4755dc5e67a83dd8e3db85151e0a2b2f725b5494c13e16b219f98d3fdbaebcd617c40702ac40f79caac202ceedd153f611f684a8e9fdb39f54;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4077c429f003a3fdd041c9b7144b9258ec4a8f5332383c7a11ca3f05f2f64e23736d4a86b4b379444ead15611d398bcd8d1228cd87b004a24c97c9970fb9aac017bc6a69e0e3b53e51705a0a00d4f7c8e89dd94c686d6de8335344204ef5773034dc0b369c71bf6d34123c77eb53387a4e72e81329fe3fbd584b7ceaab5289cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24ef89efe612c50ab3a65ba92cc620de32ac92198381f53fa8c14fbdb24da145a2d5782eb68440439ede25625f8e1288950a2d8740fa7803004b332212b74c1d36dcf69941ee2784f7435eb9399fdbfbab6be825a8d8454831d6c6eb9e21ec17d7cdc39a023da6b40a5453fd587b08a0488bd0bfe8a410d400679fde44844a87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9aa52818ccc0e000d6d723f27bf7e590cca3ba411afd5808124830c43d7e7db6927a35e4a733e3573e825411bb1c1dda82a032976670a6f5e861cdcfb95f8e2d9efe275ffe6c75889606dfae56e68973a38fc305d9f3ed796972471ad9f6abb1a22262b7d64f2d94246ea5799fa10ee331ceae51fe601f81bd041962f1852d54;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbdf6ade523601d23f8325647b0e32e8948a8a7ec4400001b4900f83b26a9763f80a2844fce8544a752bb928193577ea352ad5117ce7c6d4da11bcc1110fe77868f70557b6abaf1e376b9c65eb54174d65cfcadcc5375f81dfc5e0e3cbc6ec99ab72ac8b6792c0b86dc9678ace6de0d421e1eaa2442c3e41119c12034896ee79;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h230f0933e24ce672ebb966457a2627475fa926055cab21189722825913f527f83600ede822d8b7387c8c46eea936190ee2f0c1f5f4ac75673408a3e2abb35a658860fec6dbba34841adb08881392dddfbad6a163d6cdcb3f8b9b9b1baa0d8d116bfe5bf223ebadcda4b5e56e14933adc08fff5dc5a09fb9ea0e166f0fd5e165;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f983154399048c57603c1e931f1e736afc7469200ad40f3cdb6d08f75dc91dce97d48a85b9ea58bd336dba2828b2447df4754d4d35c04c257af1d216f91350881b731b19234c384e4fd68132f010c4b533dd0a6f56dab557f278e6bb97decb59c7f51480fb82ef2207cda6e5fbcbc63aaf475813c0ed95efdc45b5deb634054;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab64e6999f7a2bb97e1f9433a137a128d68912ed52fce76d5b900aed5e03a0ebbdf16a2e4cdadda3e4b7ad4fcf26d1cfe9b89e0a2ff9ce11443bf6a2549610fa115100cfed9fa9d43fbb949cf1487af6f24c0f772615b0d00c97fb14af0091a87f3cba924645423cfe3b7c8b62c5fc2c6be14e793b5d357ea8a31ca3f63a9693;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd89ffe636358d3c6b628dc7e6f0a39c6818bab039a0ce0bd7cb96cdc533239a08a943372b2ecdacc2743626ec2d918d1c0ebb7dd52ec8ba16b735f91b2764b6d17f3acdbd3d5a68f1a2f9b7d9b5b93d25d830b09b789d952d840af265edd0815ee0fc05f78d935949aac7bb9ec6bfb690ab7eb9ce00f3a50c0c3b5a46d57820;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6eeb6141d543ad8d523218b982a63b1e9a54dfe74c5435cb41bb02c8f5654089031c2e3acc66f29075f491b3c614d5a080a56fef19ab13fd9ab394471e2a76f183d1188a1cc8ebf0a13aff6d96144f86548e8f574fb5a5aca32200512f6382b86b290fa7b5f583fb45cf44f85094720ad699973e5f14347a7f899b630d54c28;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bced0c023e7cd57d20caa9069e4b92f99d0728730339a80256700f1cb838033f4106cbd1ba64c9bb6d4c882478bb141b3ee2044b64204a4211b6bb20b8f870313640393b38d34edcf72c399d7e6948089d0f73d7878a072a1d57e9ae17c2b2169e48a7963b77b6cde8db120e7d5a8cfa957729a04db6024049a93e84d207316;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6ea04efbf2c56ad01ce21222161731ea3ef0976c318f8ad6953b1402bb8a5076be963649e9a445d1ea70112c3e4d400d3c2921750114d10f73286be1f83237032ad234b5f902f65fa0cd316c947616d939780c87f07b64c794e51aab5f0512aa44f2e0e307916ff7e82d7816ea59b2bdd3f629f82cc77ee76210208e212ef66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94fe3565a7ecc586a44fa9cb2f1d4c228a94c7cce24a84346ac79414f8b29de515b676c912b052004f88422a55d823222687973289915afb951a170665a6a45610629817590fed51b1af197205cca37dbc6ea55147aade28fb5a9a81b13db620787febe62cdb5a81e994aab50771f3e8aa85f8898ddd9f115700108778724590;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he91de236741e139fdadec95aa4b2ab035ff792016545632bc05893c611700f8b8b303f3b837b8e8077b635f52ec060a2278a7163ef07cded84ee0f5b1f28564004bec51e130bcabc7926d0bea4c2da79bd806ea4245628da2df494a455899435dff19a674b2667ddf0ab6290572a4f130bc490e790ce47eaf21654ed3359c263;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7748eb1cde3c65eb84e3641aa8e35c19ed08f77d82e60618ef8d711250e9234baae768ed6f856ca5ba9da37c2056c1de10680440a7ba046466fade66be64645c3c736990c47ca41cf10487e2527eb85706b81a596115b3b2a22d0ceac99a3bdde368b501493cd1fd8cf5f94226200098c981f609818c1016292f679778f8e92a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h576ef24b31208e988e71a4b55695f922321c945b6c203b4b4bc02c4dd3f6f89f4486f647f85fa9c04877708da9b93ebfc9455776a4b8d67eb5616b5e299109e3d4ba803e76b52c7061eb58cd62eeaf49f9152aa5deaecc638039dda60ea9b6e44d8d2e17671cc7f1b6430fc845d6192f2a9c0b56c0afd93cad85eb9a99b20c67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha57b4706006835ba90a7f780298856c0539caf140629ab39c79874233c8d08488e3b3342715e6fe28208931ce5debbd4dfdf5a5c083d48374c224da39770d3be819024b99c3ee6a62ab163dcc4cfec65227228cc86d154240375ab0f5fcb1001241f457ee056e04ef143a6ed1ff8884d35b70a708b2c3556cc41acdbb1278296;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9081ec774c867e74687715b942623bed55b5f834123d713894e5315c25e7c029e35585846bc1d114b5aa7ffd35efea66b4eab3014a00166dbfc9df6d26046bd40543af4f53a2eb03a6777c91795a7c58d00d4bdb03a8be4d823b2e0f7513c3a75032029a25f75df1702a0b454644ab06cec9af596071b9b77215d8afb117b812;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3fe98447a46afd1df6077ebbe79666c1db65969056121c03e109d4a22b9537005e176ca91d37180100560735e6fb387519ba859413c57fd6ba785355d2bcf8ef935d4a6f4216b64f7dd640c02b5966e81bdf358bd0a75d3a80f329e979a9856456dd1bb3b0b191d2363d97d938cd3a0b90c0840d7b77316b8a45c3483ecf56bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd768f57f0bb4eb44bb738bfbe14160c1a5277aa00307376b59a3c29c93cf1957dd6b12e6c08d8937fd8e677a5c73ffc122fc2ea98ed0c1ce7a4334cf3d63a9e7d92d887f395edfbada8cd5d9631281b1a63386093da7dabbe43d03875505f80dcb1af69782d94cfb6e8fd9940657a58c43e00d2d1d986818afef3026dcb61034;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h223519c3a21315d37fac61a681fb586ae3527e9603b57bfa9518e4fab797e5fcef61394adccca100a16c931dd2d7b98a41a7107db5f6cbf8e38ac87a0cdb004596257767a88fd97c9e65ccbf4441363c1a7b44e3ea035ff6ee9727d74465af0280274c14607567997ea3b3f9d2a7237ae6bc1210696a270cba9459673efed946;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he296a972841b10a3a60b381a34657868fd3b23f562ef503c537473c297603fffcb1bacc0cc839e64ec8b4f2f25a133dee7dd35e20e71de7addbcc282707ba63dba0a3aeaa8de86796f2f4ff0a40e8eb52cd091d8d0e3849998cd12313adb0b2120abe383959681c869882bedb96d52d04321b9f1aa3a15278a4d2f5cd38b12b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3253a427c569da77da639f5948ce85b7a5b4c45a95e8e982ecc20213cebd4f3bcc72133b0aed36c90fbcba67bf3026315d2d94e3cfcd7f3f6920eab8b0744dd130cc692ee43235d5439127dc926e5e9c3d360facf8a31033466409e94d8f09b4fccff8867a81f9e6f64927a65e2cd741e550c74e6c8025826910f0d16e477dc2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75dab16be40ab27dbafdcd83429ea8dd7f28d9b96d642a55a2cbd25295f0fd3063f93097b532a8ba1af80f93b8db598f8a7709bd530310f84773f051fcc746932bc74d87102ec33277fb9848b3833ab1a873a1542285b8ddef45edfdb885bf19f81fb74174c80eae932180b6ed3d98b7d75a536100f0bb26afb2cae5d32d03c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4bc928e62524e5a351d68baeb5931996401e93e2928f52dc854abd1be5275d35202de8b8c0a707a8e15e75cdab5fdfc8a87a21b5d593223ce79ffecffa1e7ec59f71561e196e21881a0a5c8ccc8403288343fff771048238dfc821279f7865ca83d7eaf7a54d223c9ae161adcafeb80bbe3302bde39ad18fc8f2c37c0c8bf708;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61d234254220b78d41d4813926eb15f88a304a3429069933f07cd0b83736f4ba4d84f5833a7d03a3be223461c30b78e78d4c3da090e5a169f3e37183b6949e61734ddc466a87c6ea73bd5cc4d1d4840ba25bbdc4e14f969b8fa0c6207381640fd12169d9356de3e36d2c5915f2ca65a9fc3b9c48ced1f859ef6fbc9fdca54140;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h114f1dc35c60c52a8be6ed01fdab87edd1323f72f2f7546e14995b3ca088abb369abf25d8f7fad5244c8ad1f94b8291080f6c0c28136faff52f0c6c9ed08721620114c57cc7a1175debfdfa11a04e10b3d09d0b9663623cc3896705a55512e0d47629e89d6af280afd63550efb9b613143bd5cf80fddfbf486b6779a75f993aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4ade128b244d5716076566ea468f99e6427ed175e54cbf50c79d259547382a3ce60e5da197d5b10304b2a1d3a0b03819d428f436bab971ade8eb2c9eb70eb68de018216026a2c03282d2dcfdd53211c8e15cd31c1a5717b3cb4ed9b0be18923ea19819a89e303dedba364b4de5b99f534b1b3c0472005b5d44bad578a5b05972;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53215811b2f11c6c34cce1b9390054969a4c09f2b416cdf21611164f1eaa373a4942a7113e265336a28762565d53510994596abff88c0716f640673a6a688fdcbc535c77717b2663b1061a5f2e7ec25a1812bacc53be5fc054b3fc05a624f163772a5159b2df064e8fd0404ec0acac02947a13246fab13483927a84509bf2a4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4813aec3c53f95691d95adf41ae7add54e61628666e69a6b8fa6ec1b1d3ffe203ddb2609ce4289e26f74d5bd0e3bb3f9d26861f9c7ca68c5bbf20a53105802b47c52669815d313ad365bfdff13994e7c7566b1beaeffe470d58179867d8dc531d5cd805875de40d26dc712ba8752667fa534c8dd14495d2f4c2d9b90448032d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbbe6d20aa42e212b2db64759987fb74c388eb49ffc6784f8e8a1cc48b49b981b209f758ee4e114bcc904e8aa30e714a4775f810ac11d0009a5b48fb386c22cbb9d2391136fc37c0d9a7e9d02efcf40d1083535df0417be3c1542f47ff02798a382855fb0f739465f08e10cd4fb160d8bc989db9d68cb2c406e76c006903794d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf74030b8423a659b8658ab7d3993c3067ede52e042fb6d6f20a79ffad3d89758f39c44b803ed450ae21392893db40ddff43c7b5c04d3ec2fa8ff9785a166d83d4da86304709149e5838ce47103d71d1e12bae754f1db414ef4f7ac8cf92902f83adfff9edec87fd98d4000838f40721aae12973e5c4351121394ed9957fc657b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c673674991b774553278774d3025d4b71d75a40570a125e805be24a0244cf408e08af98d8de0559c9b5b4c652013c05ea777f2a6cd5f0a865845546482de05516464b407ac48df03854ab3900c16f29ebe66a9629315ed101dacd1a421e3edb3106e25fe69cf27e80c651a17fd4cb6fd4a6cdd68262a57cf0bcc797c417e692;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4371c7f10a6291ba8bc51d412763d8dafc0d0431e67e6c08b620243454f746e7d03e4a990702f6eccfee04f00b5de85ccc545e0928a9b308fbecb8624614c439ca3614fb2c90beaeacb342a0f2ea2e79b58917f7231aa826b8812004e214ccc0302caec6612c3b11e6543a7f088a6a3f50f92554e41947de62993a9e514fbe1a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc439f311e6ba7f83c46bbbebb6b392c3edf4e0e6d0e19971bf278e39e85aa5c20919192287b83212d278e2d82731bb23ad02a346585bee4a31630501b839511a440f9dcbb06262cae97bae4679fe5b7b6215af67b4c23c10ae313ba7f98670c36a059063e89aea80b68ae15404caf64b467672e10557f1ff20f0e7092f0b2caf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3de23ddf362acaac455a66d81fd68b8acae512e78ffad47957fb5a15cd2d3c83e1f839737a312568492a469d62c959be0cb5f46ab421175f3ab602f7ecc0dc506129ba394a92d55d4852f64c0d6180205dc38d63d6d7909023d89add58ca78cec512f2503c9b2df8086c2ba30c3d65cbbc819ae4e9e4ef84e53507dee98c2df1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd753f7e1c88fa33aabcd74dc37b98d1b8f00529f12c80cecb76c47432445ac789ad3bd94210c5e09ef1916d85996db390efc9c359e97fcd18a326811d2f001ef670519eeb05a2a7656e22c3b3ab18a7070c75e58339ca28ce4c92f653228032295d4db470484f64b61c2b728eb8e5bf242074b4bfa01f5fcc73154289db126e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3c6d94e19b57bc5735bdcf7760005d0ef7831d257515f728ebc07d5e998f7cea5d48e14547ef804d2aa356e7251df0a0b03beceefc5d6147830f1d7974f95894c8fca970279b39ec5b9fc4ed8e1cfd40832f5953957c68ccba8596340ca5353b4ff699c4f27d58f7cc9ff045d8c84774ed4a9c56bec90b0d8f37865a5d980f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b42848e73ecd722bd6c93a1d4a359ff264d3d14f2ba0e67f255f4960cc2a2e977aea341204daefdad7b45eb647d6f48b64914934e1fa8e920d9c2f3b1400044469595ab3638fff1fdac8c8db1f7f8dd86163fc89e52563ad611a60accd069e96d82255a965605f092c73b3ece8b8ce790687ee1fc25a4e0a4878e7582ec6f00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43de1de62a340a2a670e457f1541c02f20ede8df32d90f4e16330741b6d7ae0fb42db2419f99d55e1152a84174e140bc3db1f41e15ba53c236f90e0e493646480736a01b28aa787b1841a47578cbac95610ae70ca4238193afe82014ba38470712879afd1eadb9ad04db86a15222a9b507226ef1998e052e7c8ac808aceeb059;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha9c3339cd0e1a790cf2c918c6ab992c10284ecfc02607a87e44763b082ac7e3b1a3c02748713745933427e16d5559aec6f182fea1c398ff290b18879e3cd701c339e9db82916aff7fbf0361c7c7128054f16141cc7286ee4878e5ddd8f003be91fb5209287ccf51af5f141ca03ad0a7d928286cee0ce1c3914dc3818ea8611c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3963eeae5cd78a67bfcf5137871d6b2d7cd2544047d540c781e33f6e595813089710c0acdec73e45d1fc16ce36b5193c1a617d2c2d56bb9741b03b83c438663dc9c6249a3b19b958aa94bffd140be9fbdb1e1090ca904462f58a1db3378f23200254f6423867b9eac367bd864d6645b4db9ff584ff18e5cf05126f408ca460a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4acb3ca60ce4a7183656b63745af971c97c456961984c12241d19ad10aa79c76d93e68ed1660e7113c8bb3c9326e9e2f8f6464381d7c50a7b55bbbe1ecafd3e42aa27edaa0d83e8cc0c7a0c1347088043dfa106e2fe8c35271756eb8372896c1ad3ef902d5e1ed449d080e9e58bef82cf9bccfbde5bd9b93ab6c2a1dbb82eb3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h808d54f01e425a58357b476a88dfde0be0819da2bad305ba0c4327d3470f4d198e569c1b980aae655ea05b12d292304982e6aee8e44ff8cabafc7e9e452b2297a82d445af35cecd95d6cd59fc2f1efce441cea167fb418083cc52523c7ae959978c83bee881ba6dbbb0bb67055c82836ff7b286eaa2c85768ab8f53a05126dc0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14e4aa5fea9c9a94ef0c208b5872ee0678e929946ce60696f818e624aaad4e98d98b58dc927694e2e13c1be5cde3836a49d01afa7ba8792ce3c85f72fa5d2358c7e0f0d8dcc7d113567019ffbb55967fd2aba654eef8700fc0dd5c8d6c32af2e9c30c9b5b18e2bf643b624b56027a6e76f6c22417a62447bf91ce5183d8cfc93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e2307506add987ba6958bf8863f8ed6348dfc53849c636a1674a261b8bfc2b27f767da461083add157b63f93875e4e08208c4115ab1beef8a2eafd07064c83fb79cc69903c4591d590818085dac6f9bf45bdd99c25141aa771293d971fa464c61db48199ae6c5a6d95563180dae2279ad0c2065b47c0e76d3ede25f2ea75ab8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7b07aa4844bff344ce119fef7e4660c1c2b5c314b226a995c2906f7d8d17ce500d427e5a4239236f312d35b8906a848ae7eb7b3d945e88bb9a0ae0d7bcce717775a3a821e904a301757675a340d0976cedd3c4066d88f61550eef29924c6037425f9de6b62c22d3e583079b872f574c0ee7ce179c79433bd84709191e2b8641;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b2b73ca51f9e4060983e1912a8b71172e3948e8c9dea5392fa6df72bb005375723e62d09cb36cd283fceca188d56fdc678758aa75625a6b49104f7b616433475c57cadee7280ef2de61fb3db3fb8d0d2ba4ead0a389343e9773e827eb05c3d3100e6b8b9e324fb0244772c90d7e7e3b0fd96d9512ab7c4100badb059c55cfec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3f57520f637a2f7280bd9cc4facdf62299b53e4beb74cf3f26b261ac0e187a03802d1fe45b97f5d1d11decc5bbf8a31576f0a97a44372478c045da548f2c93bd927926e9cbb4607203928f9afce24febfd2c6d9c17059e66081f2aa8bf83952d474441f309e27d9458bdfcd46cc2943806d22075c642fbea3286d53d97a5d21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h802d648661fcf2320d377fff3029842aa583d2d4c4fc6ae064ed8a9744f84fa69391b542bdd5a9159711b7f3d8f5b40346326e713d47028a49cde58a4793d5ebc6423a2612c3d8f9730b07c8ec1b194b2fe8417211fa851f43b987d1610e7ed01f96746fb53b4c5abd27ae3474777d8142fb17043b43437c8ce6be946e1378af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61fe3ca72da1b2ca6c23f1de038e39acf0b5d9e95989157c4b1218b79abdc59ad35a4380de52db96491ec39070f831d40f5fb107d9ceb4ee51896b544e1164bf76cc991ecdab20378444bab36701b336b8a1c0c082106e2ae50c2c66dbd293bebb3ccd8868adabfe6cac621b5c76cc4e091d2c5edbcfda4e195db4b753dd8077;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7c2481382a5867bc19ece9784825255917b1950611ae1ff755b6d095dae794f5bef58819558c035dae7f33244ad1163f44e15f152d9e1b6a0c57ae3353f26242d9946ac8a8b1363c1a363831a8d7264e6f8b39599abaf4170ff23abd6bb1fc0aa625472731eee3e7b082f57fc9175704bdbf91844c86cdef0433ef782e3dc8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha21a6eb43a91214609d85833d454f872ab89aac4a0ba2d7d99d0ae91c548602e3e6d2ea3849e7329035dd05c2b9f3f1904b2f4663cf24dbc845430cc51c106a6dfef2d2475382ef8e028dfd0203d41180fb36137c0f53a12195f380c59ca260a2d1711cad8c68021cee0dd1abc426654fe9cf547f5f644f3e55091dd4651ce1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17c036823ba1af615385bcabd48b8242e6ccb3c226b53ba235014f8cca5ef8c68232a240b823f911b744704a76d4646d45358d15dbaca71a2620d282061037582a0d1e72adeac8028bf75d9b5f29ac5ff2d43b704ae3bd2b71f3d7bc690f038ce081cf0006e315a4e528bde63fe9e409a26dac32b5254bb224ff90d603919415;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a5e8a5d21e7bd4a656e7f8d110ec94e36469c5a6c0e1140b95d90553069301ee7e07b633f6df9399226fc5f7a1ba55fd59e8372116a6ee4de41b35032e5f8781f59c0b9e5160460145de1aac6436376c3ecc2cdef7e5469947b65246fb0a49137062f6c17958a63039499090d6ee02630021aa50a3f1d6080e94add77d65c8a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ed67abbf1f4fbc3c270c61cb4661d362bb5feb341e6cffda63842ec72fd723484f305a2c26af0e636f7aba6aa175dbe455a3d126d775ddc6b8ea5b2a2baf56e4dea90b9d4d893576cbd389b961d818b0dc9e4dbb76e9ed2fc711a2a0ecd4adcd4d87323741f377e6469450fe0e929db523b9ff67f58bd89884b17561359199b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9af26cbdc3943c80f7911efad6fd1a7de2bdf9391db4f7a7f4891c93e216f97d8fdcaca61bc7784fc2879b10b01bb8df9b76c066391149c1c4f5adad9d66992d5255732308f85f24c4c7ff5dc7c8f1a9f9f710d53e3da7e85eed724ffe4fd42fb83e08e434855de89eabeb578262c102521853417fb72f5a825148ae54ec08b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1aac6f4ffd4c63a2627d1d5658cae279c08852cb949cb395b926b3f5292a78cc578cdbf4b56988f08b5c1d91f1dd168cd50e07ea3d802a45c2c8ed01cfcb67475f50d9b925310b23414eeea039300e6e382ce42ccc8ce27f23c0bcd675b726a7c03c30727bc42d1106af8f319fde42e1a76488ce3494e3db596646c458f615b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd56f97530e0e2643a0ed332487f581caae82f382cd885731c3e94629f51c30327eba55ad613c6d75753b2fb72308a2f9fa0f17711dbadb9a9660da090a059d6bef86c54c12d7571dd20dcadd829f96fbc81e222a4f72f72dca7061f9a74112d44adaf00185088d7e54b4cc60073d700dfae768b81e6f1bcf840fad6ffa650042;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb13543427cc0d6ac98d9fedf20976d5ab7cd7a66b052404d3d0549258aea85a16c31b217f300ad38de98f24aecd01106dfd2f93f10b488da1b3f491dc4533ec9f3438cec6d219f889fb230762234b89eaf38b6f3d159aff0dee3c220bf76905a06ebe2fd61a31b436b247dbaf4e99918772d58b0d9e36929902b737dda2b391;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13fd2ad62df18685b673a0185c138bf3da6ec03ffb8d4cc5bcb70f7b0ab6cfd2595af90539e210199a9855e2836cf9b2ee663c435b4d57dda0bb10b8cec2890d60378894f46b9f5f66587aeae02c0f2b094b5546f4541226a1a25658ae65b98e26ce93c4adb837a18bb6b1e8433154551beb9db79c66c080ce631e2a84f11606;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21dd2db6a81fef0370839c3ac9e9e0e6ef3420a6cab44e8e0c97d4f3db8ef3b8151649cc2cdd5bafcb02167451a66b0e6d2374a093a633ad8cdf44b52d032256684afe0cab1e559cc94131d1c7b6dfda36ecc9412eae26238261d20133951a92ac3f329a55af13e0cc65b813209e59270cc55269b99ac15a2e16c2e0743a6ed9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28c3d4e1919bdca0390fc1b069378217f16384465b703d67735de31d4039221958d2bfe6bf9147ef4ddc67edc010b9f01ca11b9d069d9c42bf4218934954c230f907fea17a63e5fc374424b3d6a73384960df9670d0d4c5665ad64aeae7910c6fe2b07953e48952b966b031f09d3cb2316604c583cab0e940d8297e1928acbe4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e1e60b1920d40d8a0ea9ea260d928be0e8a43fa435f6a89b3847cc1a142bf8a3cf8d7e4645d6fe3a79e53f6a40da2b04b37345f3bf7bc74c62a374bed1cb1adeb16f12f7f652304a52692dc8be9bd07e121164a9e3ea1e5518d0dd1f786689444d079873462eb14e4e4295f100e97a2748d4a168d46e601b729c62b493a3d3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h930e2e92c8cc45053e692266421c9acffeba95ec78dac706c00eb67c1d3938f3c11def2bc67e7c87b43dc25f5294ab7370dad9c4f181d39c5133cbeec21e118cff1a34ac656a5010a8ecef34a28b794db0b863e01a06cb13c5896d6f82e58e56a898bf71a2373754558419d5422886a9bf6b4d47b7811ad5c87a59c8b9b48da3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2979d66e88f0b010676e6870c6fd93093b423f90fed4898f674805de8b8eaed545225164fbb6bb5600f7105e518d1d9deb060f50c3ecddf73366fc1c3689c66100905c3fe11274c0faf6f490d1586e438a86714d0b0e4cf5871df3151826b3dd7355c64deefec4c1209f144035b68afd3eef3cf2643a9cc5585646a68839df2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8d2fdea675280b76bda9e599e22769d87d7a05b94690da01aa1733c06bcbbeb67e1ef0b109421eb3f2caa200fc3b14b3f0b8e5699ca8d60de36b2000178a524cd98137aa11b536cfea4efbef6fa6e768220925f6b80ae795d2bbac4b47c566c1a7a8394d1fca5ace014245aa4f87c21907a5c8bd992d6ef8f20609ae47d5c2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6399591bd414ef985e8091988e612d8c59ee58bd451f8b19faf8c3eb00c9ddc90ddac062ef921acba1e07956c350ccb3b7a54fb6004c77dffc5ae58df62f3070bca86ef4d088ad0372f2f18e5bcec4123fc1d2b9b951602329e8e0e9700911016871940f6244c45cf75495c439551ad0e7dd628792f0f2ade7c446f62956385;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48e66c602d5507f506a9e68a344e0d6395f087adaac08018c2e3fdfcc2abe9fe2dfe3ada295fe8c961490cc87848f7d89bbe0a22685b706ed10357fc30658697832e1f6d0fbd647f9d8c029250ba77fc8a00046fc492cc413a30065bc5879d97ae34d28315d12f91a93cb8f8cbc3ed57e68e160bbda91bd3140a0d3d76f885b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2a17879a4ef52b919e2f69f349d12f6f3f725785f803ddb7d5325c877dd7b43059aec168de6c460bd80edb09650fe6d2f4fddbf6136126edc25ca07c9f1c929b2911182bacf31ce825e309836aa82ac19f40f34ab5852fadb716000e2c1e4781d671a2feb545fde472d8fb402a9d18489dac8f54393828e3d1114718a7e379c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87ba0530fe1f3ab486fadb90c08b744479f00110d14c1ead2dc7635b83bf1d8727ec7a2280e176f91e371c11d049a542e9ed5fc95f042b33f28b322783b89d27c4a650be1e4de0ca6eafe35a8ee44b27e63f7502b946c471c8193f65949fbdd8501304f92e84ed637741f5673cda79d6b83e2a75fcb49735ecda8b125d2dbfde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ab48c1ba7c9831b079931755bec8d9ff120faf82f364afc8dba7a992036045f47f8d47cc8d8f507f6ee35d036d7e95c97c3e53ec60eaea2ecd6e382303c1d04fe96b991b4f2b14b0fd482d8b0ec48b597093a5f9d5f79328da67dc740f8ebff1a9fb02b2c46e11fc8e25f4afb0c6f67a35cbf0a4587603df03bf3d5102cbab5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3b4fded290445e38c13503e26d998b8d8ba746d35ad7f9c45d0a8d822e7e391bee0d2b63262354773db58259d3b72e02209b6f3fa3fb6900e902a4839f56a27382c82a4bfa27e3d06219a8884840eb522061183c6807f14fa6f040e21ccdfc421dcf6c635c11df3d2656637e10fe31b5f16fd632827b66b9630b8b7c7932a5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd73f63808830f33fbeb8e94bc66b69f0aa797d4494712888adc2b977e749710de98a415408e4ba68cad8385d1fe178d0f51f42d587bc845990f4818364b635ea36ae0894c520593cc80d9db3f5a8270f35aaa5cc6170fd6aceda6f1076d11b53d221d3281c71da6760d7c16e0795609a7acf316af4cb7c754a523727ba3a337;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61fd8b255e1a793c37170a39d2f7013ab4157ee1409e24004e86629d7d1cd5349bd8da9c2d6394319f9a4117ba90ef1ea9a3f2de1abee85ce0ddc1b3ed8925ca84739edc7f5cd6c197a66dfd068242e5f559fccd3a448a4602c89e1582d25a8985a02b5f86f76e4458c69ced89eb6369d5c2684bbebbc846d33a218c70956e63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h431a7686ccd8f8436c002ce93765c411a4952316657cdb024588726bba0bad717171590235ad9898486350a69e28ff5dbbc0cbba174670bd6f961224a63b8de5d14b31fa808f2513d90c8487636f3d360d90162cb594ae23aaecfeda5a948fa1d56377996b0e01a28ed5396a6cf5a9aaff2bfd4af8aaaa8a37862ca73b69b03b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5804411f825cea44ee94074291dbbe7e7d3bf90cbcf4d270a3b699eb5d59bfa0dcb76e2cc3a3d4868d5392937249bdd8fb5dbe279c85a4afd8d22e1f820614b172e73f8d8fd0f1f8024ce5641410b90677a7ab92daf6af175e2f82c13f7eea9e83d8f4e4c71172b907a752c012979dfd1823783cc3fc9b70004dc12ab52934c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11b99f9a7be8cf5c4c9cc51936809c57987f4bbd156db8bd9f8b75e7194bb39f39b9d78651ad9d4cea1a427fd7581a93fbfb281f2f5cccfaf52b9232e6a08d45ff8c20e31b3c9edd7c17f3be4bce570486f1ef7cdc388416cb8c3b96813f98d8106884465087565518b79bcdf796f91ba0da917a5b4bc969911d3def77c4d3c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9e8ed825a5d8514c46e150fae03d50cbbfd12dd6865d07a12e02c16dfe516d15a3c5f3cc507ae3e8313b14febd581fb5b3fff07715409f7aca32359acabd23d8736f532a29cac05de5b689081644ed95350f088c7ac035907b1d47bf4f0aacdcb4390d9018c752d75345087f92594148fc25afbc9ddec5d1a6296d57aa30482;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h295eb3515b665491658e424b271d5e7d8d24ab7ba821c2778fa886be205ebf8be2383d3af3ba76658d2197a0dfa28ad9be25c8f7b4f0eb873f2adb747f94a2e68d84b250e28444713834e9eef6efc5e04d4b1e5f651cbcee14819b2484eb83af94eff0aa7e18dd010a6cbcb15a20f90eba4f702b0976fd8dbbef824d7f18f7a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe94be2f5a95ff1d6b162e2e0b104027e832b289b0549f7c251bcb4e797e0ca4b84798c5643f059f5c8be8312e72b4435489a0ca7fe3c4c84fcdcab28a1afcaaf70f32f37fe1d92d0f6a66c34e4ff63c5255a85f5c1fd557ce110937014c5148430dbaac216f662190dff47b18853091f57be6748bd77a9828e4ed1d6e269aad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb12de008fc7304e99c3cfde8ee859ddd3de1efe486d886ad0d6ae6aaade96db29fae38213c514660199d20c19f53a31a58774327f257b6292d86033cafbe6bfd949ef2b6fe9219543cd62fc61ee32fa25b24829551776de81b91e705b73c58306db74cc5899c6136f0ae8399bcc0d236bea3c04410456cb565f40a5222ba0ba3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8fdeb1833bb4dfbff872fa04e73b6471153bd20c908acb5b5490e71ee12f63dd47d9c15cac62becabe79863638a10bb8cb2c5c3ac7beb16b594367cc4bb0875afc1de6997bc030dc050f29a8299e7af0c4686cfac58ceae26babddc33b33bd10ba755613a5fb7d57c148e7a5e135c419c98d462f690221821ec154cc6389995;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf1c0327e00337d695c3d3de3b1106bc5b75f7e78c4f3d322c06471968766150350ae3769ea15ff52f859cc1817503266e00a6bb53d1939acb0e6487a675d9f00bbed1047df288919d028658de20a92756049433e6b6f96534c1de532a25fcd2719514cb1bbc3ed4898835ab939b46a1e041ebb7e2d1307a20b077011fedc816;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d86a4a45b4312b6c2022a2db15293247ab2f86436f61805d55c4f51637bee8e16f80aad933a69ba567a6d8fb11fb5fcd06469268c2211409b4b064b38ef2d51f36ff8af72764d1983e56f909f89b56e13b4c6d1082839d9475e8df6d9874e0ebf9c928b55b5287a83462e22dc0b951d0be05f17c5cd573f70f5d6efb1be99f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h500f221aa4a9602489a989c4f8ec962e27456a13f9fe47cca2c749b3d16e3ffde3a0c3f69a0bf5ee0b79d63260223a8212f1b17f11147c3a7d7734920e94536637a54576249610e28407432e626292e59713967336e06d2d0b6225dfc50e5cea4eccb969ef4a4f543330de1d0e5f7bfe02d255c8fb33e34ef1eb2a81ca2e9a9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21bd6084c7c08662725191649b983d2b0128846d1998264e019df1375280bc96345de830d7d9747794b4b5438d013c7194385c71a8c501f8d4e43ca799c87ba80f69973bc349049e1f7c47094f48f4940baaafd2e14b3fa91f0dd3731bb4ab5cae4bce8a3d8ff4349db6801fc64d817bea3045ff3359b43b2dc511e41cf93e71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h728ba375daba08a005530989a4044fa9859764081ee0d6da97400db02e5e54d2f879bb22064ba9bb155e1f0af726435f36b3cfab500fedb77735782650500bf588b06e3e5d5a05436faaf2a739029e0903e448e3e9b1e9a54497ae18fbe56e39a3718b6d5988bc98a2705d4aa609624e82022602883c73f19d0620a1b74d2395;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e2c18550cb7a6630b1d0aa9179721f134d980275707269e33d4cc0e325fa86f15e147418e0658e0173b8353cdff8c0590f1512d4e7afbc2878b0c631fc020541ae44613b26f4867b081d7dac4c27645c853b79b04893fca8961bde8ccb00ca22484448243fd7bcbc11ef8cfb34effde6a572f8f515e986d3102fb15f9313a99;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6648670d8a5fd0b8f5bafee3a5c5d3d756fc92346c1303b5927aab8656109f49ec244bec661c2844b3c2f7d50ba61cae1bd5de9b429cc6614bb8424f83222a4d9cfe64bbb631d754867dacfbb21f00e6ae75934abd39a5c0abb8f915b88003b0fc3a60c53977ad3bfc2286db3406e1f4f52e2ddf50258fcffeb8c856770044dd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0c56b49ff4d5c20dbfd5f6cdcf762b5a5c4af92af1c639aff9af2d79de99a54e907529b6f8c106a83141cccc2d565fcd5765ab752a66a96c45d108e420a81a35f3be474e29b4a0fdbd343ceecc528c496f6f7eb51f1907b4d4d5ea8c6e711b637f6bc6377d860ef40b34ed121c96919254223ed9a9cee1b43f974df83ced22c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4c2b242f0efe563b31b65150bd89cd70a5619f24f44179e9889a1d8f0acd5bc0293acc7f54f8c30423a7a561d56dfc47c8bfbe13bd1b11065d30e8edf16703ea3ead946b3fddbbb1904b3135afc6339315ddd7c9cf0347bfeb55fd3ed9e09dd6e9671dfd81118d4abde3277a8c494c9265668b8966196c4172562ef646d396a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he185de902a66081945a5fab12c57150be0bf81f76683be41c3d46030616408cfc97c5f6cd85c73a734d0e4018763ea2309bd5c80c64267fca24d44bc7440094daa879018df502d00083a5ae2935ca3f986ebfb0d13884da792a4e8d2b4cfa707c6af70d6f5b9a4ed3f2aaee7f35d3e0f84dbc3f286356d75a526a1d7a4fc0733;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f97330a1ff380ddc09e1213770b754fcd0ecaa967bc8e4c60ddc200474e7275ac6005596050f00b892e0fbcc128b4ea446e087754007652478d9497a52e4e5a05a66e9e46334c52f780b6701c362f45c86fb620e8db61d443f652bba6bf7fce4c19ae9068d0b3e1778425b68e369054bcc96cf831dd3b82f577fa7e655934e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h16dfadb7dd7309bfab5e4c03d0d905b8bae26998e1986ae1437012ac0bf3c923901472ca1d01042b44c8cb95f9f0a6b08f475a6ab7a17585fdcf668f5b5fa4c9be7be0d293bdbe6acfa47988fc4221437618e74726323ccda819ff90c39d14465eac2a5a2ee3542544d59686e74abab5397b3c1bf856c05989a26cccec6262f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f4319f924385dc6a99cee4205dcac5c2ae5a6104aa684c1953d6f8cf7037d64416c1d01ed1ca13950181230d5f7f1b8c32145b2f78d810a40234708106c69e8478b6fcbf936155b40887e05d48eab1011dce08176463d8592d61416ba9b324b0de3d794450f04b48944330d826f3d964000d87b2f370b20a59172e329aad0c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61035de8ee163895904bf22924144cf64f1f547ad65b79f976d8db127b7c25f6dfbb71f6c795d69245454a782bfccac693fe48d9d22fad5811cd92e9524802784aef0adb20f55be7e3ece08ce2e88df8d744568c0c8f837f578ec2263cd748f4032931726312fa0c0185aa919f8cc4ddb5d21f5c7df112238fff5fb84250baf7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf97b6ae63f3c899b677a1fc5a61029c7179265f4dc8b4128ebcc72b9aa0032dbf4a95238fdd5795e017145814bb75c0b32b2b28ac0a236f1bf3baa3e94b01bfe7e86d7c9f8d85f9dd998d32c93538e54591b6c83d9ff3e3d6d12c65332fa5034e84caf78df93b35238705b150e2e2b11e09df96bb8bfcd8ac5c7a033366318a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf33b9c71a23ebefd932f089eafa84542c911bd9c39dfb5cb1ea7f4f28c55d4ff0c78e5992da074e07f57b34515e2da131908aeab0aca45b464f64378b5c18541ef63b55fd44bdf7a4cd072d3d1375d9aa29f251966a535980e02d5de72f7f2bced82d868f8a6c6163881745a6873bd499b23eb84dc2476a9ee476868f2676992;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a5d81e2f63083132fc226b8cb45af3b13fed84e649e1842be43efc5ac136f14b4253674dbeb8ace9156a6015b0768e91205567637f86885628f1d2f7c3ceccb3300fee4fc6903d17c64832ac3780c4e8a7d824f9cb9a33d5e8c7abd616d3aa6ad0080287ac5071bf191c78a41acbfa2ad6c6fc70a25470b6fa78d2acf1c98f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a6c1cea4a0b2ef860a42560d8b6115b9c40a9c4cf147bcabdd4f300a0310b5d5b46d289cc164e2f09a0bb53f228c0c156ed06c2ebc83a77c7aff3a34be0ffaa2039a9051ce249cbc2f251d151e0ac25635048fa7988ecf275c7fdb1aae09711708827e334972b9cf8290e9c91754491a8d9a9e264833f32439402847b5e7689;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he78ac9aceceea0fc4e733add63d440b69c8dee7d520d5b261da253d0a89a1496f576b862e256c5cb4a22b08764c542e6a4f4b6ef065c95db436dd45b7a4492176d29c188d091f3652087cd6fc52bab6e8eedf16945ac2d32c38d6a8170b79fa3802cba71b613badbb99238fd360ed3910f3ee8645fcd5ca8b23b3bd9de4be57f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4546ff3f2f55e3de929c853f736034b606de44458f0707faf1fc64a31804c4fbf9b08b1df3197d114e8c98ec086ff957f6057351627e33a630212dacfed1b1aef42ea48e0d51ff9138b169607faca3c0472d0d82d61cc439df12073b14c1121d94e6295b8790fed28ee36f967266d1a10f0e3be5212f9edf9f51a79a47c47ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h159a28d0fee8670c11976844461192f547c01cc852aea598a06920661a259ff7866876bec9e13c76859863a2b85da0f9695d3a57a607c7602c1e5de1cd84d5bc07b0e9e72c2dcc4e43ef276fe0066b48fb2d1fff7155c2ae53ce20e2007c8ebe277285ef39182b57ae6e71da4392c1a61a29007d4168bbadc93302b91069d996;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c2e121881d53dd9167227521be776a13263b2700adebba3a6623be85f8a703ea67d76d2e587ace92064533c3b78af830a3f82921b02cfa8d9189aa22e930b76fe26d4b37d950a87597ba9a0a60311c3ab05f18fa12973826a08dcbea4c3811f1e1c19f86774066fae1086a1da0f74262c78d763e44e94ef459c11d5bfe55b24;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e5078c364dca65bc81bc6d8cba07ab84e9a5ad7fd97cf3eb700c19b204a0474b351daf2ffa1dd777e3a7a55d2e45bff9140a2f9e9e29adca3c3df28d6eda431669f5b7f6333a451e00c8bcc53bd31544fdd43cc3d96db1ffb311d2e3c42ca4823eba68391483b3f5613ca73df5d81fe590cc33b754a84cdaf598cb7c73a0888;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd5406df09f43d02ccc507c37a8f2a31015fc4e1a491252b748f756a774868f896cccb155a3c54899dcda953628cdffbad3be1ee5fd0c84d7ac4d367d031ff0a4b72cb579b94fd53003340ed976dd2897eab714ae3787ac3fbf891e7871c118ed89486766e57382f387cd750b2f7159a138cdbe8b3c3dc8e5b9535a46f89ab41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff8caaa175162b887ea5c0d0f043d9dcb68d196e403d8e88013a5b9d1e93edad05d40ca2b9880d2cb281ad631d8380cbdd28cb4bb7c41899af825fe350e5842037890ea28b69f4f8888271c9a1d4d12e448f575f3277cf07c5ca36cc9363a7b596d409a35b50b73e140c2624afd32c03c3194e635cb943025b876f9ad7a9cf05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heba7b47e07427d10f00dc99445fb42032c1244c35178f36753820d51f768a0525684058485c9a8a8dfec9ecfda5ed8cf1244e00988a1de6a998b847044f2feedb55ece8e1be601bc873c903f616aa076f4c7365cf310374b11a7f81e06b80c0611eb236dfd546a2fea71d4510478f1f13e0292041224332087a504bd0fe2f750;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a3d086a95789724b8a8125945ef005fdd0d074ffc4de521450a12b17401d1b820db1ac9f1523e333c567881f0f8322c60f95e2aaa05da7afa56ee9175dc20972cb6c89a9fc1b2e0b0f3d871fb8318909f5eda996190b4f769871655fb82f8173831419dddc559188409442ecd2bea1afd57fa1575c30156f37b254eeaa5fd00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22e915cec2cdc0ea5016f11739d351e809dbf956259cd68ee8f4b010674a1cc6afad28541ce78093203b5e4097dfba195a31030fd5cf6874461ea78f584a52be33b813ab4c24b8a72cf3c9f052cd1dc7cdf815fce747bc8348cda7e7ff663716d46d41106d143c548a5b61f197ec9dce760616f2913bcd2b4a1f76c98bd115fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c643b9c15fc18b48c9999d31a31c1552f528d2e3e8d80b0407cdad2abc502fd05bc871762b178d6af45b5f0dc01146746d8518d774c3d707ab16d2df9a062c24f75ed48ef4cd5f6486bf414a239c914c80269d08fe57742a755b0538988036ea50e77b964483d173b078d9b31bc08ede2331b9b4a55a674a9af65f840cb5984;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9151ae62e2bff74745da2666af5ec807313e2fb3fa27dfc2f00fc0da2e8a578b52180cc4d1240702adf3fbc908d9f5c452740cd6c2e44c5ec160977ae41b99b267d7221b4934dc511a7b36e23bbe8fc4951a1b9881092c7d9fea729731c580781b9e2dcf28b9bf5bcd7ed5472b4082533eb9a01e89eedcf179a560658621930e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h362a656f7f088905f5ea39d130017fbfef32023ec793fa1c6313599373aeba4385c7c07ec8801f4d7d3f0de8f4f4d4e4c53b86b2dff43268dc309b7123a671263bfe9118344a005b22d68575bb3483f55faddaa476567373a8f7603c30ce5aee0ca55368ddd638c4eb88e76fac9f02560c099c6ade3f51906c0f18399b7cb38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73dab077c99c51359564808073a37e455cff60d2a73f23eac5d6b6895c6749add9b51a07fe92ec7a067d815f62085a194eafdc34fb6e6ea23da4bfc67afb7a1080ecd7ab003ed1f38c412e711a6d7ea29077a52313cb4248abb35de5045e7a9cb3e50649a3726e2a92b525af059ec024daa73e193db77bdbaabf9b9ccaf1867d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he401b28f29d7037fe00767ceb93689745e451688800bb880aa6aea866f5aad701ebbdf2e7f923be45506cc3f1c00924babafea0674f3c1f756f656c1e5f41d488d7f59d180cbc9b41ca0f821653cda3332b8cd3dcd01a8215c2382c9e6b2bf03403c3a4e18af12a18032a3524d36daf3e96ce356aac934977c4ae82c1b7891ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he965f4254fe8595f6fad79fc1d1d8517b3b5d0dba2793eae7045d808b6c5b59dcb8457d019e6f44bc29b2c4e03316882f1c8d974234f180f2e6173d891ccf59812ba924453ef8c1283ca9e008f9e5c3d253d71b5605445024c836b5afb401b1a1288a51bcb95aba66e20b374ba0ed35893abea2b00ef1bbf96aef6900e5aed28;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf37e5cc83750c61fa0af0c4afcf8ccaf6259f40274565c4213c5221a25ae86b9709384af0d77d2b01388528a0bc1fd016a4cd128fc019310761862e13d173096ae9936225e3cb1f573bd05c3cd103783befa5295fda8e3de658baa6cebd7a159326026a9c63730bff1f593f7019654564086a80c569e6efd27f549e00651b540;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd2f4f5f9e2c9d759d49666d7ac884153186bc7bd572ca21acdfd8f1be26bcb68196161e6793db6871faf0590eaf069d0a960c3ac705cc6aa5ec530da6c2105e3b042e1b21a2046913e5f43e4fa8e01a650abd3ffab6e88f9e5cc883476b72f766c6b03c9f4fe2ae02c9558ae6e76735eecf1d5e6bcfd68dbec4acf2ec59129d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5294ba2e57095710731481743b53cf36c21f0fe2eaa9ab654b01d728eb2f94071e1b3ced78666307902574e16636639dff4fdfee95c0c249ea5e93313d8c569fe2b5cf2c4138c04e6c385367618c8b52cb20d5cf98fcac95138f3bc8a41bb163eb4807ed612cc37f5b9134ca6728d6b8d237f02567e4574706e7fc7c5a796dbe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h475b58b0fcc31fae0cfa3194766fd30532747905e3c09bed7a7a962ec8041fe40bf565c4a37f63eeee815a6e6f30d7c8e665517b55179c3c81a5857d3120b45431d277b7b8249f94e6185f80540908573ee8487f7c0d6545f52c2a116ce0ab8f5e8ecff947b2fb1cccef5907a0f96b3ebff83bc1a3e34d4a00c7b4ce738813a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf71e3504cc1fd7af588c5fa8dc553a498b5344c4cfdceed191ea330a1d70c35656a2937a19c5c2928e0fd90e6ee0b32004caf3b1cc3bf23c2ad66a0e9616d8ecb3b0257d64c1d9ba8e194478eb834b0f8a32e433c80255474e170b9be23c56a2575ad83ede2f16fe33fb6023d7549ebd3192b986efda9271cf0db3a8f7c2b603;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfee9262708dc373bffcd19484371d18cf5dcb379b32f87a854c3959c7ab2295cf5a089f6e3fd4df7be17ef85aae154f8fb06f4ec0c8cc2f13f621700565bc89c2a7d7fe6486d2a114c5567a57f43da9bd5feca2db63dc2b0e1b119b9ea0577467ae5a8880f8c8304926266caca082d4c5b586c0af261e52da50ac6c8ad9a61e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf980926c14ac4cdec7b981e2713c2b5d02c07cd0c6cd173ffa6275e3a994d063e8501320513f629b7db15901512b51dd1d11a1a6215716d478a9a506bd87af56b9bb4dd5e34eaef76954490826f47345bc0b1c0b95aa64c35b8e5fb25f3c0035f5e7e1e416e623df8abe2ed8b80d41abbf510e0a5e56cf6c74a1c8edd7b1761;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6921d5fcb0823c2174ab3bb8ad026ce0cda6b920d15b4550242317ffb8f95bdfe134b52b2d72b4d3cea244bbb7a904de0f24f05cd8dd3a9133c1d7aaba1a8cd444c78a973beae4923053bdde4dcfd61b04188429df71cc0c44cb6a6cda2d9a673eaa972788845346a45d2eaa79c3dcdc5d70664271cf4d490489efeb16628837;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7f7a86eba836119247752e2827a92d4bdcb117ea97690c56dab0c424651b118c199b2ebc217860f0a9b90a61285ecbc0da2471e97dad912a80d1b971d9b71b1a166a7541885d57e1cdf7529f040e160c6a49557e929de0d0820374eba515ac2d7596ffb8e4a3a8a0cb6a1d011bfd4fe5aedf7b2de172e12723de2efe8e8f7f5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcbea41651ad22bd04f967381f45c9bbee8174b6bd190673ccfac673024fbe4929824af6f0b352b763a8e7468eef3537ad889e1d2717fad6a7716174e8cab3935c4f769dfa16c2d10583cfab0017e541ae561881b12786a00e430cf67b6b8584a954927d104ee3d2d8cc20c5b7f1d34d5d957465b4296357fca6ef8c1c0aed06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69cd94df71695d31904c5c2c00aa1d17e663537ab50d6e9a32cd2e3b159c9bd83bdc8cf738205c5f85a1b78f69ccaff442c448d7e807fdcd28fd72e847701387543c4ff45378bfdc89feb2ebe9d198b13e60c0520f431478f3a27b6d856b5fb86a336a8d02c7589df00a42e83c1e37446aed0d80128e7c0bffb883e4051af456;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58802f69e589332ef02c49bfed9f1968798966c2cf1fc9b1adf24156161da04b9cdd47f7e7a3b7bead9f815eeee701cee86f674a0bb9a8f5a62dafa54ab948f85265095754ef5123c3f296e237bbf77e0e7de1b3f892f0f5b1826cfdb1530aced97e354ab9e3b3d5d8f25c57bcfbdbba5d7fe096e81d6a67255e13b4dd44d309;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46de3fc00e512f9d965ec505cbfd086079775c6e116c08cc12e4e97ab94272807a620ddb591ac754a5916a833f5a453faad0a088750255081da17b1bf142d1e353ffe1815f05aabde773502abe3b02ff5f389850aff72b8d6c28964526bcb042b61c61d19369e9b8bf8dde0259abb0a0e628635489d9aa2545ae16277c6d4a9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bfba5b2d073a1eef0ebcb2f11ca338670f660ba75827044d155199b4308e653f7d46313592e90e6897e3f67f941b8055e8e132e3fddf5b33bed7290b43af6d5e72580cec3a3ab2717b942018088a2a4d8fc42c16dd03990c8c75531548d94f83896a4a427b9c18ce708e32bae4955af9b9d1a92919c1c8c71c01c147333c0bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2213ed4acc969aeda862850239936a91749a17f2e1fda870e688188054ba554921e13d0ab870a3c2185a250e999514f9e04feb8a160e74dc093f9c3f11e7a7dc45f87a1a3881a30ac37ee53e8ab9230afd0af904242c0d8588ad7b14afb503282da51368fd67f24689a7f46dab96035c75de5cedcf56e657119f67036c3632c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2ad73dbbf564189d6b0ffd690d925eb283cc8f8d0d5b876b455e8cf9d1a361154e7be43f6c8ee5061b1f55bd0c30b99769585e729c10188377f5d716a52f66989f221f4cc6fd06d756c98cf0a0fb6f36335230e3ff61a4fb5d9def8565db8722537f8a11dec9e2a532b264f05c27f438206673ce9d8625faa14ffb30f0e7553;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ccd06c9b16b96e5808699661a2153e69a1492051528f1d5b407898962fd9c1295ce9356aee15226771deee6c07ef630891cac6f8d248b4adc53cf405c9e86566fe006dea788080b476b3a30d90431ea69d3e3a29eeaab08a9c233a77b4e53b54d075ca790e90abc02ad6e537434f3c52ec4ed135038fabbd86b1b44c24a3e4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35f7400e906f3e80e518ac524e8b8fe141aa3961147ea01065991495512dd054a765958c019a4f8168123883f66c7ec1b6f88bf9116c42c56a11e46fe8713b297a8d351ef25898d04e8244c61d5cf3ef3eb54ba1488208ee7355cce75323c68ccc5ce0c58562c8cf42d843897d73c013116f2d0a699172dc213dc96aea7a68c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6ced9aa3251cc13190fc3b61ad8de5baafed3cd638409b6c9c502928e9dccf3279302bcb74a898be04f6729f9e821d48166f8da97198c0217c7d7e53f3939adab20b67140384812f25165e420750494f63559d7574cf23c60e294c6b7d315388bd33f03a3da74c34464be9cec023f3072e865684abdeb91529cc24b599389b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19c1b4c0e4dbd2721b14f89ce8559badb2efdd8dfb310dd0f2a45f6b12272f2dbca28f6db4203e781516e39044a6e305a303bef3ec5c76a3ec935d7fb93c4071bf0b8bf11d7d6fe21dd3160af56a411ad210a38d64e0ce9a0eda4a54ae4af0fbf8b07aa5554029aaee579e2497510ce23bd4b984061f05e2b80e98fa91dc627;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0b90fc9cf824b72812672721eb87e9e0f11a194ba2e90236939c93cd6e5ab71705c3abfc4d21166a5f2be2b75d17625458f61e77d16ec45b80c24609d7929be15989e28282fc12a1b5f4981725cc47c9a8799fccbb5dafddc10ff0988e40f30dcf0ce63de057471318789248049401af2c18a5b1f1e81d357db9ecfae2d26e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca44e256de8d99f70db235e9cf4459c1adc25d2a7c642e4fdb5e7611b20c16f2d53072066fd090e1143f8e6c34ace8b9f7829f7555cedbdbe9859549e3a63648d824ce0568c785b020c6f509f318cf3b3d1d9ebd0b33f1b514c41d89d868bf4b087962df895073487d85a0e668e3dfbc23e4000771e5e4844e1068b2d6c20604;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd305f9b96eb7a2c6da74bcee15e818fb1accf105083ce8e3411e49ac38184eb44aa8286e1c19a33575400568aa35ab7d288f219ef84f4b238d4745a644f325f1bb0e16d7685aae1b35b0ac162adf16b1da1cd7b4b5d48963d126ccbddc3cb9576b1f6c0d194a98f4b020612f8ab61715e517b63b355838fb87063585d07f22;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b3b6e38eab1e277a0c0196fc26c4b5f759ac28692c358f2e4555656b22069599a5099403f15914c28822f634a80cdeeb0290aed190ba7515d3b31ddfecc271badbb6b3a6145d488f6cccf2b23e7a09ef51ea82eeb6ac0ac251524680d6f03aa016e03faa20bc20d030ea3d89c907e148b75bc45e005795cceea7470a59fe825;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h845493244e784f68a722b5ae6e0fa1c42486a0910087ae17f4f4b0bb46b5e291c74ffd539eab66be4a985d9e44285f5f204f4ebd7cd7679507993209643b02b463511b9c6cc1a245fcadf9a196934d1d48b78e620c063dea4716af951e70532d4da6a390a0e6bdf21cd5ce3e43454bc54b3e5bc19499e3af051ae0e72534ca0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d8315c3e657867e108ee09f9839241ef55a957edd7f9d5fe4a78b0f60903f1a446da736100f3e840983024eab0104b4b9b1306a35f4ecd30db799ba84eb94a27ad6fad50b7aeef12c41a0e4f53ff081d6cccec9cdb211a01d14747c5b577ac9e48e481aab2c9280e4be661d76bde01ebd7933715bd87e2fd03da9508a209a62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e6639293047dbdd9ea1bbba8cf24ac84748a1b7e766579daacc188176710e703a34cdb7c12cc1024150689c461cf40c736171e9880a00da35638ddb78e616a387c2e92f746eb84454f63d03ead6ff020ac0eee311deb600e96c4caf3d238370dc7b4f05b66a1ed4f69fcdacca17cb6fd720eb1b477f05d14e80b4f8bc68134c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b1ae9cb8a7ae1412d0c29d817b698a4e7c0ee947fde64129dc341a4960b0e087dffb786395d8af0e4f49aa51ccaf7d3ff21fd4ac9df0438feac3bac6bd72bb16e05335ef8e3b635f1717e88e6b712ef834499310c6586a0a88bc0aa173c8edd3e235f7f56e76b6fa8a0a2fe6fc2a953aa76cb091eba1d0b83e3741ede043c55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef9e999fe8eb40943f76453b43a0fec628aa0846d80c1f10aa3bbb103c9dcdad61195bd8cccd98e801e0599054dc67e9f8fbdac8e7fb1ce4d1499a8dbcea1a9bcd5d65a4e465d101570d4e79873bc28ff2fe3fa5373a1fd97bcaece6801c42a3f6b7611a1f2faef1cfe84c5b2bd73074a52d1856e4da47fe8b26d802d44f1cb4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac2d2978d920ad644594db57606edef7018e018971a4d417f54446a2ce533b456aca610354322843990c2e2a43563b555aca46b1f43fd1f0502ff558252bfab3f268f01dcb87cdd2b186c8bf0cafccbf8a34dfa73936ec72eee06c30f0e0ae4ae6d14c59d6f30b37504b24f1210081eff2628eb45740234d8226e2199c7b6454;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc35ed77c928cb19fed312b000a5ae24f0eab5d2388da09cac767d3e4e5f9c0b26c344885bdfb10d97f6d8428432c64f2c52b64e22e6fb67499a08cf52569e646ea845d61ef5a509d2fac7faf2db63796618cabce3c9350a6b4181a0259d561efcaaa09d6764bf935fdf91d3dd4e5725234f6466be2404a5fe410c2449b44903f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19e8eba54e957b20e68d4fc069bd2dafc58e24b1008697f3b87e39d2a95f71fdd2bbc1982208affe03490f14e0acf6c1600902b75c1f919a0e29c3da3511f6eb0c901cd7e31aa3f0c6aa88e91feda745a3dcca05fff74549fc4a65a757780d10fe571a17f48631372eff9667e6d21b6611f16b325faa670366b197764c9bd463;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb234fe4ac602ede62626777574502506f5334a6799e47be7a5716194d39a1ee9ab5b13e4439fd74b55f29c85973c9980657871e6effae33b70c9aa8e784527fb9e0cfd57e86997fc60823944a3c03a54c05ff87db047a791f307ce93f5cf9fb261941aa8904014d3b75ae43f177b64fd568e247256dfe450c5dc509824bd680a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4944980c58acfdc9ea082a4f4cb7d48b06b318c8f2f6ed5584fc2aab9b506f2c12d4a66e10efc443566b17350b9af31a84b22c4955250b18a4304ba67d3df83e0cd0e2211e31733b8e4a3cf47bd3d8212fab8ef019c5d4f9d7adc8893e962023e4435c7c5f42fe0a7ce39e50c7b6563b2ce35e2936d3eb297a8fdf383016e686;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d3d7dbc6413182dcb0c5e07c7de5333a45c7074b4b3f9b8e3a5a1f2e35638e44cf08727cbab5f14f577ceba8bfcf1b2d82e42e998052b1c9b91fd749613eda74e4ee72d920ef41e0c714d4e960e724d2e16b024a6072983b2b13bee06eefc380b82af6bd3d25786b15fe96b8f24888c645e3e0c0718aea3f68afc4e6ebf05aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee8b0712825159e332d23b2415cd911648870f69847d1c1f28cc6142d43933f89475b5cd10b03d00793dd0ede66de6d1122af584e0efe14d099cbe52f55e3461643f653f1bcc74d132594ca040b0352d04f68f0f3e3492648617948b0ec6017ddf780e0da8eefa6e2dc82c64e4a84fabb4789a68154b6a337c55a71792c5c14a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d9fb40b1135743ea32d808296b379633c2fc86ac8ad9857d1cfed044d8b7f1a5f67168bf2a69d089ca354ba39c9530679a2adb517c744a49026a71bb399d1f56e02d91e258b1477c8d39231b3774c75099d818223358c7600aade11b471bf60dc8f227d7e1a348cda6a62bb492ef0d623701b6281ac84e56025eef198f7dceb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7486c7b5f739321a05440d3d031342d62501529070762750c9acc6a6b18f31a54ef49d2fd0eece957b041859c6508c6c6bad3c39a25834298c18e3e28121785d0b97007167bcf06c5e02f2aa8795073cb8bd88b0890b95b805d17e9f66320e91010ac9f0fd2af0d9e7e839ce76ec72455de9b7a315cb1ab93ebf1aa7eb8636c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c93c9a7685f23ab4bcc84e190a3168913632535c466d4adb41648a263ae896178780155b2f3a32b519b369c7fb842ef2e2bc4098f89a75abc1ce4715ac83d0db74233cdb1f8b6815874e233e382e493a06ae35c07e55ef01a40ef6cc13a59057b70b7e815f4bbb55d34261457c857131dbe6d1e58eb7678a0f0b69c3b4ce013;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc96dd3fd0c5f9a5bb09f4d72e417fd55f5c2dc9999bac7afd5c231b5351a25fbccb7ed7157c859ed07bbac846249a82e455e47d08fb5a0f25aaa26bac2cf6bfb8ce66712d54884e1303979d3a10e66426f19308e51bbbe75ca194ef1b766b3a262e4180a9d3b598bfc7f7fd33dbb1b60e62414a7254f5fdbbd5f4b4b5291d490;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87d2595919b6943f8a1f67a1988a2c44f36c0ddb795fd3f994b48f7290d69e8c268004662a755662a4345b8f8627b5562ce3a0fbecede0f559a78541f4c47dd35020efbc70f7512e8d4dd2bec65f8ca0feaa75f6ee2ffcae7074205ae8ce1340f5e0d8910188b6acf39736367414232cf237a2d03418dc931e30a30d4aa0f88a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3da6309657b1f309c9fd79fc584aa5ad7db11fad6c1fb48979eb38a2d23c0279992676632d9a9093f0bc264458ef265a6e94a6882b08d54026ef470462701db497c0bf81b7b9b8565a2b913aa6bd5c3eca9a801da5caef3e2088b9613a8f12d2b9ce95b1b286c1cb01d37d07fd56196e146e96ed6ab9764fae680f3f971e8fb2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49f84adafd4b58a06eb18b280a48987291c7701418bc79f129ddcb4a10499677f5c0b6421711e12f9a9285514930365a8ded8a459a24a5996947256e3870c54355f9b4e66ca5d147a609d3a1830b765a21640d9aab61339fd6d9c85c2fce0803458d3723ff695c0762286abbdfe832fcccf54257417b2740eb19766bb1f8ff6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab205ce9365525730dd651dd6159cf16301074e022252c59731e20f7fc46f980293852db1fb37ccb8622d204e6f9b9356897adcc21a628b5e16dcdb700510d6059473e449f7aafafac21a8469d6aa2e0910c145096f1bd18d4db8f36f1baaaf02bf5797e57009634ee2442e5d56c2f62887ef219827eb9d83ed4efe33d7562aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a563c75f54abb3e39ce6536832b6ae0318143a4de8bd2a907fb7187dc1bc8e77a5f67ccf361144ad66db185a1291a387353fc4c2b92332b0780c69ace34fd11db601ad53673b3ff5d38341de20503a465ce60d9121808cefc340e5003f7a33148216588640732256dee51bd224560333035ad3d31b213cc1fb056c4f2cf8b8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc548681fb089e3bdd6f8070d110b646d917fca08d935241e2f0ad344f74099cf74a1010f7cf04937b95f1daa1130d8004e9e7721044dee5374c9f14ab27172ce81061ede068eb9341f128882ea219d6d6f1a526fe7c34bdf99aa4beb0bce900f2d357daca81471423bb49850d9c4efb1876fc984b5543039a458f1c67e39b90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc321126879682318d9a8075c5a1d6bc135ad64df57ea53d066969d7ecf2536672a7098743206e9b768dce5ad0987b50a0b221955007cff079913ac7dcc48904d5030234eb4998f9dcd3df5c3a4c4bf710345fc1219fa1c9bce3d8d1353d7d908df7a6006a23720f90b1ba5ae7b0d40f64e168c514c4794e936501f080efab2ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd425e4924cc5a9b11b63c74e8314b2873ac1636197221c46ebc89af66b10db935394f962acebff7108d9598cd85ea293a9fbe5053287f14788e51753b679cd88ff4ecdbcc7264427b15a0a694bb822cd6fb35f0dbd2fbee3715e04cbf15f2d8f9dd6cabc8c64da5d3f2d9ff7ad285571e6e698f6809a446a63c64c4a63316aee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h514156a680e4de8d04cb40086797963403186130fffba95f436eb8057aa81fde499e1c9bc3872681097d2b3dc8f8c759ea2c3c33d037623e9139d4590b4063844bb10347f80caa1c615b93953e670aead56a3822a0e3f17065903991fdc1346f2fd9711230a35e01f6b198ddf33db551c8f7b0e15930a7a89c02183525e5813d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37bd990b331d3fa8cbba68c98e17287c946a88ab751e584459fdb33bc87ec83a470e6a5506c75a1e0278fbd90d346f09d8079e9a6d61858d8e5a9539c399fbf5026a548ef984cc8f82521e9eafdaac48dcc22c6e99514d69eb51595c83e41d92a2d3cbec9102e37ff57f13dead59f308381385b81c1faac22374e8cf527ec9e8;
        #1
        $finish();
    end
endmodule
