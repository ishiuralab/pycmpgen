module compressor2_1_32_12_shiftregister(input clk, input in_data0, input in_data1, input in_data2, input in_data3, input in_data4, input in_data5, input in_data6, input in_data7, input in_data8, input in_data9, input in_data10, input in_data11, input in_data12, input in_data13, input in_data14, input in_data15, input in_data16, input in_data17, input in_data18, input in_data19, input in_data20, input in_data21, input in_data22, input in_data23, input in_data24, input in_data25, input in_data26, input in_data27, input in_data28, input in_data29, input in_data30, input in_data31, output [16:0]dst);
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    compressor2_1_32_12 compressor2_1_32_12(.src0(src0), .src1(src1), .src2(src2), .src3(src3), .src4(src4), .src5(src5), .src6(src6), .src7(src7), .src8(src8), .src9(src9), .src10(src10), .src11(src11), .src12(src12), .src13(src13), .src14(src14), .src15(src15), .src16(src16), .src17(src17), .src18(src18), .src19(src19), .src20(src20), .src21(src21), .src22(src22), .src23(src23), .src24(src24), .src25(src25), .src26(src26), .src27(src27), .src28(src28), .src29(src29), .src30(src30), .src31(src31), .dst(dst));
    initial begin
        src0 <= 0;
        src1 <= 0;
        src2 <= 0;
        src3 <= 0;
        src4 <= 0;
        src5 <= 0;
        src6 <= 0;
        src7 <= 0;
        src8 <= 0;
        src9 <= 0;
        src10 <= 0;
        src11 <= 0;
        src12 <= 0;
        src13 <= 0;
        src14 <= 0;
        src15 <= 0;
        src16 <= 0;
        src17 <= 0;
        src18 <= 0;
        src19 <= 0;
        src20 <= 0;
        src21 <= 0;
        src22 <= 0;
        src23 <= 0;
        src24 <= 0;
        src25 <= 0;
        src26 <= 0;
        src27 <= 0;
        src28 <= 0;
        src29 <= 0;
        src30 <= 0;
        src31 <= 0;
    end
    always @(posedge clk) begin
        src0 <= {src0[10:0], in_data0};
        src1 <= {src1[10:0], in_data1};
        src2 <= {src2[10:0], in_data2};
        src3 <= {src3[10:0], in_data3};
        src4 <= {src4[10:0], in_data4};
        src5 <= {src5[10:0], in_data5};
        src6 <= {src6[10:0], in_data6};
        src7 <= {src7[10:0], in_data7};
        src8 <= {src8[10:0], in_data8};
        src9 <= {src9[10:0], in_data9};
        src10 <= {src10[10:0], in_data10};
        src11 <= {src11[10:0], in_data11};
        src12 <= {src12[10:0], in_data12};
        src13 <= {src13[10:0], in_data13};
        src14 <= {src14[10:0], in_data14};
        src15 <= {src15[10:0], in_data15};
        src16 <= {src16[10:0], in_data16};
        src17 <= {src17[10:0], in_data17};
        src18 <= {src18[10:0], in_data18};
        src19 <= {src19[10:0], in_data19};
        src20 <= {src20[10:0], in_data20};
        src21 <= {src21[10:0], in_data21};
        src22 <= {src22[10:0], in_data22};
        src23 <= {src23[10:0], in_data23};
        src24 <= {src24[10:0], in_data24};
        src25 <= {src25[10:0], in_data25};
        src26 <= {src26[10:0], in_data26};
        src27 <= {src27[10:0], in_data27};
        src28 <= {src28[10:0], in_data28};
        src29 <= {src29[10:0], in_data29};
        src30 <= {src30[10:0], in_data30};
        src31 <= {src31[10:0], in_data31};
    end
endmodule

module compressor2_1_32_12(
    input [11:0]src0,
    input [11:0]src1,
    input [11:0]src2,
    input [11:0]src3,
    input [11:0]src4,
    input [11:0]src5,
    input [11:0]src6,
    input [11:0]src7,
    input [11:0]src8,
    input [11:0]src9,
    input [11:0]src10,
    input [11:0]src11,
    input [11:0]src12,
    input [11:0]src13,
    input [11:0]src14,
    input [11:0]src15,
    input [11:0]src16,
    input [11:0]src17,
    input [11:0]src18,
    input [11:0]src19,
    input [11:0]src20,
    input [11:0]src21,
    input [11:0]src22,
    input [11:0]src23,
    input [11:0]src24,
    input [11:0]src25,
    input [11:0]src26,
    input [11:0]src27,
    input [11:0]src28,
    input [11:0]src29,
    input [11:0]src30,
    input [11:0]src31,
    output [16:0]dst);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [0:0] comp_out15;
    wire [0:0] comp_out16;
    wire [17:0] out;
    compressor compressor_inst(
        .src0({src31[0], src30[0], src29[0], src28[0], src27[0], src26[0], src25[0], src24[0], src23[0], src22[0], src21[0], src20[0], src19[0], src18[0], src17[0], src16[0], src15[0], src14[0], src13[0], src12[0], src11[0], src10[0], src9[0], src8[0], src7[0], src6[0], src5[0], src4[0], src3[0], src2[0], src1[0], src0[0]}),
        .src1({src31[1], src30[1], src29[1], src28[1], src27[1], src26[1], src25[1], src24[1], src23[1], src22[1], src21[1], src20[1], src19[1], src18[1], src17[1], src16[1], src15[1], src14[1], src13[1], src12[1], src11[1], src10[1], src9[1], src8[1], src7[1], src6[1], src5[1], src4[1], src3[1], src2[1], src1[1], src0[1]}),
        .src2({src31[2], src30[2], src29[2], src28[2], src27[2], src26[2], src25[2], src24[2], src23[2], src22[2], src21[2], src20[2], src19[2], src18[2], src17[2], src16[2], src15[2], src14[2], src13[2], src12[2], src11[2], src10[2], src9[2], src8[2], src7[2], src6[2], src5[2], src4[2], src3[2], src2[2], src1[2], src0[2]}),
        .src3({src31[3], src30[3], src29[3], src28[3], src27[3], src26[3], src25[3], src24[3], src23[3], src22[3], src21[3], src20[3], src19[3], src18[3], src17[3], src16[3], src15[3], src14[3], src13[3], src12[3], src11[3], src10[3], src9[3], src8[3], src7[3], src6[3], src5[3], src4[3], src3[3], src2[3], src1[3], src0[3]}),
        .src4({src31[4], src30[4], src29[4], src28[4], src27[4], src26[4], src25[4], src24[4], src23[4], src22[4], src21[4], src20[4], src19[4], src18[4], src17[4], src16[4], src15[4], src14[4], src13[4], src12[4], src11[4], src10[4], src9[4], src8[4], src7[4], src6[4], src5[4], src4[4], src3[4], src2[4], src1[4], src0[4]}),
        .src5({src31[5], src30[5], src29[5], src28[5], src27[5], src26[5], src25[5], src24[5], src23[5], src22[5], src21[5], src20[5], src19[5], src18[5], src17[5], src16[5], src15[5], src14[5], src13[5], src12[5], src11[5], src10[5], src9[5], src8[5], src7[5], src6[5], src5[5], src4[5], src3[5], src2[5], src1[5], src0[5]}),
        .src6({src31[6], src30[6], src29[6], src28[6], src27[6], src26[6], src25[6], src24[6], src23[6], src22[6], src21[6], src20[6], src19[6], src18[6], src17[6], src16[6], src15[6], src14[6], src13[6], src12[6], src11[6], src10[6], src9[6], src8[6], src7[6], src6[6], src5[6], src4[6], src3[6], src2[6], src1[6], src0[6]}),
        .src7({src31[7], src30[7], src29[7], src28[7], src27[7], src26[7], src25[7], src24[7], src23[7], src22[7], src21[7], src20[7], src19[7], src18[7], src17[7], src16[7], src15[7], src14[7], src13[7], src12[7], src11[7], src10[7], src9[7], src8[7], src7[7], src6[7], src5[7], src4[7], src3[7], src2[7], src1[7], src0[7]}),
        .src8({src31[8], src30[8], src29[8], src28[8], src27[8], src26[8], src25[8], src24[8], src23[8], src22[8], src21[8], src20[8], src19[8], src18[8], src17[8], src16[8], src15[8], src14[8], src13[8], src12[8], src11[8], src10[8], src9[8], src8[8], src7[8], src6[8], src5[8], src4[8], src3[8], src2[8], src1[8], src0[8]}),
        .src9({src31[9], src30[9], src29[9], src28[9], src27[9], src26[9], src25[9], src24[9], src23[9], src22[9], src21[9], src20[9], src19[9], src18[9], src17[9], src16[9], src15[9], src14[9], src13[9], src12[9], src11[9], src10[9], src9[9], src8[9], src7[9], src6[9], src5[9], src4[9], src3[9], src2[9], src1[9], src0[9]}),
        .src10({src31[10], src30[10], src29[10], src28[10], src27[10], src26[10], src25[10], src24[10], src23[10], src22[10], src21[10], src20[10], src19[10], src18[10], src17[10], src16[10], src15[10], src14[10], src13[10], src12[10], src11[10], src10[10], src9[10], src8[10], src7[10], src6[10], src5[10], src4[10], src3[10], src2[10], src1[10], src0[10]}),
        .src11({src31[11], src30[11], src29[11], src28[11], src27[11], src26[11], src25[11], src24[11], src23[11], src22[11], src21[11], src20[11], src19[11], src18[11], src17[11], src16[11], src15[11], src14[11], src13[11], src12[11], src11[11], src10[11], src9[11], src8[11], src7[11], src6[11], src5[11], src4[11], src3[11], src2[11], src1[11], src0[11]}),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16)
    );
    rowadder2_1_17 rowadder2_1inst(
        .src0({comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst0(out)
    );
    assign dst = out[16:0];
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [0:0] dst15,
      output wire [0:0] dst16);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [17:0] stage1_0;
   wire [8:0] stage1_1;
   wire [11:0] stage1_2;
   wire [11:0] stage1_3;
   wire [13:0] stage1_4;
   wire [14:0] stage1_5;
   wire [16:0] stage1_6;
   wire [10:0] stage1_7;
   wire [21:0] stage1_8;
   wire [28:0] stage1_9;
   wire [24:0] stage1_10;
   wire [29:0] stage1_11;
   wire [2:0] stage1_12;
   wire [0:0] stage1_13;
   wire [7:0] stage2_0;
   wire [10:0] stage2_1;
   wire [1:0] stage2_2;
   wire [5:0] stage2_3;
   wire [6:0] stage2_4;
   wire [3:0] stage2_5;
   wire [5:0] stage2_6;
   wire [12:0] stage2_7;
   wire [5:0] stage2_8;
   wire [12:0] stage2_9;
   wire [11:0] stage2_10;
   wire [11:0] stage2_11;
   wire [8:0] stage2_12;
   wire [5:0] stage2_13;
   wire [7:0] stage3_0;
   wire [5:0] stage3_1;
   wire [2:0] stage3_2;
   wire [0:0] stage3_3;
   wire [2:0] stage3_4;
   wire [5:0] stage3_5;
   wire [0:0] stage3_6;
   wire [8:0] stage3_7;
   wire [3:0] stage3_8;
   wire [2:0] stage3_9;
   wire [3:0] stage3_10;
   wire [5:0] stage3_11;
   wire [5:0] stage3_12;
   wire [2:0] stage3_13;
   wire [1:0] stage3_14;
   wire [0:0] stage3_15;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [0:0] stage4_15;
   wire [0:0] stage4_16;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;

   gpc606_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_2[0], stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc615_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[0]},
      {stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc606_5 gpc3 (
      {stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3]}
   );
   gpc606_5 gpc4 (
      {stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12]},
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11]},
      {stage1_5[1],stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4]}
   );
   gpc606_5 gpc5 (
      {stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18]},
      {stage0_3[12], stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17]},
      {stage1_5[2],stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[3],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[4],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc606_5 gpc8 (
      {stage0_2[18], stage0_2[19], stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[5],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc606_5 gpc9 (
      {stage0_2[24], stage0_2[25], stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[6],stage1_4[9],stage1_3[9],stage1_2[9]}
   );
   gpc2135_5 gpc10 (
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16]},
      {stage0_5[0], stage0_5[1], stage0_5[2]},
      {stage0_6[0]},
      {stage0_7[0], stage0_7[1]},
      {stage1_8[0],stage1_7[0],stage1_6[2],stage1_5[7],stage1_4[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_6[1]},
      {stage0_7[2]},
      {stage1_8[1],stage1_7[1],stage1_6[3],stage1_5[8],stage1_4[11]}
   );
   gpc606_5 gpc12 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25]},
      {stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7]},
      {stage1_8[2],stage1_7[2],stage1_6[4],stage1_5[9],stage1_4[12]}
   );
   gpc606_5 gpc13 (
      {stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31]},
      {stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11], stage0_6[12], stage0_6[13]},
      {stage1_8[3],stage1_7[3],stage1_6[5],stage1_5[10],stage1_4[13]}
   );
   gpc606_5 gpc14 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6], stage0_7[7], stage0_7[8]},
      {stage1_9[0],stage1_8[4],stage1_7[4],stage1_6[6],stage1_5[11]}
   );
   gpc606_5 gpc15 (
      {stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20]},
      {stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12], stage0_7[13], stage0_7[14]},
      {stage1_9[1],stage1_8[5],stage1_7[5],stage1_6[7],stage1_5[12]}
   );
   gpc606_5 gpc16 (
      {stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26]},
      {stage0_7[15], stage0_7[16], stage0_7[17], stage0_7[18], stage0_7[19], stage0_7[20]},
      {stage1_9[2],stage1_8[6],stage1_7[6],stage1_6[8],stage1_5[13]}
   );
   gpc615_5 gpc17 (
      {stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage0_6[14]},
      {stage0_7[21], stage0_7[22], stage0_7[23], stage0_7[24], stage0_7[25], stage0_7[26]},
      {stage1_9[3],stage1_8[7],stage1_7[7],stage1_6[9],stage1_5[14]}
   );
   gpc606_5 gpc18 (
      {stage0_6[15], stage0_6[16], stage0_6[17], stage0_6[18], stage0_6[19], stage0_6[20]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[8],stage1_7[8],stage1_6[10]}
   );
   gpc606_5 gpc19 (
      {stage0_6[21], stage0_6[22], stage0_6[23], stage0_6[24], stage0_6[25], stage0_6[26]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[5],stage1_8[9],stage1_7[9],stage1_6[11]}
   );
   gpc615_5 gpc20 (
      {stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30], stage0_7[31]},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[6],stage1_8[10],stage1_7[10]}
   );
   gpc615_5 gpc21 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage0_9[6]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[1],stage1_10[3],stage1_9[7],stage1_8[11]}
   );
   gpc615_5 gpc22 (
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22]},
      {stage0_9[7]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[2],stage1_10[4],stage1_9[8],stage1_8[12]}
   );
   gpc615_5 gpc23 (
      {stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11], stage0_9[12]},
      {stage0_10[12]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[2],stage1_11[3],stage1_10[5],stage1_9[9]}
   );
   gpc1_1 gpc24 (
      {stage0_0[17]},
      {stage1_0[3]}
   );
   gpc1_1 gpc25 (
      {stage0_0[18]},
      {stage1_0[4]}
   );
   gpc1_1 gpc26 (
      {stage0_0[19]},
      {stage1_0[5]}
   );
   gpc1_1 gpc27 (
      {stage0_0[20]},
      {stage1_0[6]}
   );
   gpc1_1 gpc28 (
      {stage0_0[21]},
      {stage1_0[7]}
   );
   gpc1_1 gpc29 (
      {stage0_0[22]},
      {stage1_0[8]}
   );
   gpc1_1 gpc30 (
      {stage0_0[23]},
      {stage1_0[9]}
   );
   gpc1_1 gpc31 (
      {stage0_0[24]},
      {stage1_0[10]}
   );
   gpc1_1 gpc32 (
      {stage0_0[25]},
      {stage1_0[11]}
   );
   gpc1_1 gpc33 (
      {stage0_0[26]},
      {stage1_0[12]}
   );
   gpc1_1 gpc34 (
      {stage0_0[27]},
      {stage1_0[13]}
   );
   gpc1_1 gpc35 (
      {stage0_0[28]},
      {stage1_0[14]}
   );
   gpc1_1 gpc36 (
      {stage0_0[29]},
      {stage1_0[15]}
   );
   gpc1_1 gpc37 (
      {stage0_0[30]},
      {stage1_0[16]}
   );
   gpc1_1 gpc38 (
      {stage0_0[31]},
      {stage1_0[17]}
   );
   gpc1_1 gpc39 (
      {stage0_1[31]},
      {stage1_1[8]}
   );
   gpc1_1 gpc40 (
      {stage0_2[30]},
      {stage1_2[10]}
   );
   gpc1_1 gpc41 (
      {stage0_2[31]},
      {stage1_2[11]}
   );
   gpc1_1 gpc42 (
      {stage0_3[30]},
      {stage1_3[10]}
   );
   gpc1_1 gpc43 (
      {stage0_3[31]},
      {stage1_3[11]}
   );
   gpc1_1 gpc44 (
      {stage0_6[27]},
      {stage1_6[12]}
   );
   gpc1_1 gpc45 (
      {stage0_6[28]},
      {stage1_6[13]}
   );
   gpc1_1 gpc46 (
      {stage0_6[29]},
      {stage1_6[14]}
   );
   gpc1_1 gpc47 (
      {stage0_6[30]},
      {stage1_6[15]}
   );
   gpc1_1 gpc48 (
      {stage0_6[31]},
      {stage1_6[16]}
   );
   gpc1_1 gpc49 (
      {stage0_8[23]},
      {stage1_8[13]}
   );
   gpc1_1 gpc50 (
      {stage0_8[24]},
      {stage1_8[14]}
   );
   gpc1_1 gpc51 (
      {stage0_8[25]},
      {stage1_8[15]}
   );
   gpc1_1 gpc52 (
      {stage0_8[26]},
      {stage1_8[16]}
   );
   gpc1_1 gpc53 (
      {stage0_8[27]},
      {stage1_8[17]}
   );
   gpc1_1 gpc54 (
      {stage0_8[28]},
      {stage1_8[18]}
   );
   gpc1_1 gpc55 (
      {stage0_8[29]},
      {stage1_8[19]}
   );
   gpc1_1 gpc56 (
      {stage0_8[30]},
      {stage1_8[20]}
   );
   gpc1_1 gpc57 (
      {stage0_8[31]},
      {stage1_8[21]}
   );
   gpc1_1 gpc58 (
      {stage0_9[13]},
      {stage1_9[10]}
   );
   gpc1_1 gpc59 (
      {stage0_9[14]},
      {stage1_9[11]}
   );
   gpc1_1 gpc60 (
      {stage0_9[15]},
      {stage1_9[12]}
   );
   gpc1_1 gpc61 (
      {stage0_9[16]},
      {stage1_9[13]}
   );
   gpc1_1 gpc62 (
      {stage0_9[17]},
      {stage1_9[14]}
   );
   gpc1_1 gpc63 (
      {stage0_9[18]},
      {stage1_9[15]}
   );
   gpc1_1 gpc64 (
      {stage0_9[19]},
      {stage1_9[16]}
   );
   gpc1_1 gpc65 (
      {stage0_9[20]},
      {stage1_9[17]}
   );
   gpc1_1 gpc66 (
      {stage0_9[21]},
      {stage1_9[18]}
   );
   gpc1_1 gpc67 (
      {stage0_9[22]},
      {stage1_9[19]}
   );
   gpc1_1 gpc68 (
      {stage0_9[23]},
      {stage1_9[20]}
   );
   gpc1_1 gpc69 (
      {stage0_9[24]},
      {stage1_9[21]}
   );
   gpc1_1 gpc70 (
      {stage0_9[25]},
      {stage1_9[22]}
   );
   gpc1_1 gpc71 (
      {stage0_9[26]},
      {stage1_9[23]}
   );
   gpc1_1 gpc72 (
      {stage0_9[27]},
      {stage1_9[24]}
   );
   gpc1_1 gpc73 (
      {stage0_9[28]},
      {stage1_9[25]}
   );
   gpc1_1 gpc74 (
      {stage0_9[29]},
      {stage1_9[26]}
   );
   gpc1_1 gpc75 (
      {stage0_9[30]},
      {stage1_9[27]}
   );
   gpc1_1 gpc76 (
      {stage0_9[31]},
      {stage1_9[28]}
   );
   gpc1_1 gpc77 (
      {stage0_10[13]},
      {stage1_10[6]}
   );
   gpc1_1 gpc78 (
      {stage0_10[14]},
      {stage1_10[7]}
   );
   gpc1_1 gpc79 (
      {stage0_10[15]},
      {stage1_10[8]}
   );
   gpc1_1 gpc80 (
      {stage0_10[16]},
      {stage1_10[9]}
   );
   gpc1_1 gpc81 (
      {stage0_10[17]},
      {stage1_10[10]}
   );
   gpc1_1 gpc82 (
      {stage0_10[18]},
      {stage1_10[11]}
   );
   gpc1_1 gpc83 (
      {stage0_10[19]},
      {stage1_10[12]}
   );
   gpc1_1 gpc84 (
      {stage0_10[20]},
      {stage1_10[13]}
   );
   gpc1_1 gpc85 (
      {stage0_10[21]},
      {stage1_10[14]}
   );
   gpc1_1 gpc86 (
      {stage0_10[22]},
      {stage1_10[15]}
   );
   gpc1_1 gpc87 (
      {stage0_10[23]},
      {stage1_10[16]}
   );
   gpc1_1 gpc88 (
      {stage0_10[24]},
      {stage1_10[17]}
   );
   gpc1_1 gpc89 (
      {stage0_10[25]},
      {stage1_10[18]}
   );
   gpc1_1 gpc90 (
      {stage0_10[26]},
      {stage1_10[19]}
   );
   gpc1_1 gpc91 (
      {stage0_10[27]},
      {stage1_10[20]}
   );
   gpc1_1 gpc92 (
      {stage0_10[28]},
      {stage1_10[21]}
   );
   gpc1_1 gpc93 (
      {stage0_10[29]},
      {stage1_10[22]}
   );
   gpc1_1 gpc94 (
      {stage0_10[30]},
      {stage1_10[23]}
   );
   gpc1_1 gpc95 (
      {stage0_10[31]},
      {stage1_10[24]}
   );
   gpc1_1 gpc96 (
      {stage0_11[6]},
      {stage1_11[4]}
   );
   gpc1_1 gpc97 (
      {stage0_11[7]},
      {stage1_11[5]}
   );
   gpc1_1 gpc98 (
      {stage0_11[8]},
      {stage1_11[6]}
   );
   gpc1_1 gpc99 (
      {stage0_11[9]},
      {stage1_11[7]}
   );
   gpc1_1 gpc100 (
      {stage0_11[10]},
      {stage1_11[8]}
   );
   gpc1_1 gpc101 (
      {stage0_11[11]},
      {stage1_11[9]}
   );
   gpc1_1 gpc102 (
      {stage0_11[12]},
      {stage1_11[10]}
   );
   gpc1_1 gpc103 (
      {stage0_11[13]},
      {stage1_11[11]}
   );
   gpc1_1 gpc104 (
      {stage0_11[14]},
      {stage1_11[12]}
   );
   gpc1_1 gpc105 (
      {stage0_11[15]},
      {stage1_11[13]}
   );
   gpc1_1 gpc106 (
      {stage0_11[16]},
      {stage1_11[14]}
   );
   gpc1_1 gpc107 (
      {stage0_11[17]},
      {stage1_11[15]}
   );
   gpc1_1 gpc108 (
      {stage0_11[18]},
      {stage1_11[16]}
   );
   gpc1_1 gpc109 (
      {stage0_11[19]},
      {stage1_11[17]}
   );
   gpc1_1 gpc110 (
      {stage0_11[20]},
      {stage1_11[18]}
   );
   gpc1_1 gpc111 (
      {stage0_11[21]},
      {stage1_11[19]}
   );
   gpc1_1 gpc112 (
      {stage0_11[22]},
      {stage1_11[20]}
   );
   gpc1_1 gpc113 (
      {stage0_11[23]},
      {stage1_11[21]}
   );
   gpc1_1 gpc114 (
      {stage0_11[24]},
      {stage1_11[22]}
   );
   gpc1_1 gpc115 (
      {stage0_11[25]},
      {stage1_11[23]}
   );
   gpc1_1 gpc116 (
      {stage0_11[26]},
      {stage1_11[24]}
   );
   gpc1_1 gpc117 (
      {stage0_11[27]},
      {stage1_11[25]}
   );
   gpc1_1 gpc118 (
      {stage0_11[28]},
      {stage1_11[26]}
   );
   gpc1_1 gpc119 (
      {stage0_11[29]},
      {stage1_11[27]}
   );
   gpc1_1 gpc120 (
      {stage0_11[30]},
      {stage1_11[28]}
   );
   gpc1_1 gpc121 (
      {stage0_11[31]},
      {stage1_11[29]}
   );
   gpc606_5 gpc122 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc123 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc124 (
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4]},
      {stage1_4[0]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[0],stage2_4[2],stage2_3[2]}
   );
   gpc615_5 gpc125 (
      {stage1_3[5], stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9]},
      {stage1_4[1]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[1],stage2_4[3],stage2_3[3]}
   );
   gpc2135_5 gpc126 (
      {stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5], stage1_4[6]},
      {stage1_5[12], stage1_5[13], stage1_5[14]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[0],stage2_7[2],stage2_6[2],stage2_5[2],stage2_4[4]}
   );
   gpc606_5 gpc127 (
      {stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11], stage1_4[12]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[1],stage2_7[3],stage2_6[3],stage2_5[3],stage2_4[5]}
   );
   gpc615_5 gpc128 (
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_7[2]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[2],stage2_7[4],stage2_6[4]}
   );
   gpc615_5 gpc129 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16]},
      {stage1_7[3]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[3],stage2_7[5],stage2_6[5]}
   );
   gpc615_5 gpc130 (
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16]},
      {stage1_9[0]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[0],stage2_10[2],stage2_9[2],stage2_8[4]}
   );
   gpc615_5 gpc131 (
      {stage1_8[17], stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21]},
      {stage1_9[1]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[1],stage2_10[3],stage2_9[3],stage2_8[5]}
   );
   gpc1163_5 gpc132 (
      {stage1_9[2], stage1_9[3], stage1_9[4]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_11[0]},
      {stage1_12[0]},
      {stage2_13[0],stage2_12[2],stage2_11[2],stage2_10[4],stage2_9[4]}
   );
   gpc615_5 gpc133 (
      {stage1_9[5], stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9]},
      {stage1_10[18]},
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5], stage1_11[6]},
      {stage2_13[1],stage2_12[3],stage2_11[3],stage2_10[5],stage2_9[5]}
   );
   gpc615_5 gpc134 (
      {stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13], stage1_9[14]},
      {stage1_10[19]},
      {stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11], stage1_11[12]},
      {stage2_13[2],stage2_12[4],stage2_11[4],stage2_10[6],stage2_9[6]}
   );
   gpc615_5 gpc135 (
      {stage1_9[15], stage1_9[16], stage1_9[17], stage1_9[18], stage1_9[19]},
      {stage1_10[20]},
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage2_13[3],stage2_12[5],stage2_11[5],stage2_10[7],stage2_9[7]}
   );
   gpc615_5 gpc136 (
      {stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24]},
      {stage1_10[21]},
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage2_13[4],stage2_12[6],stage2_11[6],stage2_10[8],stage2_9[8]}
   );
   gpc1_1 gpc137 (
      {stage1_0[12]},
      {stage2_0[2]}
   );
   gpc1_1 gpc138 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc139 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc140 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc141 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc142 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc143 (
      {stage1_1[0]},
      {stage2_1[2]}
   );
   gpc1_1 gpc144 (
      {stage1_1[1]},
      {stage2_1[3]}
   );
   gpc1_1 gpc145 (
      {stage1_1[2]},
      {stage2_1[4]}
   );
   gpc1_1 gpc146 (
      {stage1_1[3]},
      {stage2_1[5]}
   );
   gpc1_1 gpc147 (
      {stage1_1[4]},
      {stage2_1[6]}
   );
   gpc1_1 gpc148 (
      {stage1_1[5]},
      {stage2_1[7]}
   );
   gpc1_1 gpc149 (
      {stage1_1[6]},
      {stage2_1[8]}
   );
   gpc1_1 gpc150 (
      {stage1_1[7]},
      {stage2_1[9]}
   );
   gpc1_1 gpc151 (
      {stage1_1[8]},
      {stage2_1[10]}
   );
   gpc1_1 gpc152 (
      {stage1_3[10]},
      {stage2_3[4]}
   );
   gpc1_1 gpc153 (
      {stage1_3[11]},
      {stage2_3[5]}
   );
   gpc1_1 gpc154 (
      {stage1_4[13]},
      {stage2_4[6]}
   );
   gpc1_1 gpc155 (
      {stage1_7[4]},
      {stage2_7[6]}
   );
   gpc1_1 gpc156 (
      {stage1_7[5]},
      {stage2_7[7]}
   );
   gpc1_1 gpc157 (
      {stage1_7[6]},
      {stage2_7[8]}
   );
   gpc1_1 gpc158 (
      {stage1_7[7]},
      {stage2_7[9]}
   );
   gpc1_1 gpc159 (
      {stage1_7[8]},
      {stage2_7[10]}
   );
   gpc1_1 gpc160 (
      {stage1_7[9]},
      {stage2_7[11]}
   );
   gpc1_1 gpc161 (
      {stage1_7[10]},
      {stage2_7[12]}
   );
   gpc1_1 gpc162 (
      {stage1_9[25]},
      {stage2_9[9]}
   );
   gpc1_1 gpc163 (
      {stage1_9[26]},
      {stage2_9[10]}
   );
   gpc1_1 gpc164 (
      {stage1_9[27]},
      {stage2_9[11]}
   );
   gpc1_1 gpc165 (
      {stage1_9[28]},
      {stage2_9[12]}
   );
   gpc1_1 gpc166 (
      {stage1_10[22]},
      {stage2_10[9]}
   );
   gpc1_1 gpc167 (
      {stage1_10[23]},
      {stage2_10[10]}
   );
   gpc1_1 gpc168 (
      {stage1_10[24]},
      {stage2_10[11]}
   );
   gpc1_1 gpc169 (
      {stage1_11[25]},
      {stage2_11[7]}
   );
   gpc1_1 gpc170 (
      {stage1_11[26]},
      {stage2_11[8]}
   );
   gpc1_1 gpc171 (
      {stage1_11[27]},
      {stage2_11[9]}
   );
   gpc1_1 gpc172 (
      {stage1_11[28]},
      {stage2_11[10]}
   );
   gpc1_1 gpc173 (
      {stage1_11[29]},
      {stage2_11[11]}
   );
   gpc1_1 gpc174 (
      {stage1_12[1]},
      {stage2_12[7]}
   );
   gpc1_1 gpc175 (
      {stage1_12[2]},
      {stage2_12[8]}
   );
   gpc1_1 gpc176 (
      {stage1_13[0]},
      {stage2_13[5]}
   );
   gpc606_5 gpc177 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc606_5 gpc178 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1]}
   );
   gpc606_5 gpc179 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1],stage3_7[1]}
   );
   gpc615_5 gpc180 (
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4]},
      {stage2_9[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc181 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[1],stage3_11[2],stage3_10[2],stage3_9[2]}
   );
   gpc606_5 gpc182 (
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[2],stage3_11[3],stage3_10[3]}
   );
   gpc615_5 gpc183 (
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10]},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[2],stage3_12[3],stage3_11[4]}
   );
   gpc1_1 gpc184 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc185 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc186 (
      {stage2_0[2]},
      {stage3_0[2]}
   );
   gpc1_1 gpc187 (
      {stage2_0[3]},
      {stage3_0[3]}
   );
   gpc1_1 gpc188 (
      {stage2_0[4]},
      {stage3_0[4]}
   );
   gpc1_1 gpc189 (
      {stage2_0[5]},
      {stage3_0[5]}
   );
   gpc1_1 gpc190 (
      {stage2_0[6]},
      {stage3_0[6]}
   );
   gpc1_1 gpc191 (
      {stage2_0[7]},
      {stage3_0[7]}
   );
   gpc1_1 gpc192 (
      {stage2_1[6]},
      {stage3_1[1]}
   );
   gpc1_1 gpc193 (
      {stage2_1[7]},
      {stage3_1[2]}
   );
   gpc1_1 gpc194 (
      {stage2_1[8]},
      {stage3_1[3]}
   );
   gpc1_1 gpc195 (
      {stage2_1[9]},
      {stage3_1[4]}
   );
   gpc1_1 gpc196 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc197 (
      {stage2_2[0]},
      {stage3_2[1]}
   );
   gpc1_1 gpc198 (
      {stage2_2[1]},
      {stage3_2[2]}
   );
   gpc1_1 gpc199 (
      {stage2_4[6]},
      {stage3_4[2]}
   );
   gpc1_1 gpc200 (
      {stage2_5[0]},
      {stage3_5[2]}
   );
   gpc1_1 gpc201 (
      {stage2_5[1]},
      {stage3_5[3]}
   );
   gpc1_1 gpc202 (
      {stage2_5[2]},
      {stage3_5[4]}
   );
   gpc1_1 gpc203 (
      {stage2_5[3]},
      {stage3_5[5]}
   );
   gpc1_1 gpc204 (
      {stage2_7[6]},
      {stage3_7[2]}
   );
   gpc1_1 gpc205 (
      {stage2_7[7]},
      {stage3_7[3]}
   );
   gpc1_1 gpc206 (
      {stage2_7[8]},
      {stage3_7[4]}
   );
   gpc1_1 gpc207 (
      {stage2_7[9]},
      {stage3_7[5]}
   );
   gpc1_1 gpc208 (
      {stage2_7[10]},
      {stage3_7[6]}
   );
   gpc1_1 gpc209 (
      {stage2_7[11]},
      {stage3_7[7]}
   );
   gpc1_1 gpc210 (
      {stage2_7[12]},
      {stage3_7[8]}
   );
   gpc1_1 gpc211 (
      {stage2_8[5]},
      {stage3_8[3]}
   );
   gpc1_1 gpc212 (
      {stage2_11[11]},
      {stage3_11[5]}
   );
   gpc1_1 gpc213 (
      {stage2_12[7]},
      {stage3_12[4]}
   );
   gpc1_1 gpc214 (
      {stage2_12[8]},
      {stage3_12[5]}
   );
   gpc207_4 gpc215 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5], stage3_0[6]},
      {stage3_2[0], stage3_2[1]},
      {stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc2116_5 gpc216 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_2[2]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1]},
      {stage4_5[0],stage4_4[0],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc606_5 gpc217 (
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[0],stage4_7[0],stage4_6[0],stage4_5[1]}
   );
   gpc1343_5 gpc218 (
      {stage3_7[6], stage3_7[7], stage3_7[8]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3]},
      {stage3_9[0], stage3_9[1], stage3_9[2]},
      {stage3_10[0]},
      {stage4_11[0],stage4_10[0],stage4_9[1],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc219 (
      {stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[0]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[0],stage4_11[1],stage4_10[1]}
   );
   gpc1325_5 gpc220 (
      {stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage3_13[1], stage3_13[2]},
      {stage3_14[0], stage3_14[1], 1'b0},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1],stage4_12[1]}
   );
   gpc1_1 gpc221 (
      {stage3_0[7]},
      {stage4_0[1]}
   );
   gpc1_1 gpc222 (
      {stage3_4[2]},
      {stage4_4[1]}
   );
   gpc1_1 gpc223 (
      {stage3_6[0]},
      {stage4_6[1]}
   );
endmodule
module rowadder2_1_17(input [16:0] src0, input [16:0] src1, output [17:0] dst0);
    wire [16:0] gene;
    wire [16:0] prop;
    wire [19:0] out;
    wire [19:0] carryout;
    LUT2 #(
        .INIT(4'h8)
    ) lut_0_gene (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(gene[0])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_0_prop (
        .I0(src0[0]),
        .I1(src1[0]),
        .O(prop[0])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_1_gene (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(gene[1])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_1_prop (
        .I0(src0[1]),
        .I1(src1[1]),
        .O(prop[1])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_2_gene (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(gene[2])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_2_prop (
        .I0(src0[2]),
        .I1(src1[2]),
        .O(prop[2])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_3_gene (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(gene[3])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_3_prop (
        .I0(src0[3]),
        .I1(src1[3]),
        .O(prop[3])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_4_gene (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(gene[4])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_4_prop (
        .I0(src0[4]),
        .I1(src1[4]),
        .O(prop[4])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_5_gene (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(gene[5])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_5_prop (
        .I0(src0[5]),
        .I1(src1[5]),
        .O(prop[5])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_6_gene (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(gene[6])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_6_prop (
        .I0(src0[6]),
        .I1(src1[6]),
        .O(prop[6])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_7_gene (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(gene[7])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_7_prop (
        .I0(src0[7]),
        .I1(src1[7]),
        .O(prop[7])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_8_gene (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(gene[8])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_8_prop (
        .I0(src0[8]),
        .I1(src1[8]),
        .O(prop[8])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_9_gene (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(gene[9])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_9_prop (
        .I0(src0[9]),
        .I1(src1[9]),
        .O(prop[9])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_10_gene (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(gene[10])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_10_prop (
        .I0(src0[10]),
        .I1(src1[10]),
        .O(prop[10])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_11_gene (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(gene[11])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_11_prop (
        .I0(src0[11]),
        .I1(src1[11]),
        .O(prop[11])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_12_gene (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(gene[12])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_12_prop (
        .I0(src0[12]),
        .I1(src1[12]),
        .O(prop[12])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_13_gene (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(gene[13])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_13_prop (
        .I0(src0[13]),
        .I1(src1[13]),
        .O(prop[13])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_14_gene (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(gene[14])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_14_prop (
        .I0(src0[14]),
        .I1(src1[14]),
        .O(prop[14])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_15_gene (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(gene[15])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_15_prop (
        .I0(src0[15]),
        .I1(src1[15]),
        .O(prop[15])
    );
    LUT2 #(
        .INIT(4'h8)
    ) lut_16_gene (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(gene[16])
    );
    LUT2 #(
        .INIT(4'h6)
    ) lut_16_prop (
        .I0(src0[16]),
        .I1(src1[16]),
        .O(prop[16])
    );
    CARRY4 carry4_3_0 (
        .CO(carryout[3:0]),
        .O(out[3:0]),
        .CI(1'h0),
        .CYINIT(1'h0),
        .DI(gene[3:0]),
        .S(prop[3:0])
    );
    CARRY4 carry4_7_4 (
        .CO(carryout[7:4]),
        .O(out[7:4]),
        .CI(carryout[3]),
        .CYINIT(1'h0),
        .DI(gene[7:4]),
        .S(prop[7:4])
    );
    CARRY4 carry4_11_8 (
        .CO(carryout[11:8]),
        .O(out[11:8]),
        .CI(carryout[7]),
        .CYINIT(1'h0),
        .DI(gene[11:8]),
        .S(prop[11:8])
    );
    CARRY4 carry4_15_12 (
        .CO(carryout[15:12]),
        .O(out[15:12]),
        .CI(carryout[11]),
        .CYINIT(1'h0),
        .DI(gene[15:12]),
        .S(prop[15:12])
    );
    CARRY4 carry4_19_16 (
        .CO(carryout[19:16]),
        .O(out[19:16]),
        .CI(carryout[15]),
        .CYINIT(1'h0),
        .DI({3'h0, gene[16:16]}),
        .S({3'h0, prop[16:16]})
    );
    assign dst0 = {carryout[16], out[16:0]};
endmodule


module comp2_1test_32_12();
    reg [11:0] src0;
    reg [11:0] src1;
    reg [11:0] src2;
    reg [11:0] src3;
    reg [11:0] src4;
    reg [11:0] src5;
    reg [11:0] src6;
    reg [11:0] src7;
    reg [11:0] src8;
    reg [11:0] src9;
    reg [11:0] src10;
    reg [11:0] src11;
    reg [11:0] src12;
    reg [11:0] src13;
    reg [11:0] src14;
    reg [11:0] src15;
    reg [11:0] src16;
    reg [11:0] src17;
    reg [11:0] src18;
    reg [11:0] src19;
    reg [11:0] src20;
    reg [11:0] src21;
    reg [11:0] src22;
    reg [11:0] src23;
    reg [11:0] src24;
    reg [11:0] src25;
    reg [11:0] src26;
    reg [11:0] src27;
    reg [11:0] src28;
    reg [11:0] src29;
    reg [11:0] src30;
    reg [11:0] src31;
    reg [16:0] exp;
    wire [16:0] dst;
    assign test = dst == exp;
    compressor2_1_32_12 compressor2_1_32_12_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst(dst)
    );
    initial begin
        $monitor("0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x 0x%x %x", src0, src1, src2, src3, src4, src5, src6, src7, src8, src9, src10, src11, src12, src13, src14, src15, src16, src17, src18, src19, src20, src21, src22, src23, src24, src25, src26, src27, src28, src29, src30, src31, dst, exp, test);
        src0 <= 12'h90e;
        src1 <= 12'hd02;
        src2 <= 12'h468;
        src3 <= 12'h980;
        src4 <= 12'hfbe;
        src5 <= 12'h1ea;
        src6 <= 12'h3ae;
        src7 <= 12'he26;
        src8 <= 12'h7b3;
        src9 <= 12'h2d9;
        src10 <= 12'h9a8;
        src11 <= 12'h6c3;
        src12 <= 12'h934;
        src13 <= 12'hc42;
        src14 <= 12'hc6f;
        src15 <= 12'h117;
        src16 <= 12'h412;
        src17 <= 12'hc7c;
        src18 <= 12'h778;
        src19 <= 12'hd6;
        src20 <= 12'h3b1;
        src21 <= 12'hb92;
        src22 <= 12'hbe2;
        src23 <= 12'h576;
        src24 <= 12'hb2;
        src25 <= 12'h690;
        src26 <= 12'h2f1;
        src27 <= 12'h9d0;
        src28 <= 12'hb2e;
        src29 <= 12'hd6b;
        src30 <= 12'h1e2;
        src31 <= 12'h766;
        exp <= 17'hf4c2;
        #1
        src0 <= 12'h8d3;
        src1 <= 12'h10a;
        src2 <= 12'he93;
        src3 <= 12'h236;
        src4 <= 12'h180;
        src5 <= 12'hc0f;
        src6 <= 12'h94c;
        src7 <= 12'h205;
        src8 <= 12'h65b;
        src9 <= 12'h57c;
        src10 <= 12'h28a;
        src11 <= 12'hae;
        src12 <= 12'hc14;
        src13 <= 12'h36a;
        src14 <= 12'h5a3;
        src15 <= 12'h57e;
        src16 <= 12'h466;
        src17 <= 12'h17b;
        src18 <= 12'he2c;
        src19 <= 12'h85;
        src20 <= 12'hc33;
        src21 <= 12'ha8d;
        src22 <= 12'hea4;
        src23 <= 12'h515;
        src24 <= 12'h430;
        src25 <= 12'hd75;
        src26 <= 12'h288;
        src27 <= 12'he1d;
        src28 <= 12'hb5;
        src29 <= 12'h3ec;
        src30 <= 12'ha12;
        src31 <= 12'h89a;
        exp <= 17'hd5d6;
        #1
        src0 <= 12'h38d;
        src1 <= 12'h48e;
        src2 <= 12'h728;
        src3 <= 12'h138;
        src4 <= 12'h670;
        src5 <= 12'he88;
        src6 <= 12'h7b4;
        src7 <= 12'hcf5;
        src8 <= 12'h7ae;
        src9 <= 12'heb2;
        src10 <= 12'he30;
        src11 <= 12'h4e6;
        src12 <= 12'h5e9;
        src13 <= 12'he6a;
        src14 <= 12'ha61;
        src15 <= 12'hf76;
        src16 <= 12'h72b;
        src17 <= 12'hb4d;
        src18 <= 12'hebc;
        src19 <= 12'h288;
        src20 <= 12'hf07;
        src21 <= 12'h7e5;
        src22 <= 12'h77;
        src23 <= 12'h9dd;
        src24 <= 12'h9c3;
        src25 <= 12'h82a;
        src26 <= 12'hfd0;
        src27 <= 12'h411;
        src28 <= 12'h8f1;
        src29 <= 12'h38f;
        src30 <= 12'h902;
        src31 <= 12'h43a;
        exp <= 17'h11642;
        #1
        src0 <= 12'h265;
        src1 <= 12'hcbb;
        src2 <= 12'h433;
        src3 <= 12'h4d9;
        src4 <= 12'h66;
        src5 <= 12'hbe1;
        src6 <= 12'h1a6;
        src7 <= 12'hcb2;
        src8 <= 12'h21d;
        src9 <= 12'hf37;
        src10 <= 12'h53a;
        src11 <= 12'h5bf;
        src12 <= 12'hbd7;
        src13 <= 12'hd4f;
        src14 <= 12'h18f;
        src15 <= 12'h83f;
        src16 <= 12'he45;
        src17 <= 12'h4f1;
        src18 <= 12'h323;
        src19 <= 12'h1c3;
        src20 <= 12'he17;
        src21 <= 12'h89d;
        src22 <= 12'h371;
        src23 <= 12'h2fd;
        src24 <= 12'h74e;
        src25 <= 12'hcee;
        src26 <= 12'h8e2;
        src27 <= 12'h58e;
        src28 <= 12'h825;
        src29 <= 12'he38;
        src30 <= 12'h811;
        src31 <= 12'hc1b;
        exp <= 17'hf47f;
        #1
        src0 <= 12'h51d;
        src1 <= 12'h2b8;
        src2 <= 12'h8e2;
        src3 <= 12'hc55;
        src4 <= 12'h56c;
        src5 <= 12'h584;
        src6 <= 12'h97a;
        src7 <= 12'h736;
        src8 <= 12'h6ad;
        src9 <= 12'h598;
        src10 <= 12'h103;
        src11 <= 12'hf0d;
        src12 <= 12'hd83;
        src13 <= 12'h703;
        src14 <= 12'h4fe;
        src15 <= 12'hdd3;
        src16 <= 12'hc37;
        src17 <= 12'h9c;
        src18 <= 12'hd84;
        src19 <= 12'hfe2;
        src20 <= 12'ha3a;
        src21 <= 12'h3cc;
        src22 <= 12'h53b;
        src23 <= 12'h62e;
        src24 <= 12'h698;
        src25 <= 12'h293;
        src26 <= 12'hec7;
        src27 <= 12'h7e;
        src28 <= 12'hdce;
        src29 <= 12'he83;
        src30 <= 12'h980;
        src31 <= 12'h259;
        exp <= 17'h1009a;
        #1
        src0 <= 12'h63d;
        src1 <= 12'hfcc;
        src2 <= 12'hd17;
        src3 <= 12'h337;
        src4 <= 12'hc6;
        src5 <= 12'h1a0;
        src6 <= 12'hd4a;
        src7 <= 12'h116;
        src8 <= 12'had9;
        src9 <= 12'hb43;
        src10 <= 12'h6a7;
        src11 <= 12'hffd;
        src12 <= 12'hca7;
        src13 <= 12'h4df;
        src14 <= 12'ha91;
        src15 <= 12'h6f2;
        src16 <= 12'hba6;
        src17 <= 12'hbeb;
        src18 <= 12'hb7f;
        src19 <= 12'h111;
        src20 <= 12'he2c;
        src21 <= 12'h481;
        src22 <= 12'hd03;
        src23 <= 12'h85c;
        src24 <= 12'h349;
        src25 <= 12'h4c8;
        src26 <= 12'h9a4;
        src27 <= 12'hf47;
        src28 <= 12'hbaf;
        src29 <= 12'h9c0;
        src30 <= 12'h17e;
        src31 <= 12'h156;
        exp <= 17'h10c52;
        #1
        src0 <= 12'had1;
        src1 <= 12'hbcd;
        src2 <= 12'hd3f;
        src3 <= 12'hfa7;
        src4 <= 12'ha3c;
        src5 <= 12'hb7d;
        src6 <= 12'h3b5;
        src7 <= 12'hbf6;
        src8 <= 12'h361;
        src9 <= 12'ha29;
        src10 <= 12'h3ec;
        src11 <= 12'h190;
        src12 <= 12'h26e;
        src13 <= 12'hdc7;
        src14 <= 12'h24e;
        src15 <= 12'h783;
        src16 <= 12'h79e;
        src17 <= 12'h990;
        src18 <= 12'hef0;
        src19 <= 12'h51a;
        src20 <= 12'h1d9;
        src21 <= 12'he41;
        src22 <= 12'h8;
        src23 <= 12'hd57;
        src24 <= 12'hed4;
        src25 <= 12'hc49;
        src26 <= 12'hb57;
        src27 <= 12'hc54;
        src28 <= 12'hbf0;
        src29 <= 12'h126;
        src30 <= 12'hf47;
        src31 <= 12'hecd;
        exp <= 17'h12697;
        #1
        src0 <= 12'h7bd;
        src1 <= 12'h494;
        src2 <= 12'h8e2;
        src3 <= 12'h3d9;
        src4 <= 12'h224;
        src5 <= 12'h529;
        src6 <= 12'hdb2;
        src7 <= 12'h34;
        src8 <= 12'hf4f;
        src9 <= 12'h3ae;
        src10 <= 12'he7d;
        src11 <= 12'h978;
        src12 <= 12'head;
        src13 <= 12'hac2;
        src14 <= 12'ha86;
        src15 <= 12'hb05;
        src16 <= 12'h98f;
        src17 <= 12'haa;
        src18 <= 12'h762;
        src19 <= 12'h4f4;
        src20 <= 12'heb6;
        src21 <= 12'h87d;
        src22 <= 12'hf6a;
        src23 <= 12'hb61;
        src24 <= 12'h5ac;
        src25 <= 12'hc24;
        src26 <= 12'hb4b;
        src27 <= 12'h441;
        src28 <= 12'h83d;
        src29 <= 12'hf3f;
        src30 <= 12'hb56;
        src31 <= 12'hb63;
        exp <= 17'h12049;
        #1
        src0 <= 12'h87e;
        src1 <= 12'hcf5;
        src2 <= 12'h3e0;
        src3 <= 12'h414;
        src4 <= 12'haa8;
        src5 <= 12'hca8;
        src6 <= 12'hf5f;
        src7 <= 12'hd2b;
        src8 <= 12'h51f;
        src9 <= 12'h2a4;
        src10 <= 12'he3e;
        src11 <= 12'h3bc;
        src12 <= 12'hd4a;
        src13 <= 12'hacd;
        src14 <= 12'ha82;
        src15 <= 12'h4ad;
        src16 <= 12'h5b7;
        src17 <= 12'hd4e;
        src18 <= 12'h6c6;
        src19 <= 12'h420;
        src20 <= 12'h2b0;
        src21 <= 12'hf16;
        src22 <= 12'h32a;
        src23 <= 12'h20b;
        src24 <= 12'h9cd;
        src25 <= 12'hd9a;
        src26 <= 12'hc1c;
        src27 <= 12'hb45;
        src28 <= 12'h907;
        src29 <= 12'hb7c;
        src30 <= 12'h763;
        src31 <= 12'h501;
        exp <= 17'h116d9;
        #1
        src0 <= 12'h86b;
        src1 <= 12'h640;
        src2 <= 12'he82;
        src3 <= 12'hb7a;
        src4 <= 12'h972;
        src5 <= 12'h348;
        src6 <= 12'h320;
        src7 <= 12'h74d;
        src8 <= 12'hd97;
        src9 <= 12'h1cb;
        src10 <= 12'h3e8;
        src11 <= 12'hfc6;
        src12 <= 12'h8dd;
        src13 <= 12'h3ec;
        src14 <= 12'hda1;
        src15 <= 12'hbf6;
        src16 <= 12'h15;
        src17 <= 12'hb1a;
        src18 <= 12'hdc1;
        src19 <= 12'h882;
        src20 <= 12'h8;
        src21 <= 12'h40;
        src22 <= 12'h35c;
        src23 <= 12'hc04;
        src24 <= 12'ha7a;
        src25 <= 12'hef6;
        src26 <= 12'h80c;
        src27 <= 12'h1b6;
        src28 <= 12'h641;
        src29 <= 12'hbb4;
        src30 <= 12'h900;
        src31 <= 12'h743;
        exp <= 17'hffc2;
        #1
        src0 <= 12'he8;
        src1 <= 12'h7b0;
        src2 <= 12'hcfe;
        src3 <= 12'h7c8;
        src4 <= 12'h9b6;
        src5 <= 12'h13f;
        src6 <= 12'h62e;
        src7 <= 12'h117;
        src8 <= 12'haae;
        src9 <= 12'h10c;
        src10 <= 12'h89b;
        src11 <= 12'hced;
        src12 <= 12'h7;
        src13 <= 12'h8fb;
        src14 <= 12'hfa9;
        src15 <= 12'h485;
        src16 <= 12'he8;
        src17 <= 12'h2fa;
        src18 <= 12'h330;
        src19 <= 12'h279;
        src20 <= 12'hee9;
        src21 <= 12'hadf;
        src22 <= 12'hb55;
        src23 <= 12'h655;
        src24 <= 12'h14d;
        src25 <= 12'h74b;
        src26 <= 12'hb4c;
        src27 <= 12'h1b3;
        src28 <= 12'hf3c;
        src29 <= 12'h503;
        src30 <= 12'h89c;
        src31 <= 12'h88a;
        exp <= 17'hde03;
        #1
        src0 <= 12'h407;
        src1 <= 12'hb0f;
        src2 <= 12'hfd1;
        src3 <= 12'h76f;
        src4 <= 12'h627;
        src5 <= 12'hc7a;
        src6 <= 12'hfa7;
        src7 <= 12'hba;
        src8 <= 12'h154;
        src9 <= 12'hc74;
        src10 <= 12'h259;
        src11 <= 12'ha44;
        src12 <= 12'ha7e;
        src13 <= 12'h9bc;
        src14 <= 12'h33d;
        src15 <= 12'h7a2;
        src16 <= 12'hf1e;
        src17 <= 12'h1a3;
        src18 <= 12'h1e0;
        src19 <= 12'h935;
        src20 <= 12'h5d9;
        src21 <= 12'hb06;
        src22 <= 12'hd4;
        src23 <= 12'he14;
        src24 <= 12'hbec;
        src25 <= 12'h54c;
        src26 <= 12'hc39;
        src27 <= 12'hdeb;
        src28 <= 12'h309;
        src29 <= 12'hdbe;
        src30 <= 12'h9c;
        src31 <= 12'h632;
        exp <= 17'h10164;
        #1
        src0 <= 12'he33;
        src1 <= 12'hbef;
        src2 <= 12'h318;
        src3 <= 12'hc84;
        src4 <= 12'h5d0;
        src5 <= 12'h2ac;
        src6 <= 12'h962;
        src7 <= 12'h634;
        src8 <= 12'hfeb;
        src9 <= 12'h21c;
        src10 <= 12'h5c5;
        src11 <= 12'hb18;
        src12 <= 12'h2cb;
        src13 <= 12'ha52;
        src14 <= 12'hf9;
        src15 <= 12'ha4c;
        src16 <= 12'h75e;
        src17 <= 12'h2a8;
        src18 <= 12'hd9b;
        src19 <= 12'ha81;
        src20 <= 12'he43;
        src21 <= 12'h293;
        src22 <= 12'h15c;
        src23 <= 12'hfc8;
        src24 <= 12'h123;
        src25 <= 12'h729;
        src26 <= 12'h914;
        src27 <= 12'heac;
        src28 <= 12'h5a8;
        src29 <= 12'ha1c;
        src30 <= 12'hd7;
        src31 <= 12'h859;
        exp <= 17'hfa32;
        #1
        src0 <= 12'hc09;
        src1 <= 12'ha44;
        src2 <= 12'h6bd;
        src3 <= 12'he81;
        src4 <= 12'h1d1;
        src5 <= 12'hf90;
        src6 <= 12'h50f;
        src7 <= 12'hf53;
        src8 <= 12'hc8f;
        src9 <= 12'h28a;
        src10 <= 12'he8c;
        src11 <= 12'hc59;
        src12 <= 12'h90c;
        src13 <= 12'hdf8;
        src14 <= 12'haef;
        src15 <= 12'h680;
        src16 <= 12'hd7c;
        src17 <= 12'hb5;
        src18 <= 12'h261;
        src19 <= 12'h1f0;
        src20 <= 12'hd72;
        src21 <= 12'ha34;
        src22 <= 12'h4e9;
        src23 <= 12'he52;
        src24 <= 12'hc10;
        src25 <= 12'h89a;
        src26 <= 12'h230;
        src27 <= 12'hfac;
        src28 <= 12'hd9f;
        src29 <= 12'h790;
        src30 <= 12'h2b8;
        src31 <= 12'h5bc;
        exp <= 17'h1254b;
        #1
        src0 <= 12'h832;
        src1 <= 12'h57a;
        src2 <= 12'h723;
        src3 <= 12'h5b2;
        src4 <= 12'hadb;
        src5 <= 12'h632;
        src6 <= 12'h6bc;
        src7 <= 12'h244;
        src8 <= 12'hb7c;
        src9 <= 12'h498;
        src10 <= 12'h634;
        src11 <= 12'h1ae;
        src12 <= 12'he8c;
        src13 <= 12'h41c;
        src14 <= 12'hc3c;
        src15 <= 12'h9e0;
        src16 <= 12'h302;
        src17 <= 12'h262;
        src18 <= 12'h9df;
        src19 <= 12'h20f;
        src20 <= 12'h57d;
        src21 <= 12'h2dd;
        src22 <= 12'hcfd;
        src23 <= 12'h509;
        src24 <= 12'hc75;
        src25 <= 12'h220;
        src26 <= 12'h7f8;
        src27 <= 12'hec8;
        src28 <= 12'hb96;
        src29 <= 12'h85b;
        src30 <= 12'h3be;
        src31 <= 12'h497;
        exp <= 17'he295;
        #1
        src0 <= 12'h1ce;
        src1 <= 12'h62a;
        src2 <= 12'h2d;
        src3 <= 12'h18e;
        src4 <= 12'hf;
        src5 <= 12'he3;
        src6 <= 12'hc52;
        src7 <= 12'h7d8;
        src8 <= 12'h465;
        src9 <= 12'hc57;
        src10 <= 12'hee3;
        src11 <= 12'h13d;
        src12 <= 12'hf6a;
        src13 <= 12'hc3d;
        src14 <= 12'h35e;
        src15 <= 12'h3b7;
        src16 <= 12'hafc;
        src17 <= 12'h147;
        src18 <= 12'hafe;
        src19 <= 12'hc92;
        src20 <= 12'h95b;
        src21 <= 12'h160;
        src22 <= 12'he6a;
        src23 <= 12'h681;
        src24 <= 12'h4ec;
        src25 <= 12'h854;
        src26 <= 12'hfc8;
        src27 <= 12'ha5;
        src28 <= 12'h4bb;
        src29 <= 12'h635;
        src30 <= 12'hdc6;
        src31 <= 12'h42a;
        exp <= 17'he06d;
        #1
        src0 <= 12'h8e3;
        src1 <= 12'h453;
        src2 <= 12'hba3;
        src3 <= 12'h101;
        src4 <= 12'hac3;
        src5 <= 12'h2d7;
        src6 <= 12'h115;
        src7 <= 12'hedd;
        src8 <= 12'ha86;
        src9 <= 12'he04;
        src10 <= 12'h611;
        src11 <= 12'hdf7;
        src12 <= 12'h186;
        src13 <= 12'h6b6;
        src14 <= 12'h8c9;
        src15 <= 12'h744;
        src16 <= 12'h816;
        src17 <= 12'hd56;
        src18 <= 12'h68e;
        src19 <= 12'hf5f;
        src20 <= 12'hc23;
        src21 <= 12'h96e;
        src22 <= 12'h68d;
        src23 <= 12'h560;
        src24 <= 12'h6de;
        src25 <= 12'h14a;
        src26 <= 12'h805;
        src27 <= 12'hee5;
        src28 <= 12'h447;
        src29 <= 12'h184;
        src30 <= 12'h181;
        src31 <= 12'h400;
        exp <= 17'hf376;
        #1
        src0 <= 12'h72;
        src1 <= 12'h56;
        src2 <= 12'h592;
        src3 <= 12'h539;
        src4 <= 12'hb1f;
        src5 <= 12'hf78;
        src6 <= 12'h280;
        src7 <= 12'hc2c;
        src8 <= 12'h9ac;
        src9 <= 12'h3fb;
        src10 <= 12'h13a;
        src11 <= 12'h802;
        src12 <= 12'h592;
        src13 <= 12'h45b;
        src14 <= 12'h81b;
        src15 <= 12'hb46;
        src16 <= 12'h204;
        src17 <= 12'h831;
        src18 <= 12'he00;
        src19 <= 12'h8ee;
        src20 <= 12'h55e;
        src21 <= 12'hf4;
        src22 <= 12'h470;
        src23 <= 12'he82;
        src24 <= 12'hbbe;
        src25 <= 12'ha59;
        src26 <= 12'h55e;
        src27 <= 12'h45d;
        src28 <= 12'h93b;
        src29 <= 12'h6d;
        src30 <= 12'h77;
        src31 <= 12'h607;
        exp <= 17'hd366;
        #1
        src0 <= 12'ha98;
        src1 <= 12'h844;
        src2 <= 12'h442;
        src3 <= 12'h920;
        src4 <= 12'ha9d;
        src5 <= 12'h3f6;
        src6 <= 12'h53c;
        src7 <= 12'h2b4;
        src8 <= 12'h4ef;
        src9 <= 12'h295;
        src10 <= 12'hc9e;
        src11 <= 12'h4c1;
        src12 <= 12'h74d;
        src13 <= 12'h3d8;
        src14 <= 12'h6c4;
        src15 <= 12'h6f2;
        src16 <= 12'h40b;
        src17 <= 12'h632;
        src18 <= 12'hc5c;
        src19 <= 12'h60e;
        src20 <= 12'hd49;
        src21 <= 12'hfda;
        src22 <= 12'h232;
        src23 <= 12'hf9d;
        src24 <= 12'he5e;
        src25 <= 12'he1b;
        src26 <= 12'h662;
        src27 <= 12'he2a;
        src28 <= 12'hbc0;
        src29 <= 12'hdf0;
        src30 <= 12'hcb5;
        src31 <= 12'h227;
        exp <= 17'h10da9;
        #1
        src0 <= 12'h578;
        src1 <= 12'h2bb;
        src2 <= 12'h784;
        src3 <= 12'hd3a;
        src4 <= 12'h7eb;
        src5 <= 12'h85d;
        src6 <= 12'had6;
        src7 <= 12'h52;
        src8 <= 12'he1d;
        src9 <= 12'h7a0;
        src10 <= 12'h915;
        src11 <= 12'h72b;
        src12 <= 12'h9b;
        src13 <= 12'hea3;
        src14 <= 12'h22a;
        src15 <= 12'hd8;
        src16 <= 12'h8b0;
        src17 <= 12'hca8;
        src18 <= 12'hbf2;
        src19 <= 12'hf2c;
        src20 <= 12'hd79;
        src21 <= 12'h2ae;
        src22 <= 12'ha43;
        src23 <= 12'hf23;
        src24 <= 12'hf3e;
        src25 <= 12'h1e;
        src26 <= 12'h1a7;
        src27 <= 12'hd5f;
        src28 <= 12'h2ca;
        src29 <= 12'h2df;
        src30 <= 12'h4ab;
        src31 <= 12'h5c1;
        exp <= 17'hf918;
        #1
        src0 <= 12'h643;
        src1 <= 12'hcaa;
        src2 <= 12'h660;
        src3 <= 12'h6af;
        src4 <= 12'h321;
        src5 <= 12'hbff;
        src6 <= 12'h409;
        src7 <= 12'habd;
        src8 <= 12'h1a0;
        src9 <= 12'hbfe;
        src10 <= 12'h569;
        src11 <= 12'he13;
        src12 <= 12'h699;
        src13 <= 12'h4e8;
        src14 <= 12'h723;
        src15 <= 12'hab0;
        src16 <= 12'hf8f;
        src17 <= 12'hcf;
        src18 <= 12'hb48;
        src19 <= 12'h7f5;
        src20 <= 12'h475;
        src21 <= 12'h547;
        src22 <= 12'hd7f;
        src23 <= 12'ha76;
        src24 <= 12'hac7;
        src25 <= 12'he8a;
        src26 <= 12'h8aa;
        src27 <= 12'hb66;
        src28 <= 12'h318;
        src29 <= 12'h3e0;
        src30 <= 12'h6e3;
        src31 <= 12'h4bc;
        exp <= 17'h10194;
        #1
        src0 <= 12'h50e;
        src1 <= 12'h2fd;
        src2 <= 12'h7e3;
        src3 <= 12'h240;
        src4 <= 12'h5a6;
        src5 <= 12'h8bd;
        src6 <= 12'h675;
        src7 <= 12'had9;
        src8 <= 12'h2c1;
        src9 <= 12'h926;
        src10 <= 12'hbc5;
        src11 <= 12'h730;
        src12 <= 12'h31d;
        src13 <= 12'hb48;
        src14 <= 12'he2;
        src15 <= 12'h808;
        src16 <= 12'h9a4;
        src17 <= 12'h42d;
        src18 <= 12'h69f;
        src19 <= 12'h471;
        src20 <= 12'h248;
        src21 <= 12'hca0;
        src22 <= 12'h779;
        src23 <= 12'h812;
        src24 <= 12'h90d;
        src25 <= 12'hba3;
        src26 <= 12'he8;
        src27 <= 12'h226;
        src28 <= 12'he97;
        src29 <= 12'h182;
        src30 <= 12'h2f9;
        src31 <= 12'h290;
        exp <= 17'hccbe;
        #1
        src0 <= 12'h53b;
        src1 <= 12'h307;
        src2 <= 12'hf01;
        src3 <= 12'hc6d;
        src4 <= 12'h75b;
        src5 <= 12'hb58;
        src6 <= 12'hf2a;
        src7 <= 12'h5f3;
        src8 <= 12'h744;
        src9 <= 12'h486;
        src10 <= 12'hfc0;
        src11 <= 12'h762;
        src12 <= 12'h334;
        src13 <= 12'h8b4;
        src14 <= 12'hd9f;
        src15 <= 12'he24;
        src16 <= 12'h4a9;
        src17 <= 12'h142;
        src18 <= 12'hf82;
        src19 <= 12'h209;
        src20 <= 12'h8de;
        src21 <= 12'h341;
        src22 <= 12'h92f;
        src23 <= 12'h7f4;
        src24 <= 12'hc55;
        src25 <= 12'h8ad;
        src26 <= 12'hb1c;
        src27 <= 12'hde9;
        src28 <= 12'h249;
        src29 <= 12'h3f1;
        src30 <= 12'h4ea;
        src31 <= 12'h2e;
        exp <= 17'h10428;
        #1
        src0 <= 12'h9dd;
        src1 <= 12'hfa8;
        src2 <= 12'h887;
        src3 <= 12'hc9d;
        src4 <= 12'h2db;
        src5 <= 12'h198;
        src6 <= 12'hfe9;
        src7 <= 12'h618;
        src8 <= 12'h4d6;
        src9 <= 12'h452;
        src10 <= 12'hfb9;
        src11 <= 12'h65f;
        src12 <= 12'h233;
        src13 <= 12'h5ea;
        src14 <= 12'hc2e;
        src15 <= 12'h60e;
        src16 <= 12'hbf8;
        src17 <= 12'h800;
        src18 <= 12'ha7a;
        src19 <= 12'h3ca;
        src20 <= 12'h101;
        src21 <= 12'hc4d;
        src22 <= 12'ha08;
        src23 <= 12'ha54;
        src24 <= 12'ha1c;
        src25 <= 12'h8ff;
        src26 <= 12'h897;
        src27 <= 12'hd5b;
        src28 <= 12'he31;
        src29 <= 12'hdb5;
        src30 <= 12'h502;
        src31 <= 12'hc2b;
        exp <= 17'h11cbc;
        #1
        src0 <= 12'heeb;
        src1 <= 12'h69f;
        src2 <= 12'h218;
        src3 <= 12'h76d;
        src4 <= 12'h62b;
        src5 <= 12'h219;
        src6 <= 12'h561;
        src7 <= 12'h4c6;
        src8 <= 12'hb89;
        src9 <= 12'h1df;
        src10 <= 12'h355;
        src11 <= 12'h410;
        src12 <= 12'hffa;
        src13 <= 12'h499;
        src14 <= 12'hfcf;
        src15 <= 12'he99;
        src16 <= 12'h56b;
        src17 <= 12'h9dd;
        src18 <= 12'h8f2;
        src19 <= 12'h953;
        src20 <= 12'h2b1;
        src21 <= 12'h1da;
        src22 <= 12'h694;
        src23 <= 12'he73;
        src24 <= 12'had1;
        src25 <= 12'hfc1;
        src26 <= 12'hda0;
        src27 <= 12'had6;
        src28 <= 12'h814;
        src29 <= 12'h453;
        src30 <= 12'hf5;
        src31 <= 12'h151;
        exp <= 17'hf616;
        #1
        src0 <= 12'h79c;
        src1 <= 12'h68f;
        src2 <= 12'h710;
        src3 <= 12'he9;
        src4 <= 12'h6df;
        src5 <= 12'h4e;
        src6 <= 12'h12b;
        src7 <= 12'h56c;
        src8 <= 12'h968;
        src9 <= 12'he13;
        src10 <= 12'h728;
        src11 <= 12'h6d1;
        src12 <= 12'h7f6;
        src13 <= 12'hb53;
        src14 <= 12'hb88;
        src15 <= 12'hf35;
        src16 <= 12'h39d;
        src17 <= 12'ha3f;
        src18 <= 12'ha40;
        src19 <= 12'h9c8;
        src20 <= 12'h321;
        src21 <= 12'h412;
        src22 <= 12'he23;
        src23 <= 12'ha62;
        src24 <= 12'hf83;
        src25 <= 12'h19f;
        src26 <= 12'h45d;
        src27 <= 12'h590;
        src28 <= 12'hcee;
        src29 <= 12'hcd0;
        src30 <= 12'hcd7;
        src31 <= 12'he3a;
        exp <= 17'h108dc;
        #1
        src0 <= 12'hf0c;
        src1 <= 12'h31f;
        src2 <= 12'he;
        src3 <= 12'hfdc;
        src4 <= 12'hd26;
        src5 <= 12'hc7d;
        src6 <= 12'h7ac;
        src7 <= 12'he6f;
        src8 <= 12'h96e;
        src9 <= 12'hee3;
        src10 <= 12'haed;
        src11 <= 12'h1ec;
        src12 <= 12'h8af;
        src13 <= 12'ha7e;
        src14 <= 12'hfe9;
        src15 <= 12'h9eb;
        src16 <= 12'hf9a;
        src17 <= 12'hd91;
        src18 <= 12'h2c9;
        src19 <= 12'hedf;
        src20 <= 12'hc7d;
        src21 <= 12'hb78;
        src22 <= 12'h1d6;
        src23 <= 12'hcad;
        src24 <= 12'h34c;
        src25 <= 12'hee0;
        src26 <= 12'hd6;
        src27 <= 12'hc96;
        src28 <= 12'he5a;
        src29 <= 12'hb9e;
        src30 <= 12'h6c;
        src31 <= 12'hc36;
        exp <= 17'h13f7b;
        #1
        src0 <= 12'hf2d;
        src1 <= 12'hc9e;
        src2 <= 12'ha11;
        src3 <= 12'hc93;
        src4 <= 12'h40a;
        src5 <= 12'h45d;
        src6 <= 12'h864;
        src7 <= 12'h6fb;
        src8 <= 12'h243;
        src9 <= 12'hcc1;
        src10 <= 12'h437;
        src11 <= 12'h147;
        src12 <= 12'h31a;
        src13 <= 12'hce6;
        src14 <= 12'h656;
        src15 <= 12'h72b;
        src16 <= 12'hacb;
        src17 <= 12'h794;
        src18 <= 12'hb24;
        src19 <= 12'h946;
        src20 <= 12'h819;
        src21 <= 12'h13c;
        src22 <= 12'h3c1;
        src23 <= 12'h4bb;
        src24 <= 12'h71e;
        src25 <= 12'h34b;
        src26 <= 12'h4b6;
        src27 <= 12'h292;
        src28 <= 12'heed;
        src29 <= 12'hb88;
        src30 <= 12'hbb2;
        src31 <= 12'h9a3;
        exp <= 17'hf64d;
        #1
        src0 <= 12'h4c2;
        src1 <= 12'h1b2;
        src2 <= 12'h5cc;
        src3 <= 12'h1fa;
        src4 <= 12'h831;
        src5 <= 12'h96d;
        src6 <= 12'ha1d;
        src7 <= 12'h756;
        src8 <= 12'h5da;
        src9 <= 12'h55b;
        src10 <= 12'h5d;
        src11 <= 12'hb46;
        src12 <= 12'hb26;
        src13 <= 12'h4ce;
        src14 <= 12'h92d;
        src15 <= 12'ha44;
        src16 <= 12'hc69;
        src17 <= 12'h72c;
        src18 <= 12'h3d7;
        src19 <= 12'hd5e;
        src20 <= 12'hb59;
        src21 <= 12'hc0e;
        src22 <= 12'h187;
        src23 <= 12'h18c;
        src24 <= 12'h3f3;
        src25 <= 12'hb73;
        src26 <= 12'h113;
        src27 <= 12'hf18;
        src28 <= 12'h1a2;
        src29 <= 12'hae8;
        src30 <= 12'h60;
        src31 <= 12'hdf4;
        exp <= 17'he53b;
        #1
        src0 <= 12'h112;
        src1 <= 12'hdb;
        src2 <= 12'h8f0;
        src3 <= 12'hbcb;
        src4 <= 12'hedc;
        src5 <= 12'h386;
        src6 <= 12'h96e;
        src7 <= 12'heb3;
        src8 <= 12'h8a1;
        src9 <= 12'hc08;
        src10 <= 12'hf1e;
        src11 <= 12'h612;
        src12 <= 12'hd4b;
        src13 <= 12'h2ed;
        src14 <= 12'hc9c;
        src15 <= 12'h5e5;
        src16 <= 12'h9bc;
        src17 <= 12'h81d;
        src18 <= 12'h45f;
        src19 <= 12'he23;
        src20 <= 12'h9c2;
        src21 <= 12'ha99;
        src22 <= 12'heab;
        src23 <= 12'h34e;
        src24 <= 12'h847;
        src25 <= 12'hc4e;
        src26 <= 12'hcb4;
        src27 <= 12'h322;
        src28 <= 12'hfb9;
        src29 <= 12'h192;
        src30 <= 12'h33a;
        src31 <= 12'h3ac;
        exp <= 17'h11508;
        #1
        src0 <= 12'hb15;
        src1 <= 12'h461;
        src2 <= 12'h21f;
        src3 <= 12'h709;
        src4 <= 12'hb0a;
        src5 <= 12'hda;
        src6 <= 12'h122;
        src7 <= 12'ha0f;
        src8 <= 12'h1cb;
        src9 <= 12'h5cd;
        src10 <= 12'h506;
        src11 <= 12'h1f2;
        src12 <= 12'h24;
        src13 <= 12'hf02;
        src14 <= 12'h729;
        src15 <= 12'h4d1;
        src16 <= 12'heab;
        src17 <= 12'hb95;
        src18 <= 12'h300;
        src19 <= 12'hbec;
        src20 <= 12'h597;
        src21 <= 12'h579;
        src22 <= 12'hb56;
        src23 <= 12'h57c;
        src24 <= 12'hc25;
        src25 <= 12'hde5;
        src26 <= 12'h8a7;
        src27 <= 12'h7f1;
        src28 <= 12'hb1e;
        src29 <= 12'h710;
        src30 <= 12'h469;
        src31 <= 12'h4f7;
        exp <= 17'he4a1;
        #1
        src0 <= 12'hfc;
        src1 <= 12'h89e;
        src2 <= 12'h82;
        src3 <= 12'h751;
        src4 <= 12'hef7;
        src5 <= 12'h5a3;
        src6 <= 12'hdf9;
        src7 <= 12'hcda;
        src8 <= 12'h9b5;
        src9 <= 12'h333;
        src10 <= 12'hd19;
        src11 <= 12'h31c;
        src12 <= 12'h7fb;
        src13 <= 12'h965;
        src14 <= 12'h41b;
        src15 <= 12'h8ec;
        src16 <= 12'heb;
        src17 <= 12'h7ad;
        src18 <= 12'h425;
        src19 <= 12'hb3a;
        src20 <= 12'h869;
        src21 <= 12'h600;
        src22 <= 12'he79;
        src23 <= 12'h4ff;
        src24 <= 12'h3f8;
        src25 <= 12'h2be;
        src26 <= 12'h5e5;
        src27 <= 12'h772;
        src28 <= 12'hb6;
        src29 <= 12'h5b6;
        src30 <= 12'he74;
        src31 <= 12'h68b;
        exp <= 17'he5ae;
        #1
        src0 <= 12'h15f;
        src1 <= 12'h399;
        src2 <= 12'hd29;
        src3 <= 12'h394;
        src4 <= 12'h97a;
        src5 <= 12'haea;
        src6 <= 12'ha92;
        src7 <= 12'hd8d;
        src8 <= 12'h7bc;
        src9 <= 12'heb0;
        src10 <= 12'hafd;
        src11 <= 12'h668;
        src12 <= 12'h6e1;
        src13 <= 12'hef3;
        src14 <= 12'h129;
        src15 <= 12'h7aa;
        src16 <= 12'head;
        src17 <= 12'hb69;
        src18 <= 12'h31c;
        src19 <= 12'h3d2;
        src20 <= 12'h85a;
        src21 <= 12'h7af;
        src22 <= 12'hf6f;
        src23 <= 12'h9d7;
        src24 <= 12'hcd5;
        src25 <= 12'h3ef;
        src26 <= 12'h253;
        src27 <= 12'h351;
        src28 <= 12'h8b1;
        src29 <= 12'h13b;
        src30 <= 12'h702;
        src31 <= 12'h82a;
        exp <= 17'h10283;
        #1
        src0 <= 12'haa;
        src1 <= 12'h8f6;
        src2 <= 12'h210;
        src3 <= 12'hb80;
        src4 <= 12'h264;
        src5 <= 12'h6fc;
        src6 <= 12'h8f0;
        src7 <= 12'hb2a;
        src8 <= 12'h22c;
        src9 <= 12'h891;
        src10 <= 12'hf16;
        src11 <= 12'h939;
        src12 <= 12'hdf2;
        src13 <= 12'h2cd;
        src14 <= 12'he5d;
        src15 <= 12'h600;
        src16 <= 12'h595;
        src17 <= 12'h478;
        src18 <= 12'hf81;
        src19 <= 12'h890;
        src20 <= 12'ha0;
        src21 <= 12'he4b;
        src22 <= 12'hff1;
        src23 <= 12'hec7;
        src24 <= 12'h297;
        src25 <= 12'hdd;
        src26 <= 12'h68b;
        src27 <= 12'ha2d;
        src28 <= 12'hc32;
        src29 <= 12'h511;
        src30 <= 12'habc;
        src31 <= 12'ha44;
        exp <= 17'h10702;
        #1
        src0 <= 12'h70c;
        src1 <= 12'hdbd;
        src2 <= 12'hfcf;
        src3 <= 12'h806;
        src4 <= 12'hee4;
        src5 <= 12'he25;
        src6 <= 12'h3b;
        src7 <= 12'hf55;
        src8 <= 12'h566;
        src9 <= 12'hb6d;
        src10 <= 12'hf49;
        src11 <= 12'h4d;
        src12 <= 12'h9a1;
        src13 <= 12'haf8;
        src14 <= 12'h2fc;
        src15 <= 12'h3a2;
        src16 <= 12'h321;
        src17 <= 12'h6f7;
        src18 <= 12'ha8a;
        src19 <= 12'h6a;
        src20 <= 12'hb0f;
        src21 <= 12'hce8;
        src22 <= 12'h4e7;
        src23 <= 12'h67e;
        src24 <= 12'hef;
        src25 <= 12'h716;
        src26 <= 12'h13b;
        src27 <= 12'hf4c;
        src28 <= 12'h832;
        src29 <= 12'h117;
        src30 <= 12'ha6f;
        src31 <= 12'h520;
        exp <= 17'hfea3;
        #1
        src0 <= 12'habc;
        src1 <= 12'hcb0;
        src2 <= 12'h83;
        src3 <= 12'hbdf;
        src4 <= 12'h8cf;
        src5 <= 12'h511;
        src6 <= 12'h772;
        src7 <= 12'h251;
        src8 <= 12'h109;
        src9 <= 12'hca7;
        src10 <= 12'h10f;
        src11 <= 12'hff5;
        src12 <= 12'h7ab;
        src13 <= 12'h97d;
        src14 <= 12'hf0e;
        src15 <= 12'h86;
        src16 <= 12'h334;
        src17 <= 12'h164;
        src18 <= 12'h80b;
        src19 <= 12'ha6d;
        src20 <= 12'h3f9;
        src21 <= 12'hda1;
        src22 <= 12'haa2;
        src23 <= 12'h74a;
        src24 <= 12'h8c0;
        src25 <= 12'hb39;
        src26 <= 12'hb4b;
        src27 <= 12'hb84;
        src28 <= 12'hdb7;
        src29 <= 12'hecb;
        src30 <= 12'h599;
        src31 <= 12'h5a8;
        exp <= 17'h10802;
        #1
        src0 <= 12'hfbe;
        src1 <= 12'ha6d;
        src2 <= 12'hee1;
        src3 <= 12'hc06;
        src4 <= 12'h663;
        src5 <= 12'h81a;
        src6 <= 12'h321;
        src7 <= 12'hcd6;
        src8 <= 12'hbfe;
        src9 <= 12'h193;
        src10 <= 12'h8cc;
        src11 <= 12'h4fc;
        src12 <= 12'he5;
        src13 <= 12'hc7c;
        src14 <= 12'h9df;
        src15 <= 12'ha9b;
        src16 <= 12'hc98;
        src17 <= 12'h3d7;
        src18 <= 12'hc71;
        src19 <= 12'h82;
        src20 <= 12'hb73;
        src21 <= 12'hc7b;
        src22 <= 12'hc6b;
        src23 <= 12'hda0;
        src24 <= 12'he5f;
        src25 <= 12'h19d;
        src26 <= 12'h8b;
        src27 <= 12'h29c;
        src28 <= 12'hb02;
        src29 <= 12'hc69;
        src30 <= 12'h8a9;
        src31 <= 12'hf0e;
        exp <= 17'h1225a;
        #1
        src0 <= 12'h8af;
        src1 <= 12'hadb;
        src2 <= 12'h3ce;
        src3 <= 12'h26;
        src4 <= 12'h4fe;
        src5 <= 12'h90a;
        src6 <= 12'hce5;
        src7 <= 12'ha48;
        src8 <= 12'h273;
        src9 <= 12'h31e;
        src10 <= 12'h6dd;
        src11 <= 12'hf3f;
        src12 <= 12'h529;
        src13 <= 12'h8ad;
        src14 <= 12'h715;
        src15 <= 12'he83;
        src16 <= 12'h53c;
        src17 <= 12'h71e;
        src18 <= 12'h79a;
        src19 <= 12'h443;
        src20 <= 12'h726;
        src21 <= 12'h456;
        src22 <= 12'hc34;
        src23 <= 12'hc15;
        src24 <= 12'h186;
        src25 <= 12'hb21;
        src26 <= 12'h43b;
        src27 <= 12'h197;
        src28 <= 12'h5be;
        src29 <= 12'hdb2;
        src30 <= 12'ha84;
        src31 <= 12'h382;
        exp <= 17'hebb9;
        #1
        src0 <= 12'h2d3;
        src1 <= 12'h5cb;
        src2 <= 12'h5cb;
        src3 <= 12'h7c6;
        src4 <= 12'h51e;
        src5 <= 12'h7de;
        src6 <= 12'hac2;
        src7 <= 12'hf41;
        src8 <= 12'h78b;
        src9 <= 12'hec2;
        src10 <= 12'h15;
        src11 <= 12'ha1e;
        src12 <= 12'h935;
        src13 <= 12'h80e;
        src14 <= 12'hc40;
        src15 <= 12'hfdb;
        src16 <= 12'hb36;
        src17 <= 12'ha38;
        src18 <= 12'h1d3;
        src19 <= 12'he9c;
        src20 <= 12'h6f8;
        src21 <= 12'h245;
        src22 <= 12'h1d2;
        src23 <= 12'h78;
        src24 <= 12'h48e;
        src25 <= 12'h9cc;
        src26 <= 12'h302;
        src27 <= 12'h83;
        src28 <= 12'h8aa;
        src29 <= 12'h5ee;
        src30 <= 12'ha07;
        src31 <= 12'h340;
        exp <= 17'hea2e;
        #1
        src0 <= 12'he45;
        src1 <= 12'hb40;
        src2 <= 12'h75f;
        src3 <= 12'hfae;
        src4 <= 12'h23e;
        src5 <= 12'hdb4;
        src6 <= 12'h795;
        src7 <= 12'h9ac;
        src8 <= 12'h2e8;
        src9 <= 12'ha68;
        src10 <= 12'h7d9;
        src11 <= 12'h387;
        src12 <= 12'h312;
        src13 <= 12'h7fc;
        src14 <= 12'hc21;
        src15 <= 12'hb7d;
        src16 <= 12'h68;
        src17 <= 12'h2e9;
        src18 <= 12'hcf1;
        src19 <= 12'hcaa;
        src20 <= 12'h383;
        src21 <= 12'hf02;
        src22 <= 12'h236;
        src23 <= 12'h858;
        src24 <= 12'h748;
        src25 <= 12'h8cf;
        src26 <= 12'hda;
        src27 <= 12'haaf;
        src28 <= 12'h547;
        src29 <= 12'h26b;
        src30 <= 12'h6a2;
        src31 <= 12'h140;
        exp <= 17'hf254;
        #1
        src0 <= 12'h6ef;
        src1 <= 12'hae8;
        src2 <= 12'hf68;
        src3 <= 12'hdd5;
        src4 <= 12'h7d7;
        src5 <= 12'hca;
        src6 <= 12'h7e7;
        src7 <= 12'h3a8;
        src8 <= 12'hd7f;
        src9 <= 12'hf8b;
        src10 <= 12'hc2e;
        src11 <= 12'heb6;
        src12 <= 12'h6c7;
        src13 <= 12'h665;
        src14 <= 12'hadb;
        src15 <= 12'hcc7;
        src16 <= 12'hf74;
        src17 <= 12'h58b;
        src18 <= 12'h83f;
        src19 <= 12'h452;
        src20 <= 12'h203;
        src21 <= 12'hf5e;
        src22 <= 12'h115;
        src23 <= 12'h464;
        src24 <= 12'h354;
        src25 <= 12'h1c7;
        src26 <= 12'hde9;
        src27 <= 12'h4f1;
        src28 <= 12'h1cb;
        src29 <= 12'hda1;
        src30 <= 12'hd6b;
        src31 <= 12'h2c2;
        exp <= 17'h10ff8;
        #1
        src0 <= 12'hcf1;
        src1 <= 12'h664;
        src2 <= 12'hca8;
        src3 <= 12'h657;
        src4 <= 12'hbd;
        src5 <= 12'h7b9;
        src6 <= 12'h360;
        src7 <= 12'hb69;
        src8 <= 12'h14;
        src9 <= 12'h592;
        src10 <= 12'hb31;
        src11 <= 12'h24c;
        src12 <= 12'h556;
        src13 <= 12'hd5a;
        src14 <= 12'h513;
        src15 <= 12'ha93;
        src16 <= 12'h764;
        src17 <= 12'h630;
        src18 <= 12'h786;
        src19 <= 12'he83;
        src20 <= 12'he47;
        src21 <= 12'hb72;
        src22 <= 12'h129;
        src23 <= 12'hdb;
        src24 <= 12'h4d8;
        src25 <= 12'hee5;
        src26 <= 12'hd42;
        src27 <= 12'h92a;
        src28 <= 12'h8fa;
        src29 <= 12'h662;
        src30 <= 12'h264;
        src31 <= 12'h7b0;
        exp <= 17'hf5ff;
        #1
        src0 <= 12'hc6a;
        src1 <= 12'h26d;
        src2 <= 12'h829;
        src3 <= 12'h3a5;
        src4 <= 12'hbe0;
        src5 <= 12'hdf0;
        src6 <= 12'ha06;
        src7 <= 12'h990;
        src8 <= 12'h593;
        src9 <= 12'hc0f;
        src10 <= 12'h648;
        src11 <= 12'h457;
        src12 <= 12'h665;
        src13 <= 12'he4c;
        src14 <= 12'h40d;
        src15 <= 12'h824;
        src16 <= 12'h85f;
        src17 <= 12'ha5f;
        src18 <= 12'h35e;
        src19 <= 12'ha35;
        src20 <= 12'hc73;
        src21 <= 12'ha8f;
        src22 <= 12'h8f1;
        src23 <= 12'hbc1;
        src24 <= 12'hbc;
        src25 <= 12'h34b;
        src26 <= 12'h48f;
        src27 <= 12'h94f;
        src28 <= 12'h8a8;
        src29 <= 12'h8da;
        src30 <= 12'h3f0;
        src31 <= 12'hb20;
        exp <= 17'h103aa;
        #1
        src0 <= 12'haa0;
        src1 <= 12'h788;
        src2 <= 12'hb5b;
        src3 <= 12'h4d7;
        src4 <= 12'h2a9;
        src5 <= 12'h2a1;
        src6 <= 12'h728;
        src7 <= 12'h278;
        src8 <= 12'ha82;
        src9 <= 12'h439;
        src10 <= 12'h257;
        src11 <= 12'h4c9;
        src12 <= 12'ha19;
        src13 <= 12'h512;
        src14 <= 12'h8d1;
        src15 <= 12'hbdc;
        src16 <= 12'h171;
        src17 <= 12'h705;
        src18 <= 12'hbc1;
        src19 <= 12'h4b0;
        src20 <= 12'he4a;
        src21 <= 12'h787;
        src22 <= 12'h378;
        src23 <= 12'h48;
        src24 <= 12'hc4;
        src25 <= 12'hc69;
        src26 <= 12'h649;
        src27 <= 12'hc4f;
        src28 <= 12'h8fb;
        src29 <= 12'h85a;
        src30 <= 12'h5b3;
        src31 <= 12'hb3;
        exp <= 17'hd4ef;
        #1
        src0 <= 12'h946;
        src1 <= 12'hffd;
        src2 <= 12'h281;
        src3 <= 12'hf9;
        src4 <= 12'he21;
        src5 <= 12'hd79;
        src6 <= 12'h5fc;
        src7 <= 12'hc3f;
        src8 <= 12'h530;
        src9 <= 12'he8e;
        src10 <= 12'he09;
        src11 <= 12'h8cb;
        src12 <= 12'h9b9;
        src13 <= 12'hc47;
        src14 <= 12'h7ce;
        src15 <= 12'h76;
        src16 <= 12'he66;
        src17 <= 12'h486;
        src18 <= 12'h121;
        src19 <= 12'hc6e;
        src20 <= 12'h4d5;
        src21 <= 12'hf16;
        src22 <= 12'hdf;
        src23 <= 12'h9ee;
        src24 <= 12'h75a;
        src25 <= 12'hb28;
        src26 <= 12'h5be;
        src27 <= 12'h5b7;
        src28 <= 12'h20b;
        src29 <= 12'h13c;
        src30 <= 12'h53b;
        src31 <= 12'h778;
        exp <= 17'h1008c;
        #1
        src0 <= 12'h8bf;
        src1 <= 12'h7c4;
        src2 <= 12'h191;
        src3 <= 12'h7cf;
        src4 <= 12'h3ec;
        src5 <= 12'h37d;
        src6 <= 12'hfe9;
        src7 <= 12'hfb2;
        src8 <= 12'h285;
        src9 <= 12'hda7;
        src10 <= 12'hfd4;
        src11 <= 12'hf77;
        src12 <= 12'h539;
        src13 <= 12'hf2c;
        src14 <= 12'h77;
        src15 <= 12'hc1f;
        src16 <= 12'h9b2;
        src17 <= 12'h327;
        src18 <= 12'h48e;
        src19 <= 12'hfd3;
        src20 <= 12'h3c9;
        src21 <= 12'hf49;
        src22 <= 12'h25c;
        src23 <= 12'hb63;
        src24 <= 12'he63;
        src25 <= 12'haab;
        src26 <= 12'hdfa;
        src27 <= 12'h499;
        src28 <= 12'hb37;
        src29 <= 12'h2a2;
        src30 <= 12'h254;
        src31 <= 12'h9c8;
        exp <= 17'h118fa;
        #1
        src0 <= 12'h3e0;
        src1 <= 12'hbfa;
        src2 <= 12'he60;
        src3 <= 12'h87a;
        src4 <= 12'h1bc;
        src5 <= 12'h9fe;
        src6 <= 12'h59b;
        src7 <= 12'h6f3;
        src8 <= 12'h5a2;
        src9 <= 12'h2dd;
        src10 <= 12'hfd3;
        src11 <= 12'h290;
        src12 <= 12'hc5f;
        src13 <= 12'hc34;
        src14 <= 12'h408;
        src15 <= 12'he63;
        src16 <= 12'h854;
        src17 <= 12'h987;
        src18 <= 12'h3a8;
        src19 <= 12'ha6c;
        src20 <= 12'h71b;
        src21 <= 12'hfca;
        src22 <= 12'h4b0;
        src23 <= 12'hbad;
        src24 <= 12'h495;
        src25 <= 12'h5cd;
        src26 <= 12'h42c;
        src27 <= 12'h8bf;
        src28 <= 12'h572;
        src29 <= 12'h397;
        src30 <= 12'h5b1;
        src31 <= 12'hd11;
        exp <= 17'hff25;
        #1
        src0 <= 12'h732;
        src1 <= 12'haeb;
        src2 <= 12'h90;
        src3 <= 12'h7a4;
        src4 <= 12'h9b9;
        src5 <= 12'had0;
        src6 <= 12'h119;
        src7 <= 12'h922;
        src8 <= 12'hd51;
        src9 <= 12'hf4e;
        src10 <= 12'h5ba;
        src11 <= 12'hb9c;
        src12 <= 12'h98f;
        src13 <= 12'h26;
        src14 <= 12'hef8;
        src15 <= 12'h140;
        src16 <= 12'hd7b;
        src17 <= 12'hcb2;
        src18 <= 12'hc3f;
        src19 <= 12'h848;
        src20 <= 12'h15e;
        src21 <= 12'hbb2;
        src22 <= 12'hca9;
        src23 <= 12'h30c;
        src24 <= 12'h1ee;
        src25 <= 12'ha0d;
        src26 <= 12'h371;
        src27 <= 12'hd5c;
        src28 <= 12'hdf;
        src29 <= 12'hfb;
        src30 <= 12'hdcf;
        src31 <= 12'hd1a;
        exp <= 17'h105fb;
        #1
        src0 <= 12'h9fa;
        src1 <= 12'h495;
        src2 <= 12'h2b2;
        src3 <= 12'h383;
        src4 <= 12'h82d;
        src5 <= 12'h110;
        src6 <= 12'h9e2;
        src7 <= 12'hf41;
        src8 <= 12'hf9d;
        src9 <= 12'h9b4;
        src10 <= 12'h85a;
        src11 <= 12'h23e;
        src12 <= 12'h290;
        src13 <= 12'h1ff;
        src14 <= 12'hdb6;
        src15 <= 12'hfb2;
        src16 <= 12'ha1a;
        src17 <= 12'hbc3;
        src18 <= 12'h1b9;
        src19 <= 12'hbf2;
        src20 <= 12'h62c;
        src21 <= 12'hb41;
        src22 <= 12'he29;
        src23 <= 12'h4f5;
        src24 <= 12'hf0f;
        src25 <= 12'hbad;
        src26 <= 12'hc32;
        src27 <= 12'h82a;
        src28 <= 12'h1cf;
        src29 <= 12'hcbf;
        src30 <= 12'hd3b;
        src31 <= 12'hf9;
        exp <= 17'h110f1;
        #1
        src0 <= 12'h7da;
        src1 <= 12'hf6a;
        src2 <= 12'h510;
        src3 <= 12'h1e3;
        src4 <= 12'h30;
        src5 <= 12'h59f;
        src6 <= 12'hb4;
        src7 <= 12'h308;
        src8 <= 12'hc10;
        src9 <= 12'h4bd;
        src10 <= 12'hc7;
        src11 <= 12'hbcb;
        src12 <= 12'h474;
        src13 <= 12'hccb;
        src14 <= 12'hacc;
        src15 <= 12'haeb;
        src16 <= 12'hbe8;
        src17 <= 12'h4d;
        src18 <= 12'h4a9;
        src19 <= 12'h177;
        src20 <= 12'h9df;
        src21 <= 12'he34;
        src22 <= 12'hd9e;
        src23 <= 12'hddf;
        src24 <= 12'hd03;
        src25 <= 12'hd61;
        src26 <= 12'h8b4;
        src27 <= 12'h2d1;
        src28 <= 12'h4eb;
        src29 <= 12'hc62;
        src30 <= 12'h175;
        src31 <= 12'hf6f;
        exp <= 17'hfa16;
        #1
        src0 <= 12'h4d1;
        src1 <= 12'h1;
        src2 <= 12'hfee;
        src3 <= 12'hd09;
        src4 <= 12'ha8d;
        src5 <= 12'hc51;
        src6 <= 12'hb79;
        src7 <= 12'ha54;
        src8 <= 12'h2a4;
        src9 <= 12'he15;
        src10 <= 12'h496;
        src11 <= 12'h8d5;
        src12 <= 12'hc9d;
        src13 <= 12'hdf4;
        src14 <= 12'h180;
        src15 <= 12'h63f;
        src16 <= 12'h142;
        src17 <= 12'he25;
        src18 <= 12'hff0;
        src19 <= 12'h7f9;
        src20 <= 12'had3;
        src21 <= 12'h157;
        src22 <= 12'he2f;
        src23 <= 12'hc04;
        src24 <= 12'h6ba;
        src25 <= 12'h995;
        src26 <= 12'h863;
        src27 <= 12'h7ce;
        src28 <= 12'hbcf;
        src29 <= 12'hbea;
        src30 <= 12'h64d;
        src31 <= 12'h69c;
        exp <= 17'h121b7;
        #1
        src0 <= 12'ha1;
        src1 <= 12'h98c;
        src2 <= 12'h7a1;
        src3 <= 12'h397;
        src4 <= 12'he4c;
        src5 <= 12'hae3;
        src6 <= 12'hd59;
        src7 <= 12'ha56;
        src8 <= 12'h5d0;
        src9 <= 12'h5b4;
        src10 <= 12'he79;
        src11 <= 12'h516;
        src12 <= 12'hab9;
        src13 <= 12'hb4f;
        src14 <= 12'h49d;
        src15 <= 12'hc85;
        src16 <= 12'hc3;
        src17 <= 12'h993;
        src18 <= 12'h555;
        src19 <= 12'h7a7;
        src20 <= 12'h985;
        src21 <= 12'hb10;
        src22 <= 12'ha97;
        src23 <= 12'h88;
        src24 <= 12'hbae;
        src25 <= 12'h5d2;
        src26 <= 12'hbc9;
        src27 <= 12'hcc7;
        src28 <= 12'hee0;
        src29 <= 12'h5a5;
        src30 <= 12'h17f;
        src31 <= 12'h134;
        exp <= 17'h104ce;
        #1
        src0 <= 12'he0;
        src1 <= 12'he75;
        src2 <= 12'h4bb;
        src3 <= 12'h833;
        src4 <= 12'hb1;
        src5 <= 12'h714;
        src6 <= 12'h88f;
        src7 <= 12'hb02;
        src8 <= 12'hadc;
        src9 <= 12'h5ec;
        src10 <= 12'h8e6;
        src11 <= 12'h197;
        src12 <= 12'h943;
        src13 <= 12'h7ba;
        src14 <= 12'h5fd;
        src15 <= 12'h7a5;
        src16 <= 12'hadc;
        src17 <= 12'h848;
        src18 <= 12'h2ec;
        src19 <= 12'hd76;
        src20 <= 12'h748;
        src21 <= 12'h45f;
        src22 <= 12'hd22;
        src23 <= 12'h8b4;
        src24 <= 12'h9bb;
        src25 <= 12'h9ab;
        src26 <= 12'h227;
        src27 <= 12'h50e;
        src28 <= 12'h31;
        src29 <= 12'h2bf;
        src30 <= 12'h1e3;
        src31 <= 12'hcfa;
        exp <= 17'he2e8;
        #1
        src0 <= 12'hc1a;
        src1 <= 12'h719;
        src2 <= 12'hfe1;
        src3 <= 12'ha94;
        src4 <= 12'h4ae;
        src5 <= 12'h200;
        src6 <= 12'h1b7;
        src7 <= 12'h1ed;
        src8 <= 12'hfca;
        src9 <= 12'hea5;
        src10 <= 12'h53f;
        src11 <= 12'h894;
        src12 <= 12'hf7a;
        src13 <= 12'h3a4;
        src14 <= 12'h514;
        src15 <= 12'h28d;
        src16 <= 12'h7e7;
        src17 <= 12'h581;
        src18 <= 12'h4a3;
        src19 <= 12'hced;
        src20 <= 12'hdde;
        src21 <= 12'h40c;
        src22 <= 12'h28c;
        src23 <= 12'hcb1;
        src24 <= 12'h2a0;
        src25 <= 12'hfa5;
        src26 <= 12'hf21;
        src27 <= 12'h151;
        src28 <= 12'hff4;
        src29 <= 12'h550;
        src30 <= 12'h306;
        src31 <= 12'h7c0;
        exp <= 17'h101db;
        #1
        src0 <= 12'h8fe;
        src1 <= 12'ha8;
        src2 <= 12'h9c8;
        src3 <= 12'hd79;
        src4 <= 12'ha5c;
        src5 <= 12'h1b8;
        src6 <= 12'hf7e;
        src7 <= 12'h91d;
        src8 <= 12'h8a8;
        src9 <= 12'ha49;
        src10 <= 12'h45b;
        src11 <= 12'h70c;
        src12 <= 12'hb87;
        src13 <= 12'hac5;
        src14 <= 12'h13d;
        src15 <= 12'hc9e;
        src16 <= 12'h53d;
        src17 <= 12'h273;
        src18 <= 12'hac8;
        src19 <= 12'hc4d;
        src20 <= 12'hc88;
        src21 <= 12'h1d4;
        src22 <= 12'hf77;
        src23 <= 12'ha2a;
        src24 <= 12'h860;
        src25 <= 12'h403;
        src26 <= 12'h2ed;
        src27 <= 12'h690;
        src28 <= 12'h276;
        src29 <= 12'h485;
        src30 <= 12'hc95;
        src31 <= 12'hb1e;
        exp <= 17'h10365;
        #1
        src0 <= 12'h5c8;
        src1 <= 12'h75;
        src2 <= 12'h2af;
        src3 <= 12'h11d;
        src4 <= 12'h91a;
        src5 <= 12'hbe4;
        src6 <= 12'h45a;
        src7 <= 12'hd15;
        src8 <= 12'hf07;
        src9 <= 12'h652;
        src10 <= 12'hd9e;
        src11 <= 12'h1dc;
        src12 <= 12'hbcf;
        src13 <= 12'ha8a;
        src14 <= 12'h40c;
        src15 <= 12'hebc;
        src16 <= 12'h42f;
        src17 <= 12'hc03;
        src18 <= 12'hf6b;
        src19 <= 12'h10e;
        src20 <= 12'h6ec;
        src21 <= 12'hdb1;
        src22 <= 12'hdf8;
        src23 <= 12'h7;
        src24 <= 12'haa3;
        src25 <= 12'h5b5;
        src26 <= 12'h111;
        src27 <= 12'hfe9;
        src28 <= 12'h2f5;
        src29 <= 12'ha16;
        src30 <= 12'he04;
        src31 <= 12'h168;
        exp <= 17'hff7a;
        #1
        src0 <= 12'hacf;
        src1 <= 12'h268;
        src2 <= 12'ha51;
        src3 <= 12'he98;
        src4 <= 12'hd25;
        src5 <= 12'ha46;
        src6 <= 12'h71a;
        src7 <= 12'h82a;
        src8 <= 12'hdcf;
        src9 <= 12'ha16;
        src10 <= 12'h9c4;
        src11 <= 12'h22a;
        src12 <= 12'h967;
        src13 <= 12'h7f6;
        src14 <= 12'h3e7;
        src15 <= 12'ha0b;
        src16 <= 12'hc40;
        src17 <= 12'hdba;
        src18 <= 12'h2c2;
        src19 <= 12'h631;
        src20 <= 12'h8aa;
        src21 <= 12'hdce;
        src22 <= 12'h8d;
        src23 <= 12'ha1f;
        src24 <= 12'h1ea;
        src25 <= 12'h63a;
        src26 <= 12'h392;
        src27 <= 12'ha04;
        src28 <= 12'h886;
        src29 <= 12'ha67;
        src30 <= 12'hbd9;
        src31 <= 12'h72f;
        exp <= 17'h10fb1;
        #1
        src0 <= 12'h1a4;
        src1 <= 12'he3b;
        src2 <= 12'h48a;
        src3 <= 12'heef;
        src4 <= 12'hd57;
        src5 <= 12'haf7;
        src6 <= 12'hd1a;
        src7 <= 12'h8ab;
        src8 <= 12'ha5a;
        src9 <= 12'h83e;
        src10 <= 12'h158;
        src11 <= 12'hfd7;
        src12 <= 12'h257;
        src13 <= 12'h26b;
        src14 <= 12'h6b2;
        src15 <= 12'ha47;
        src16 <= 12'h38c;
        src17 <= 12'h8ab;
        src18 <= 12'hdb3;
        src19 <= 12'h239;
        src20 <= 12'hd3a;
        src21 <= 12'h9d3;
        src22 <= 12'ha4d;
        src23 <= 12'h8e8;
        src24 <= 12'h7ef;
        src25 <= 12'hde;
        src26 <= 12'he3d;
        src27 <= 12'h506;
        src28 <= 12'h142;
        src29 <= 12'h40;
        src30 <= 12'h302;
        src31 <= 12'h78a;
        exp <= 17'hf970;
        #1
        src0 <= 12'h231;
        src1 <= 12'ha9c;
        src2 <= 12'hfa5;
        src3 <= 12'h8e9;
        src4 <= 12'h2d8;
        src5 <= 12'h4f7;
        src6 <= 12'he4b;
        src7 <= 12'hfe0;
        src8 <= 12'h682;
        src9 <= 12'h233;
        src10 <= 12'h83b;
        src11 <= 12'h41f;
        src12 <= 12'hcce;
        src13 <= 12'h426;
        src14 <= 12'hc88;
        src15 <= 12'h9ee;
        src16 <= 12'h18b;
        src17 <= 12'ha96;
        src18 <= 12'h602;
        src19 <= 12'h418;
        src20 <= 12'ha69;
        src21 <= 12'h14d;
        src22 <= 12'h6f8;
        src23 <= 12'h60c;
        src24 <= 12'h774;
        src25 <= 12'hae9;
        src26 <= 12'h18f;
        src27 <= 12'he60;
        src28 <= 12'h295;
        src29 <= 12'h5fd;
        src30 <= 12'h909;
        src31 <= 12'hf94;
        exp <= 17'hfa3e;
        #1
        src0 <= 12'h49;
        src1 <= 12'hadc;
        src2 <= 12'heb3;
        src3 <= 12'h53c;
        src4 <= 12'h9be;
        src5 <= 12'h63e;
        src6 <= 12'hf3c;
        src7 <= 12'h6d4;
        src8 <= 12'hd6f;
        src9 <= 12'h968;
        src10 <= 12'h63d;
        src11 <= 12'h8b5;
        src12 <= 12'h39a;
        src13 <= 12'h1e3;
        src14 <= 12'ha27;
        src15 <= 12'hbcd;
        src16 <= 12'h105;
        src17 <= 12'h24f;
        src18 <= 12'h272;
        src19 <= 12'h159;
        src20 <= 12'h634;
        src21 <= 12'h376;
        src22 <= 12'hd7c;
        src23 <= 12'h973;
        src24 <= 12'hcec;
        src25 <= 12'hf78;
        src26 <= 12'ha92;
        src27 <= 12'h559;
        src28 <= 12'ha77;
        src29 <= 12'h3e5;
        src30 <= 12'h63d;
        src31 <= 12'hcab;
        exp <= 17'hfba5;
        #1
        src0 <= 12'h8e9;
        src1 <= 12'hb71;
        src2 <= 12'h3c2;
        src3 <= 12'ha2f;
        src4 <= 12'h286;
        src5 <= 12'he0d;
        src6 <= 12'h96d;
        src7 <= 12'h73;
        src8 <= 12'hc03;
        src9 <= 12'h6e3;
        src10 <= 12'he82;
        src11 <= 12'hd36;
        src12 <= 12'h22d;
        src13 <= 12'h554;
        src14 <= 12'hc37;
        src15 <= 12'hb90;
        src16 <= 12'heec;
        src17 <= 12'hbcf;
        src18 <= 12'hac3;
        src19 <= 12'hb3d;
        src20 <= 12'h3ca;
        src21 <= 12'heb8;
        src22 <= 12'he5a;
        src23 <= 12'h595;
        src24 <= 12'h34d;
        src25 <= 12'hd5e;
        src26 <= 12'hbf8;
        src27 <= 12'h598;
        src28 <= 12'hbb5;
        src29 <= 12'hd76;
        src30 <= 12'hc53;
        src31 <= 12'h84a;
        exp <= 17'h131d3;
        #1
        src0 <= 12'ha1a;
        src1 <= 12'h1b0;
        src2 <= 12'h100;
        src3 <= 12'h6af;
        src4 <= 12'h7f2;
        src5 <= 12'hec3;
        src6 <= 12'hc52;
        src7 <= 12'h38f;
        src8 <= 12'he55;
        src9 <= 12'haff;
        src10 <= 12'ha0d;
        src11 <= 12'h151;
        src12 <= 12'h3;
        src13 <= 12'h778;
        src14 <= 12'hd55;
        src15 <= 12'hcca;
        src16 <= 12'h6b;
        src17 <= 12'hfdc;
        src18 <= 12'hd15;
        src19 <= 12'h576;
        src20 <= 12'h89a;
        src21 <= 12'h1e3;
        src22 <= 12'h884;
        src23 <= 12'h3d4;
        src24 <= 12'hd90;
        src25 <= 12'h373;
        src26 <= 12'h971;
        src27 <= 12'h755;
        src28 <= 12'h86;
        src29 <= 12'hb3c;
        src30 <= 12'h3e0;
        src31 <= 12'h84;
        exp <= 17'hebf1;
        #1
        src0 <= 12'hbf3;
        src1 <= 12'h154;
        src2 <= 12'ha4d;
        src3 <= 12'h3fb;
        src4 <= 12'hdb8;
        src5 <= 12'he43;
        src6 <= 12'hf8f;
        src7 <= 12'h1a4;
        src8 <= 12'h98d;
        src9 <= 12'h3fc;
        src10 <= 12'ha8f;
        src11 <= 12'h681;
        src12 <= 12'h21a;
        src13 <= 12'h941;
        src14 <= 12'h912;
        src15 <= 12'h5c2;
        src16 <= 12'h157;
        src17 <= 12'he1b;
        src18 <= 12'hde;
        src19 <= 12'hd8a;
        src20 <= 12'h993;
        src21 <= 12'hae1;
        src22 <= 12'h72d;
        src23 <= 12'h4a4;
        src24 <= 12'h518;
        src25 <= 12'h8f6;
        src26 <= 12'h1d5;
        src27 <= 12'h4a0;
        src28 <= 12'h5c1;
        src29 <= 12'h645;
        src30 <= 12'h466;
        src31 <= 12'h260;
        exp <= 17'he6f3;
        #1
        src0 <= 12'h9fc;
        src1 <= 12'h81b;
        src2 <= 12'hf95;
        src3 <= 12'h62b;
        src4 <= 12'h6ed;
        src5 <= 12'hbf;
        src6 <= 12'h51;
        src7 <= 12'he40;
        src8 <= 12'hb81;
        src9 <= 12'h939;
        src10 <= 12'h78b;
        src11 <= 12'hf88;
        src12 <= 12'h8de;
        src13 <= 12'hdbc;
        src14 <= 12'h555;
        src15 <= 12'h1db;
        src16 <= 12'h126;
        src17 <= 12'h6f9;
        src18 <= 12'hcb2;
        src19 <= 12'h3a4;
        src20 <= 12'hd11;
        src21 <= 12'h4c5;
        src22 <= 12'h119;
        src23 <= 12'h14;
        src24 <= 12'h9f0;
        src25 <= 12'h5b2;
        src26 <= 12'hf1c;
        src27 <= 12'h475;
        src28 <= 12'h85c;
        src29 <= 12'h565;
        src30 <= 12'h7e6;
        src31 <= 12'h2ff;
        exp <= 17'heefc;
        #1
        src0 <= 12'h55;
        src1 <= 12'h47c;
        src2 <= 12'h6e7;
        src3 <= 12'h8c7;
        src4 <= 12'h37a;
        src5 <= 12'he34;
        src6 <= 12'h85;
        src7 <= 12'h676;
        src8 <= 12'hdd1;
        src9 <= 12'hfc9;
        src10 <= 12'hf4a;
        src11 <= 12'hcf1;
        src12 <= 12'had1;
        src13 <= 12'h7;
        src14 <= 12'h693;
        src15 <= 12'h408;
        src16 <= 12'h32f;
        src17 <= 12'h579;
        src18 <= 12'hae;
        src19 <= 12'h16a;
        src20 <= 12'hf44;
        src21 <= 12'h607;
        src22 <= 12'h274;
        src23 <= 12'haed;
        src24 <= 12'h243;
        src25 <= 12'h93e;
        src26 <= 12'h563;
        src27 <= 12'hf8a;
        src28 <= 12'h50d;
        src29 <= 12'h3e3;
        src30 <= 12'hc9e;
        src31 <= 12'h7c8;
        exp <= 17'he7a0;
        #1
        src0 <= 12'h849;
        src1 <= 12'h5e3;
        src2 <= 12'h230;
        src3 <= 12'hec7;
        src4 <= 12'hf34;
        src5 <= 12'h764;
        src6 <= 12'h31;
        src7 <= 12'h9db;
        src8 <= 12'hdf5;
        src9 <= 12'h10f;
        src10 <= 12'h37c;
        src11 <= 12'h584;
        src12 <= 12'h3c1;
        src13 <= 12'h2c4;
        src14 <= 12'h362;
        src15 <= 12'haca;
        src16 <= 12'hf54;
        src17 <= 12'h96a;
        src18 <= 12'hf8f;
        src19 <= 12'hb79;
        src20 <= 12'h33;
        src21 <= 12'he78;
        src22 <= 12'h7f3;
        src23 <= 12'h4c;
        src24 <= 12'h44c;
        src25 <= 12'h343;
        src26 <= 12'h9b4;
        src27 <= 12'h1e;
        src28 <= 12'h13e;
        src29 <= 12'h42c;
        src30 <= 12'h8df;
        src31 <= 12'h465;
        exp <= 17'hdb3b;
        #1
        src0 <= 12'h514;
        src1 <= 12'hf84;
        src2 <= 12'hb7b;
        src3 <= 12'hab8;
        src4 <= 12'h42c;
        src5 <= 12'h73;
        src6 <= 12'h697;
        src7 <= 12'h3d3;
        src8 <= 12'h8cb;
        src9 <= 12'hce;
        src10 <= 12'hc30;
        src11 <= 12'hacb;
        src12 <= 12'h1c7;
        src13 <= 12'h224;
        src14 <= 12'he03;
        src15 <= 12'h6f1;
        src16 <= 12'hee0;
        src17 <= 12'h3a3;
        src18 <= 12'hf5d;
        src19 <= 12'hb82;
        src20 <= 12'he19;
        src21 <= 12'h313;
        src22 <= 12'hfe9;
        src23 <= 12'h631;
        src24 <= 12'h55e;
        src25 <= 12'h4e4;
        src26 <= 12'h9d7;
        src27 <= 12'hce4;
        src28 <= 12'h5db;
        src29 <= 12'h423;
        src30 <= 12'h430;
        src31 <= 12'h461;
        exp <= 17'hfb7b;
        #1
        src0 <= 12'h409;
        src1 <= 12'h64b;
        src2 <= 12'h63a;
        src3 <= 12'ha73;
        src4 <= 12'h6e0;
        src5 <= 12'h8d0;
        src6 <= 12'h7d1;
        src7 <= 12'ha23;
        src8 <= 12'h306;
        src9 <= 12'h261;
        src10 <= 12'h921;
        src11 <= 12'h89e;
        src12 <= 12'h5d0;
        src13 <= 12'h27e;
        src14 <= 12'he19;
        src15 <= 12'h41a;
        src16 <= 12'h208;
        src17 <= 12'ha0e;
        src18 <= 12'h7d1;
        src19 <= 12'h208;
        src20 <= 12'h335;
        src21 <= 12'h8f6;
        src22 <= 12'hde9;
        src23 <= 12'h2fd;
        src24 <= 12'h1e8;
        src25 <= 12'h704;
        src26 <= 12'h901;
        src27 <= 12'h542;
        src28 <= 12'h9e6;
        src29 <= 12'h3b;
        src30 <= 12'hffa;
        src31 <= 12'h9b;
        exp <= 17'hd331;
        #1
        src0 <= 12'h62e;
        src1 <= 12'h803;
        src2 <= 12'h7c1;
        src3 <= 12'h8c3;
        src4 <= 12'h50b;
        src5 <= 12'hd7a;
        src6 <= 12'ha77;
        src7 <= 12'h8f8;
        src8 <= 12'h7cb;
        src9 <= 12'h588;
        src10 <= 12'h82b;
        src11 <= 12'hbfe;
        src12 <= 12'hafa;
        src13 <= 12'h2a6;
        src14 <= 12'h528;
        src15 <= 12'h60d;
        src16 <= 12'h7a9;
        src17 <= 12'hf12;
        src18 <= 12'h6f3;
        src19 <= 12'hb5f;
        src20 <= 12'h81;
        src21 <= 12'h635;
        src22 <= 12'h138;
        src23 <= 12'he8a;
        src24 <= 12'h1ed;
        src25 <= 12'h2f5;
        src26 <= 12'h2b7;
        src27 <= 12'h591;
        src28 <= 12'h7cb;
        src29 <= 12'hab9;
        src30 <= 12'h346;
        src31 <= 12'h265;
        exp <= 17'he3d8;
        #1
        src0 <= 12'h99a;
        src1 <= 12'h816;
        src2 <= 12'h8de;
        src3 <= 12'he4;
        src4 <= 12'had1;
        src5 <= 12'h26c;
        src6 <= 12'h37f;
        src7 <= 12'h41a;
        src8 <= 12'h7ac;
        src9 <= 12'h758;
        src10 <= 12'h42f;
        src11 <= 12'hd8a;
        src12 <= 12'h954;
        src13 <= 12'h5da;
        src14 <= 12'ha90;
        src15 <= 12'ha87;
        src16 <= 12'h9c0;
        src17 <= 12'hb59;
        src18 <= 12'he00;
        src19 <= 12'h175;
        src20 <= 12'h825;
        src21 <= 12'habe;
        src22 <= 12'h8f1;
        src23 <= 12'hb73;
        src24 <= 12'h8ec;
        src25 <= 12'h124;
        src26 <= 12'hec;
        src27 <= 12'h929;
        src28 <= 12'hc40;
        src29 <= 12'h13b;
        src30 <= 12'h9f6;
        src31 <= 12'h6ec;
        exp <= 17'hf3a1;
        #1
        src0 <= 12'h3e6;
        src1 <= 12'h753;
        src2 <= 12'h8c9;
        src3 <= 12'h30b;
        src4 <= 12'h436;
        src5 <= 12'h365;
        src6 <= 12'hcc6;
        src7 <= 12'h505;
        src8 <= 12'h428;
        src9 <= 12'h9be;
        src10 <= 12'hf82;
        src11 <= 12'h701;
        src12 <= 12'hca9;
        src13 <= 12'hb63;
        src14 <= 12'hab5;
        src15 <= 12'hc2b;
        src16 <= 12'h868;
        src17 <= 12'h1cb;
        src18 <= 12'h176;
        src19 <= 12'hfeb;
        src20 <= 12'h9e3;
        src21 <= 12'h98a;
        src22 <= 12'h475;
        src23 <= 12'h62c;
        src24 <= 12'hb42;
        src25 <= 12'h875;
        src26 <= 12'h328;
        src27 <= 12'h29b;
        src28 <= 12'hd21;
        src29 <= 12'he96;
        src30 <= 12'h974;
        src31 <= 12'h3be;
        exp <= 17'hffcd;
        #1
        src0 <= 12'h4e4;
        src1 <= 12'h651;
        src2 <= 12'hd38;
        src3 <= 12'h3e9;
        src4 <= 12'h2ce;
        src5 <= 12'hef0;
        src6 <= 12'hf86;
        src7 <= 12'hfc5;
        src8 <= 12'hcef;
        src9 <= 12'h766;
        src10 <= 12'hb52;
        src11 <= 12'h18b;
        src12 <= 12'hbe9;
        src13 <= 12'h946;
        src14 <= 12'h7f2;
        src15 <= 12'hbba;
        src16 <= 12'h65e;
        src17 <= 12'h261;
        src18 <= 12'h358;
        src19 <= 12'h727;
        src20 <= 12'ha56;
        src21 <= 12'hca;
        src22 <= 12'h91b;
        src23 <= 12'hb51;
        src24 <= 12'hec8;
        src25 <= 12'h500;
        src26 <= 12'hfdf;
        src27 <= 12'h811;
        src28 <= 12'h52c;
        src29 <= 12'hcb7;
        src30 <= 12'h4d4;
        src31 <= 12'h7e2;
        exp <= 17'h11487;
        #1
        src0 <= 12'hb6e;
        src1 <= 12'h8b4;
        src2 <= 12'h21b;
        src3 <= 12'hbc9;
        src4 <= 12'h68d;
        src5 <= 12'hf07;
        src6 <= 12'h884;
        src7 <= 12'h187;
        src8 <= 12'h613;
        src9 <= 12'h448;
        src10 <= 12'hd9b;
        src11 <= 12'h500;
        src12 <= 12'h213;
        src13 <= 12'h77e;
        src14 <= 12'h755;
        src15 <= 12'h43d;
        src16 <= 12'ha5a;
        src17 <= 12'ha8d;
        src18 <= 12'h250;
        src19 <= 12'ha6d;
        src20 <= 12'h688;
        src21 <= 12'h323;
        src22 <= 12'h799;
        src23 <= 12'h8d5;
        src24 <= 12'h826;
        src25 <= 12'h607;
        src26 <= 12'he42;
        src27 <= 12'hc35;
        src28 <= 12'h8bb;
        src29 <= 12'h9d7;
        src30 <= 12'h3e6;
        src31 <= 12'h636;
        exp <= 17'hf4cd;
        #1
        src0 <= 12'h33f;
        src1 <= 12'h44f;
        src2 <= 12'h8ff;
        src3 <= 12'hed8;
        src4 <= 12'h8c2;
        src5 <= 12'h81c;
        src6 <= 12'hdc8;
        src7 <= 12'hd9d;
        src8 <= 12'h396;
        src9 <= 12'hd11;
        src10 <= 12'h690;
        src11 <= 12'h61f;
        src12 <= 12'hd1a;
        src13 <= 12'hebf;
        src14 <= 12'h8d0;
        src15 <= 12'hf70;
        src16 <= 12'h6ef;
        src17 <= 12'h784;
        src18 <= 12'hb0;
        src19 <= 12'h45d;
        src20 <= 12'hee3;
        src21 <= 12'h832;
        src22 <= 12'h3df;
        src23 <= 12'hda5;
        src24 <= 12'h26c;
        src25 <= 12'had4;
        src26 <= 12'h985;
        src27 <= 12'h109;
        src28 <= 12'h85b;
        src29 <= 12'hc0a;
        src30 <= 12'hea5;
        src31 <= 12'h3e0;
        exp <= 17'h117e8;
        #1
        src0 <= 12'h282;
        src1 <= 12'hbcb;
        src2 <= 12'h33e;
        src3 <= 12'h854;
        src4 <= 12'h5e8;
        src5 <= 12'hc40;
        src6 <= 12'ha00;
        src7 <= 12'h81a;
        src8 <= 12'h154;
        src9 <= 12'h799;
        src10 <= 12'h55d;
        src11 <= 12'h70f;
        src12 <= 12'h531;
        src13 <= 12'hc50;
        src14 <= 12'hfd8;
        src15 <= 12'h74b;
        src16 <= 12'hc22;
        src17 <= 12'h289;
        src18 <= 12'hccc;
        src19 <= 12'h1ee;
        src20 <= 12'h6d4;
        src21 <= 12'hd1e;
        src22 <= 12'hd67;
        src23 <= 12'h484;
        src24 <= 12'h332;
        src25 <= 12'hedc;
        src26 <= 12'h2f2;
        src27 <= 12'h37;
        src28 <= 12'h360;
        src29 <= 12'h491;
        src30 <= 12'hdea;
        src31 <= 12'h8fc;
        exp <= 17'hf36e;
        #1
        src0 <= 12'hd72;
        src1 <= 12'hbd6;
        src2 <= 12'hc7c;
        src3 <= 12'h823;
        src4 <= 12'h1c8;
        src5 <= 12'h72e;
        src6 <= 12'h1ca;
        src7 <= 12'h2a;
        src8 <= 12'hdf1;
        src9 <= 12'h49d;
        src10 <= 12'h2ba;
        src11 <= 12'h82c;
        src12 <= 12'h881;
        src13 <= 12'h46b;
        src14 <= 12'h52d;
        src15 <= 12'h525;
        src16 <= 12'h2e9;
        src17 <= 12'h5d1;
        src18 <= 12'h404;
        src19 <= 12'h186;
        src20 <= 12'h8be;
        src21 <= 12'h224;
        src22 <= 12'h98c;
        src23 <= 12'hf87;
        src24 <= 12'h5f;
        src25 <= 12'hd4a;
        src26 <= 12'hc54;
        src27 <= 12'hd36;
        src28 <= 12'hb1b;
        src29 <= 12'h78b;
        src30 <= 12'hbf3;
        src31 <= 12'hd9d;
        exp <= 17'hf325;
        #1
        src0 <= 12'hcf7;
        src1 <= 12'h313;
        src2 <= 12'hd9;
        src3 <= 12'h258;
        src4 <= 12'h5f2;
        src5 <= 12'h208;
        src6 <= 12'h7e1;
        src7 <= 12'h38b;
        src8 <= 12'h79b;
        src9 <= 12'hed2;
        src10 <= 12'h6de;
        src11 <= 12'h7c4;
        src12 <= 12'h3a1;
        src13 <= 12'h6a3;
        src14 <= 12'h9e6;
        src15 <= 12'h600;
        src16 <= 12'h916;
        src17 <= 12'he37;
        src18 <= 12'hc7c;
        src19 <= 12'hadb;
        src20 <= 12'h56f;
        src21 <= 12'h7e6;
        src22 <= 12'h906;
        src23 <= 12'h2b3;
        src24 <= 12'h8b3;
        src25 <= 12'h43f;
        src26 <= 12'he9b;
        src27 <= 12'he8c;
        src28 <= 12'h1de;
        src29 <= 12'hfcc;
        src30 <= 12'h733;
        src31 <= 12'h529;
        exp <= 17'hf5ab;
        #1
        src0 <= 12'hbf8;
        src1 <= 12'h79c;
        src2 <= 12'h976;
        src3 <= 12'ha52;
        src4 <= 12'h855;
        src5 <= 12'h67c;
        src6 <= 12'h990;
        src7 <= 12'h141;
        src8 <= 12'hf3f;
        src9 <= 12'h76e;
        src10 <= 12'hc61;
        src11 <= 12'h6ee;
        src12 <= 12'h951;
        src13 <= 12'h2f2;
        src14 <= 12'hcd3;
        src15 <= 12'h445;
        src16 <= 12'h833;
        src17 <= 12'h5;
        src18 <= 12'hdab;
        src19 <= 12'h106;
        src20 <= 12'h533;
        src21 <= 12'h45f;
        src22 <= 12'h627;
        src23 <= 12'h585;
        src24 <= 12'hdfe;
        src25 <= 12'hf1d;
        src26 <= 12'h758;
        src27 <= 12'h827;
        src28 <= 12'hd99;
        src29 <= 12'hf77;
        src30 <= 12'h9bc;
        src31 <= 12'hb50;
        exp <= 17'h11332;
        #1
        src0 <= 12'h6f0;
        src1 <= 12'h77d;
        src2 <= 12'h1da;
        src3 <= 12'hf57;
        src4 <= 12'hef0;
        src5 <= 12'h392;
        src6 <= 12'hd0a;
        src7 <= 12'h615;
        src8 <= 12'hcfd;
        src9 <= 12'hb86;
        src10 <= 12'h7cd;
        src11 <= 12'h3b7;
        src12 <= 12'h7ff;
        src13 <= 12'he7f;
        src14 <= 12'hbd4;
        src15 <= 12'h9f0;
        src16 <= 12'h7a9;
        src17 <= 12'hcf9;
        src18 <= 12'h3ea;
        src19 <= 12'h6d6;
        src20 <= 12'hb2f;
        src21 <= 12'h90;
        src22 <= 12'h971;
        src23 <= 12'h963;
        src24 <= 12'h8c4;
        src25 <= 12'haef;
        src26 <= 12'h3c0;
        src27 <= 12'hae;
        src28 <= 12'h7e2;
        src29 <= 12'h108;
        src30 <= 12'hc62;
        src31 <= 12'h1d3;
        exp <= 17'h102bd;
        #1
        src0 <= 12'hef7;
        src1 <= 12'h241;
        src2 <= 12'hfc0;
        src3 <= 12'hbb4;
        src4 <= 12'h920;
        src5 <= 12'h20b;
        src6 <= 12'hc65;
        src7 <= 12'hb04;
        src8 <= 12'h4b7;
        src9 <= 12'hcbe;
        src10 <= 12'h629;
        src11 <= 12'h1;
        src12 <= 12'hc61;
        src13 <= 12'h1ef;
        src14 <= 12'he83;
        src15 <= 12'hda8;
        src16 <= 12'h992;
        src17 <= 12'h7bf;
        src18 <= 12'h7f;
        src19 <= 12'h45e;
        src20 <= 12'h545;
        src21 <= 12'hb61;
        src22 <= 12'h276;
        src23 <= 12'h5bc;
        src24 <= 12'h855;
        src25 <= 12'h97e;
        src26 <= 12'h8dd;
        src27 <= 12'hff2;
        src28 <= 12'h9da;
        src29 <= 12'he19;
        src30 <= 12'h341;
        src31 <= 12'hdd5;
        exp <= 17'h1140b;
        #1
        src0 <= 12'h73a;
        src1 <= 12'h522;
        src2 <= 12'h4e4;
        src3 <= 12'hf01;
        src4 <= 12'h522;
        src5 <= 12'hcd3;
        src6 <= 12'h176;
        src7 <= 12'hfab;
        src8 <= 12'ha49;
        src9 <= 12'h5d0;
        src10 <= 12'h512;
        src11 <= 12'h171;
        src12 <= 12'ha38;
        src13 <= 12'h9b0;
        src14 <= 12'h1b1;
        src15 <= 12'hc19;
        src16 <= 12'hb7f;
        src17 <= 12'he60;
        src18 <= 12'h96d;
        src19 <= 12'hbf2;
        src20 <= 12'hb00;
        src21 <= 12'h80f;
        src22 <= 12'he7c;
        src23 <= 12'ha62;
        src24 <= 12'h9d1;
        src25 <= 12'h108;
        src26 <= 12'h6be;
        src27 <= 12'he78;
        src28 <= 12'hcfa;
        src29 <= 12'h176;
        src30 <= 12'heff;
        src31 <= 12'ha6e;
        exp <= 17'h11ebc;
        #1
        src0 <= 12'hd06;
        src1 <= 12'h24e;
        src2 <= 12'h7ec;
        src3 <= 12'hdef;
        src4 <= 12'hf6f;
        src5 <= 12'hf17;
        src6 <= 12'h29f;
        src7 <= 12'h1fd;
        src8 <= 12'h788;
        src9 <= 12'hf38;
        src10 <= 12'hf47;
        src11 <= 12'h398;
        src12 <= 12'h5d5;
        src13 <= 12'he8a;
        src14 <= 12'hcef;
        src15 <= 12'h95f;
        src16 <= 12'hcbb;
        src17 <= 12'h5eb;
        src18 <= 12'hab4;
        src19 <= 12'h713;
        src20 <= 12'h65d;
        src21 <= 12'h943;
        src22 <= 12'hcb0;
        src23 <= 12'h7e1;
        src24 <= 12'h83c;
        src25 <= 12'h500;
        src26 <= 12'h9fe;
        src27 <= 12'h388;
        src28 <= 12'h980;
        src29 <= 12'h5e2;
        src30 <= 12'h1dc;
        src31 <= 12'h615;
        exp <= 17'h11750;
        #1
        src0 <= 12'h100;
        src1 <= 12'h494;
        src2 <= 12'h7fb;
        src3 <= 12'hb68;
        src4 <= 12'h8f8;
        src5 <= 12'h41a;
        src6 <= 12'h8b7;
        src7 <= 12'h11a;
        src8 <= 12'hc74;
        src9 <= 12'h5ee;
        src10 <= 12'ha35;
        src11 <= 12'h255;
        src12 <= 12'h9e5;
        src13 <= 12'h589;
        src14 <= 12'hd9f;
        src15 <= 12'h630;
        src16 <= 12'h8ca;
        src17 <= 12'h34e;
        src18 <= 12'h694;
        src19 <= 12'hf2c;
        src20 <= 12'hfd8;
        src21 <= 12'h1d4;
        src22 <= 12'hc7a;
        src23 <= 12'ha1b;
        src24 <= 12'h246;
        src25 <= 12'hebf;
        src26 <= 12'hf01;
        src27 <= 12'h25;
        src28 <= 12'h45c;
        src29 <= 12'h36d;
        src30 <= 12'hdd4;
        src31 <= 12'hda4;
        exp <= 17'hff88;
        #1
        src0 <= 12'h549;
        src1 <= 12'h43f;
        src2 <= 12'h3b1;
        src3 <= 12'h6a4;
        src4 <= 12'h4f5;
        src5 <= 12'h6df;
        src6 <= 12'h104;
        src7 <= 12'h180;
        src8 <= 12'he6;
        src9 <= 12'ha36;
        src10 <= 12'ha0e;
        src11 <= 12'h8af;
        src12 <= 12'hb10;
        src13 <= 12'h65;
        src14 <= 12'hb10;
        src15 <= 12'haa7;
        src16 <= 12'h64c;
        src17 <= 12'h81a;
        src18 <= 12'hb70;
        src19 <= 12'h335;
        src20 <= 12'hcd3;
        src21 <= 12'he76;
        src22 <= 12'h673;
        src23 <= 12'hc98;
        src24 <= 12'hff0;
        src25 <= 12'h877;
        src26 <= 12'hc33;
        src27 <= 12'ha10;
        src28 <= 12'ha67;
        src29 <= 12'hca2;
        src30 <= 12'h206;
        src31 <= 12'h51;
        exp <= 17'hf4a3;
        #1
        src0 <= 12'hb4d;
        src1 <= 12'h671;
        src2 <= 12'hc80;
        src3 <= 12'h501;
        src4 <= 12'hf3a;
        src5 <= 12'h608;
        src6 <= 12'hc8f;
        src7 <= 12'h4dd;
        src8 <= 12'hfd8;
        src9 <= 12'h83f;
        src10 <= 12'h3c5;
        src11 <= 12'h777;
        src12 <= 12'h96d;
        src13 <= 12'h592;
        src14 <= 12'ha04;
        src15 <= 12'hcfb;
        src16 <= 12'h6a4;
        src17 <= 12'hf59;
        src18 <= 12'hf47;
        src19 <= 12'hd7f;
        src20 <= 12'h8e3;
        src21 <= 12'h8da;
        src22 <= 12'hf12;
        src23 <= 12'h44;
        src24 <= 12'h761;
        src25 <= 12'h347;
        src26 <= 12'h84c;
        src27 <= 12'h622;
        src28 <= 12'h296;
        src29 <= 12'hb1c;
        src30 <= 12'h7b7;
        src31 <= 12'h1bd;
        exp <= 17'h11750;
        #1
        src0 <= 12'h72c;
        src1 <= 12'hb57;
        src2 <= 12'h4cc;
        src3 <= 12'h320;
        src4 <= 12'h161;
        src5 <= 12'hd69;
        src6 <= 12'h84b;
        src7 <= 12'h79d;
        src8 <= 12'h3c9;
        src9 <= 12'h45f;
        src10 <= 12'hf74;
        src11 <= 12'h2c0;
        src12 <= 12'h935;
        src13 <= 12'h38c;
        src14 <= 12'h3cc;
        src15 <= 12'h2c4;
        src16 <= 12'h39c;
        src17 <= 12'h992;
        src18 <= 12'h2d8;
        src19 <= 12'h5e4;
        src20 <= 12'ha0c;
        src21 <= 12'hc62;
        src22 <= 12'h3ca;
        src23 <= 12'h421;
        src24 <= 12'hc81;
        src25 <= 12'hde6;
        src26 <= 12'h57d;
        src27 <= 12'he97;
        src28 <= 12'h988;
        src29 <= 12'hb62;
        src30 <= 12'h556;
        src31 <= 12'hf7b;
        exp <= 17'hf347;
        #1
        src0 <= 12'h5be;
        src1 <= 12'hee7;
        src2 <= 12'h733;
        src3 <= 12'h646;
        src4 <= 12'h882;
        src5 <= 12'h930;
        src6 <= 12'hc6f;
        src7 <= 12'h586;
        src8 <= 12'h807;
        src9 <= 12'h830;
        src10 <= 12'hb9;
        src11 <= 12'h94d;
        src12 <= 12'hd8c;
        src13 <= 12'h331;
        src14 <= 12'h11e;
        src15 <= 12'h9da;
        src16 <= 12'hcb;
        src17 <= 12'he8e;
        src18 <= 12'h586;
        src19 <= 12'hccd;
        src20 <= 12'h91d;
        src21 <= 12'h7ee;
        src22 <= 12'hb40;
        src23 <= 12'hc73;
        src24 <= 12'hcea;
        src25 <= 12'h2c1;
        src26 <= 12'h539;
        src27 <= 12'h2f5;
        src28 <= 12'h587;
        src29 <= 12'h681;
        src30 <= 12'h267;
        src31 <= 12'h2dc;
        exp <= 17'hef45;
        #1
        src0 <= 12'hac1;
        src1 <= 12'hca6;
        src2 <= 12'hdbf;
        src3 <= 12'h247;
        src4 <= 12'ha52;
        src5 <= 12'h895;
        src6 <= 12'hfaa;
        src7 <= 12'he97;
        src8 <= 12'h898;
        src9 <= 12'h3fe;
        src10 <= 12'h4d9;
        src11 <= 12'h205;
        src12 <= 12'h5c8;
        src13 <= 12'h520;
        src14 <= 12'h82b;
        src15 <= 12'h62f;
        src16 <= 12'h62e;
        src17 <= 12'h885;
        src18 <= 12'h505;
        src19 <= 12'h2ec;
        src20 <= 12'he08;
        src21 <= 12'h7f7;
        src22 <= 12'h2a6;
        src23 <= 12'hfa9;
        src24 <= 12'h497;
        src25 <= 12'h7a5;
        src26 <= 12'hdcd;
        src27 <= 12'he13;
        src28 <= 12'hdc1;
        src29 <= 12'h7fd;
        src30 <= 12'hd56;
        src31 <= 12'hf3e;
        exp <= 17'h11eab;
        #1
        src0 <= 12'h22b;
        src1 <= 12'hc3a;
        src2 <= 12'hb10;
        src3 <= 12'h167;
        src4 <= 12'h84c;
        src5 <= 12'h4aa;
        src6 <= 12'h2c8;
        src7 <= 12'h35e;
        src8 <= 12'hd90;
        src9 <= 12'h2f7;
        src10 <= 12'h6ca;
        src11 <= 12'h733;
        src12 <= 12'h575;
        src13 <= 12'h451;
        src14 <= 12'h8ac;
        src15 <= 12'had1;
        src16 <= 12'h247;
        src17 <= 12'h7af;
        src18 <= 12'h30a;
        src19 <= 12'h2d;
        src20 <= 12'h45b;
        src21 <= 12'h8a;
        src22 <= 12'h1c8;
        src23 <= 12'h6a9;
        src24 <= 12'heaa;
        src25 <= 12'h7b7;
        src26 <= 12'hf2f;
        src27 <= 12'h3da;
        src28 <= 12'hb7e;
        src29 <= 12'hf17;
        src30 <= 12'h97b;
        src31 <= 12'h9e9;
        exp <= 17'hdba5;
        #1
        src0 <= 12'h97f;
        src1 <= 12'hda1;
        src2 <= 12'h8a0;
        src3 <= 12'h98c;
        src4 <= 12'h256;
        src5 <= 12'hbde;
        src6 <= 12'h2bd;
        src7 <= 12'h96;
        src8 <= 12'h3c7;
        src9 <= 12'h3be;
        src10 <= 12'h266;
        src11 <= 12'h831;
        src12 <= 12'hc77;
        src13 <= 12'h54e;
        src14 <= 12'h7e7;
        src15 <= 12'h381;
        src16 <= 12'h687;
        src17 <= 12'h460;
        src18 <= 12'h232;
        src19 <= 12'h96f;
        src20 <= 12'h254;
        src21 <= 12'h7f2;
        src22 <= 12'he02;
        src23 <= 12'h22;
        src24 <= 12'h915;
        src25 <= 12'h534;
        src26 <= 12'h906;
        src27 <= 12'h9fb;
        src28 <= 12'h945;
        src29 <= 12'h14c;
        src30 <= 12'ha14;
        src31 <= 12'h8e4;
        exp <= 17'hd7e1;
        #1
        src0 <= 12'h4fb;
        src1 <= 12'hed5;
        src2 <= 12'he7d;
        src3 <= 12'hccb;
        src4 <= 12'h119;
        src5 <= 12'hb51;
        src6 <= 12'hbcb;
        src7 <= 12'h61;
        src8 <= 12'h2f3;
        src9 <= 12'hb82;
        src10 <= 12'h91;
        src11 <= 12'h268;
        src12 <= 12'h6b5;
        src13 <= 12'h430;
        src14 <= 12'h54d;
        src15 <= 12'h68e;
        src16 <= 12'h94a;
        src17 <= 12'he4f;
        src18 <= 12'hd0;
        src19 <= 12'hb82;
        src20 <= 12'h243;
        src21 <= 12'h8e7;
        src22 <= 12'h139;
        src23 <= 12'hd21;
        src24 <= 12'h2e6;
        src25 <= 12'hd64;
        src26 <= 12'h6d3;
        src27 <= 12'h26;
        src28 <= 12'h7e4;
        src29 <= 12'h13b;
        src30 <= 12'h25e;
        src31 <= 12'h436;
        exp <= 17'hd441;
        #1
        src0 <= 12'h8e5;
        src1 <= 12'h30d;
        src2 <= 12'h290;
        src3 <= 12'h94;
        src4 <= 12'h1b6;
        src5 <= 12'hdc3;
        src6 <= 12'h30d;
        src7 <= 12'h539;
        src8 <= 12'hae7;
        src9 <= 12'hbdb;
        src10 <= 12'hc81;
        src11 <= 12'h14c;
        src12 <= 12'h203;
        src13 <= 12'hb4b;
        src14 <= 12'h8ac;
        src15 <= 12'h21f;
        src16 <= 12'h1c5;
        src17 <= 12'h4fd;
        src18 <= 12'h116;
        src19 <= 12'h805;
        src20 <= 12'ha21;
        src21 <= 12'h8d;
        src22 <= 12'h8cc;
        src23 <= 12'h707;
        src24 <= 12'h73;
        src25 <= 12'hac6;
        src26 <= 12'h294;
        src27 <= 12'hd9b;
        src28 <= 12'h961;
        src29 <= 12'hd94;
        src30 <= 12'h8a2;
        src31 <= 12'h795;
        exp <= 17'hd06f;
        #1
        src0 <= 12'h903;
        src1 <= 12'h2cc;
        src2 <= 12'h8fb;
        src3 <= 12'h241;
        src4 <= 12'hb20;
        src5 <= 12'hb17;
        src6 <= 12'hf15;
        src7 <= 12'h47b;
        src8 <= 12'h4f0;
        src9 <= 12'h5c6;
        src10 <= 12'h60d;
        src11 <= 12'hfd;
        src12 <= 12'h666;
        src13 <= 12'h5e7;
        src14 <= 12'h94b;
        src15 <= 12'h356;
        src16 <= 12'h723;
        src17 <= 12'h84e;
        src18 <= 12'h858;
        src19 <= 12'hc98;
        src20 <= 12'hef3;
        src21 <= 12'hadd;
        src22 <= 12'hc90;
        src23 <= 12'h580;
        src24 <= 12'h9e0;
        src25 <= 12'h5b2;
        src26 <= 12'h4fe;
        src27 <= 12'h370;
        src28 <= 12'hf94;
        src29 <= 12'hdff;
        src30 <= 12'h671;
        src31 <= 12'h827;
        exp <= 17'hffec;
        #1
        src0 <= 12'h58e;
        src1 <= 12'h73d;
        src2 <= 12'hb3a;
        src3 <= 12'h5b6;
        src4 <= 12'hf82;
        src5 <= 12'hf6d;
        src6 <= 12'h1c8;
        src7 <= 12'h67a;
        src8 <= 12'h745;
        src9 <= 12'hc6a;
        src10 <= 12'h85;
        src11 <= 12'he6c;
        src12 <= 12'h6a7;
        src13 <= 12'h924;
        src14 <= 12'ha76;
        src15 <= 12'h569;
        src16 <= 12'h240;
        src17 <= 12'h525;
        src18 <= 12'h878;
        src19 <= 12'h966;
        src20 <= 12'h637;
        src21 <= 12'h131;
        src22 <= 12'h2d7;
        src23 <= 12'hfeb;
        src24 <= 12'h4b8;
        src25 <= 12'h963;
        src26 <= 12'h934;
        src27 <= 12'h652;
        src28 <= 12'h259;
        src29 <= 12'h942;
        src30 <= 12'hff6;
        src31 <= 12'h81a;
        exp <= 17'hfbef;
        #1
        src0 <= 12'h279;
        src1 <= 12'hd8c;
        src2 <= 12'h7da;
        src3 <= 12'hab4;
        src4 <= 12'h4a3;
        src5 <= 12'h272;
        src6 <= 12'h588;
        src7 <= 12'h6d;
        src8 <= 12'hc21;
        src9 <= 12'ha1;
        src10 <= 12'hf1f;
        src11 <= 12'h76b;
        src12 <= 12'h4c7;
        src13 <= 12'h1a4;
        src14 <= 12'hd85;
        src15 <= 12'h100;
        src16 <= 12'h5d3;
        src17 <= 12'h417;
        src18 <= 12'h926;
        src19 <= 12'h125;
        src20 <= 12'h1d9;
        src21 <= 12'hacb;
        src22 <= 12'hefa;
        src23 <= 12'h50f;
        src24 <= 12'h99f;
        src25 <= 12'h65a;
        src26 <= 12'hd87;
        src27 <= 12'hc21;
        src28 <= 12'he27;
        src29 <= 12'h949;
        src30 <= 12'h871;
        src31 <= 12'h630;
        exp <= 17'hec6d;
        #1
        src0 <= 12'hf4;
        src1 <= 12'hea3;
        src2 <= 12'hc22;
        src3 <= 12'hbd5;
        src4 <= 12'h522;
        src5 <= 12'h2f9;
        src6 <= 12'h7ab;
        src7 <= 12'hbd4;
        src8 <= 12'h18d;
        src9 <= 12'h71;
        src10 <= 12'hc34;
        src11 <= 12'h1d7;
        src12 <= 12'h6d1;
        src13 <= 12'hafb;
        src14 <= 12'hb62;
        src15 <= 12'he37;
        src16 <= 12'h64d;
        src17 <= 12'h3f8;
        src18 <= 12'h1f3;
        src19 <= 12'h318;
        src20 <= 12'ha5f;
        src21 <= 12'ha0f;
        src22 <= 12'hec3;
        src23 <= 12'he94;
        src24 <= 12'h1a0;
        src25 <= 12'hf1;
        src26 <= 12'h45a;
        src27 <= 12'h3be;
        src28 <= 12'h900;
        src29 <= 12'h1d7;
        src30 <= 12'h349;
        src31 <= 12'h247;
        exp <= 17'hdabb;
        #1
        src0 <= 12'hd41;
        src1 <= 12'hcc0;
        src2 <= 12'h193;
        src3 <= 12'h167;
        src4 <= 12'h511;
        src5 <= 12'hb32;
        src6 <= 12'h416;
        src7 <= 12'haf8;
        src8 <= 12'hcd3;
        src9 <= 12'ha2a;
        src10 <= 12'h801;
        src11 <= 12'h330;
        src12 <= 12'h699;
        src13 <= 12'ha1e;
        src14 <= 12'h4c6;
        src15 <= 12'h66d;
        src16 <= 12'h28b;
        src17 <= 12'h25d;
        src18 <= 12'h86c;
        src19 <= 12'hf3;
        src20 <= 12'h9fc;
        src21 <= 12'hc5f;
        src22 <= 12'hc68;
        src23 <= 12'hf0;
        src24 <= 12'h325;
        src25 <= 12'h5b8;
        src26 <= 12'h4c2;
        src27 <= 12'hf2;
        src28 <= 12'hbd4;
        src29 <= 12'h750;
        src30 <= 12'h6d2;
        src31 <= 12'h4b3;
        exp <= 17'hd998;
        #1
        src0 <= 12'h4d9;
        src1 <= 12'hbec;
        src2 <= 12'h362;
        src3 <= 12'h9e;
        src4 <= 12'h41b;
        src5 <= 12'h239;
        src6 <= 12'h967;
        src7 <= 12'h312;
        src8 <= 12'heaf;
        src9 <= 12'h86d;
        src10 <= 12'h994;
        src11 <= 12'hc37;
        src12 <= 12'h91b;
        src13 <= 12'hf;
        src14 <= 12'h565;
        src15 <= 12'hdcb;
        src16 <= 12'hf8c;
        src17 <= 12'hc71;
        src18 <= 12'had7;
        src19 <= 12'hc5;
        src20 <= 12'ha7a;
        src21 <= 12'h225;
        src22 <= 12'h9de;
        src23 <= 12'hf2a;
        src24 <= 12'hb4b;
        src25 <= 12'h1a5;
        src26 <= 12'hcb6;
        src27 <= 12'ha25;
        src28 <= 12'h5be;
        src29 <= 12'h637;
        src30 <= 12'h520;
        src31 <= 12'haaf;
        exp <= 17'hfda2;
        #1
        src0 <= 12'h89c;
        src1 <= 12'h5a7;
        src2 <= 12'h889;
        src3 <= 12'hdd1;
        src4 <= 12'h482;
        src5 <= 12'h1a4;
        src6 <= 12'h6f1;
        src7 <= 12'ha32;
        src8 <= 12'had2;
        src9 <= 12'h8f4;
        src10 <= 12'h419;
        src11 <= 12'h554;
        src12 <= 12'h950;
        src13 <= 12'h5a8;
        src14 <= 12'hacf;
        src15 <= 12'h29;
        src16 <= 12'h129;
        src17 <= 12'h726;
        src18 <= 12'hf33;
        src19 <= 12'h607;
        src20 <= 12'hefa;
        src21 <= 12'h46e;
        src22 <= 12'h5ee;
        src23 <= 12'h4e;
        src24 <= 12'h9a6;
        src25 <= 12'h8f3;
        src26 <= 12'hac6;
        src27 <= 12'hb6d;
        src28 <= 12'h730;
        src29 <= 12'h8e5;
        src30 <= 12'hb27;
        src31 <= 12'h9c7;
        exp <= 17'hf805;
        #1
        src0 <= 12'h958;
        src1 <= 12'hac0;
        src2 <= 12'h5b1;
        src3 <= 12'h899;
        src4 <= 12'hf07;
        src5 <= 12'he74;
        src6 <= 12'hf9d;
        src7 <= 12'h6a5;
        src8 <= 12'h13;
        src9 <= 12'hae7;
        src10 <= 12'h8b0;
        src11 <= 12'h58f;
        src12 <= 12'hb21;
        src13 <= 12'h21a;
        src14 <= 12'he3c;
        src15 <= 12'ha60;
        src16 <= 12'h602;
        src17 <= 12'h670;
        src18 <= 12'hceb;
        src19 <= 12'h37;
        src20 <= 12'h5f5;
        src21 <= 12'h312;
        src22 <= 12'habe;
        src23 <= 12'hfcd;
        src24 <= 12'h36c;
        src25 <= 12'h1af;
        src26 <= 12'heae;
        src27 <= 12'h178;
        src28 <= 12'h27e;
        src29 <= 12'h6;
        src30 <= 12'h3ba;
        src31 <= 12'hdb0;
        exp <= 17'hfb84;
        #1
        $finish;
    end
endmodule

