module testbench();
    reg [12:0] src0;
    reg [12:0] src1;
    reg [12:0] src2;
    reg [12:0] src3;
    reg [12:0] src4;
    reg [12:0] src5;
    reg [12:0] src6;
    reg [12:0] src7;
    reg [12:0] src8;
    reg [12:0] src9;
    reg [12:0] src10;
    reg [12:0] src11;
    reg [12:0] src12;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73d661ae79c49f9846318aa5f5513096661eac0ba3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af8335e88e210694e3cc995e760cbe677cdc5c0b70;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'habb45068ea80b01f2d4c56cfe4f7e45f629da7234c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd759a9a3839e13f81d74dd93e617d72913180d6030;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bf7b029dd0387192fea0954700c4a789f7784be65c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1128dc8ef815747b7801151818f8bc484e6b26fb1b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he800fb910e58a8390109d644b20690db34c8dc8bde;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4752c1e5969a11bbf0e2e37ef332f72cf65cc9966;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1454e21cd7226b14b2839e0f4ad1186477f239875af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165f0872f9134de9c7bb9bf71b23ad530ce3aa8f6e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd4a5c647708cce2019fbbc7bf57fc400fe574f44d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1110e543f2c9ada2633aa55d9debc17ace195ee982a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a8af51c54c6247aa540b2bcf1c33414ede4c36903;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b90ea5d45e12657032e668bf8e917c9111a627f9a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7b4f9e71e8cd381696583ee9bb4ea985f86044ce69;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1526259ba73520a80f2a250418eff26c44d4123ca9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1855286b0e526af9b56cd0b11371f4800886af42ba5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12083c73979a4a04cb7d278320b04f428f58f587177;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'habb870f80db2eabc4dfcf67b0e3b73f3d98265b657;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166ab190126dccbaa82a3d4eaef3f1bb9ad0cb74523;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1281bb8ec4b39d9256a7f0e149a5c7ec147376bc49b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea72237e50c9caacbc1374d6cc1003604c1368b4ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1563ae7e88d13f023d8fefa376bff41e4799c96b00a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2b157c9a1c84e3c6685af00f8c0e18a02bb1e7c367;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb45b46f1376fcfc81f4fa1b0d54917f2ee2700ed5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b1248b2858b510989bcfdfdcb70287ec904db2d3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h522e6bb4a34b80e5e9f5c645e75f938ec34975e08f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117f3687f397adb9d6cb2ae132eb2456f73b12bd084;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1759077c714687b6ecf7df2c1b6214d63c8b04e62fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17ea94f1f986b4f7c08ab1d80e40be6edd30e760a58;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b48b1c96829abb062783324a0aeb4c431311e30033;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b996d02d0c51cdc4a1521c84549c2fbfd0b2eeaffa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h27db5c24e6f22c8b4a872ff77c58256bf936b9bef6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c0de26a3c9f2c752ec813d99afb582414978dab81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda33c1377f064df9e49ffa89138a0113402e67d587;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h932dd11241c77e89ee3fe1ac8b311cf0147a57dff0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11a88be1c8485dfe76996ada070747b8c10792e7a18;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dcb86a7ff85ae99fd099a88e947953201cb28720f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f5b7188b5c846f2831ba0d0b84b3bdb819ba95896;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1126525f0417435d243f9b216f29e6c77dd8e442290;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15875001223ac353330208535c2b154888428c51dc8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1409bfffc1361546e10e0c0b7a9442ec9e08615b76d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbfd039bfedf9d34c6d468b5a54e3b4bab528778111;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8cb04dc59f20764cf3ab2fa473cc09b664b7e3f7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h999928db3ca6aba915f8ef6fbeea118104897ca7df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb8d4d81f8cc08c03735ac35bf3e8ba450b8707183;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119a19e020e58f5e965db4700d3f6ca5fbd7b283d2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16760c2ac972cd50ecdeec170df380f4e83e6722270;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h149c2bf9c7c607509db87734b6a25f9ecbef2a8555a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ce0e07656e1e704d9636761dae7df07318755c233a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ee880f7380bd6cf9235087b2b3162d30d2504ae721;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2cc3193766858abe31221d1f2b4070dd0dbaf89d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he8db399c12c4e646623874191dc3e7965801b6ff67;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf008299c155fd9a512dd37fcca8bed261df5a13fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6bccb88856bd141ba47e58c519159579fcabb2ada;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a10eaab545c7a495fb2550ccd585595e574326518;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ce4a4e38429ec7577c2daaf894690f69c02325b72;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c7f693339559b0e41ffff5bbfa4f8456d6623966f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc18c740cd7e3e1fcedc9c0807e976d3a9587a5a3ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12755409af2f802b8163b15d5d9a2662de9f136bb05;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9760ff9aebe52ede245847bb089832578d36bd5ed4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfea6ad16e2feef22d8de9f47538dd1e1681841864c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7512cadc67906315b73fee8635c27a932428b43d6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f1d99ee0089b7a339f4f2a09071495d439dc41eae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e899663e8532fdfa7c47d3b76b8f01981fc2c6d11;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c277f6701dbc2dbd3110513bce3c531827ce20eece;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14bf75e8c47ed92031169ae31786c05a46629c705c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c48cc599f2bcc06a1a8125e16293408a399c05124a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17cafb1026e812e49164d4ab13103eb78960cc13959;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hddfad2d16b75e68a4e0cfb77de198d7d5786a91faa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf8112cde543bd5c1758cd9673abf1fc63873d0854;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c982bf5b6d8466367f5e2f1d56a8d276e651c07f82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1acb19c7fbdc8fed2193355d26689ea0cfbd0d0fd4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1421ce26e7b01c7db42ad518005dc8c0b68f4bceca9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h48e8a0393d522df74aacd4aed796f4117e696669d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80e3012faa1e1450f740d193c69e238b62c626e01e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h162e95c050a4d5fbc4b387602094d1c56545a2c3cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he90be427d8364c45d3cecf897868c14c67d6837e55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7892a016b35975d929113f2400123f82e327071ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50f42c07600f844274361a91fb849091535b4fb578;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h29c78d259dfc57838d208d1fa6323f5a4fd3b60eb4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ad5a1ac5bf47250afcf13da4639f89bf386202194;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11036f376927476ac47b2f969626e70bb19a2bf0d56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16fa7677cb8c634b364d4a663cd4adf9320ffbd04db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53d267c773c3b9beace6d82eaa20fb7e565b84211d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h144e4a5d05875eb91846696526054510947df1daf82;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb0841bffa521e16472f675a71e4dcfd3d87f8f6246;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80c4cea5316395a1fbb8eb0a9a693586bd199106f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h903a37d20bece19580a0445e8fa00a2db3694155;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ab54fcafc63a897f457f19bb2926b1a837129cbf41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h274b42bb003870690eddb78b254cbc32e6020b6984;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f877907c92ceeddad85675958481234effdbb4982;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12bf701e413c15ee4a5bf1c3463181e4b2e277b1737;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ee7940f6a1afa428fe088fcceb9c0e3d7f82c83b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6872bf66254d676bc6f4fa2db41365648663330cc8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha4589042df75f41fa6ee7ecff464467b0aae1bcf78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heaa284d9d2a6fb29564d091a6e999afa39d6add3ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f9254b660c812697b8f44376a8c7e809669c044b5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h124ccb9173bf21b8037f1d2831d91aeb128a5a0cc16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he51bf82891fb9f5fae5067bd36f92ac136444073e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b6e6fbe305d2713af6d23e19162733ae81840a979;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15dcc7a4d2c17e1bbe864feea54e0e139d73ba48d6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0b507f9c1490c94ae93a855197ed4b9c557e65de3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1db880977a19db7d990b7a381bf889be24d3cca56bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd1e18cbc352f6fcdca3b43f5aa64ca46bb806f9b93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a5e53aa455f2e6cee0655a5d6dd3e8b112a6436030;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8ae84694173cc43f4d2bcd478e0a8e34e2e973a634;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11df41a0e791ff15caa1f1c4f07e1173fc40be13e97;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141ec11154c184ee04296dab14e9fd6ec8bd6ae6d71;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ed5061b2feba5b46d9dd18514973e87fefcf1ff009;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13649d7a24bc2a919e10f4e34402707846e70455378;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h27132175d0b7ab43f0dd71c8c92ac153d73b1519c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7a3204e214324dbaa8df6f085b3bde15ba17ce2f9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2bcd3f7170b535e4be17d4f05bd51a1d7477500a78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h115d2f92e1213abc94d474d6857dc2c05a564f08afa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb59a4ed540954a4f98f881fb551fc030f8f56f065d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1339b19534131705fcaf478ab95284a30e3d591ab8b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1daad8cc5beec9174147abeff173593909748437c9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0fde4967284c570db28374f05db76a5f5a51dae05;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1013da0b656e661c08b47fff9ee0113ec1e346b4d7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h115c39832d86c2a92a3a6f646551a94dfb815570278;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h26fc329f0e848f7159b38359c36d7d1a0320f04274;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h98612044c694b4168133c3a30e3f41af6f17b4d615;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f0535c3eb935912d00dcb27649d3f22d34c2e8ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1326e91d3629b97d43ebd47729481a93bc7b34bbd99;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c8b123bb23224457e4c06537a024310863f618b52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4dc4548da9da0b7ddd1a39c14958eb490361eedfe0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7cd63f7d09111c1ae7748756aef560f1fdc5189bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d33537e25aad6eed68e1d56cb1db7aa5b5c02c880f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15a4232112e1f6a9bb61aaaf38fd1c45605dd825184;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h91e9ba7f31efb504b4375ca5fa50f71ec7a68eabbf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17b06936e26436b7cda1d9e4a5b421ee91349c196ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h190465f66fe7705134f63e066bc1d802f482848cc9c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d30e234e6732898891525035ca565dcc9eee09fac3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h121fd1b305dc8e6d60c6c3ca8b91986a6af406cee44;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1844d95e46703d77b0e39df06a9355a8f65a14beb38;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f55148ec25a6a8713de05489e42af69274219ed197;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10efc2d30f786e8aa5c7ac35126fe871a3109bbd3e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10678a55659691701ea359244385339ed7c610f6bb5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf66ffeb9f752a228062bd0493e746f6a2c3f9c3da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bdbd9e96924b30e12d8dd9a872d6937f0094f71417;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c2d5ab35d29764950e47124bac222534b2b8f41169;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172fe6f3c8dde6c8cdc568d89e41f2b212810ff9b6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b983107603b9de773aee5d67f288cd624ea0a1990d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9fd42f6329960bfc2863671e0e5002023163959e43;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e7d2104a8a9d30fca2d12aa4b7e72c7f1479e336e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6411079a1e396c2907f1a9046281907af4cf47d603;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd43727bd24b179cf5030b7d6cbca8d03dad6277c4c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a27778735ed449d2bdc28e8ddca1767967cb2a1604;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc3eadc4f63958155171a6e1668e7d4af93b72f079;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6bdd80cd7097b9673e0c18b1a0e9eec3e81d12ab5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b90bb8ed093b3836e795788e1666c1f5b140c98622;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12032f0febc95fb9e87ed3a67f07c728184dbdab09a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he9a1bcf78e55e063375bb808772df72c527177fc88;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha1d7469b1ce41493cb1c02ca9f9a2a9f06fe0679ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c0f95e54acd26d0021708b8cfc7323a234714caf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2aa7afc4a707a769af742248aa0c2385b7f723d4e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha51ae749d3d34fa3d7da0924189a564f4012479ce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h325982102acad59e46b77d91be0d649c26f8afe15d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfc4c74ee2fc3477abee11c44e6346dbcdc9ee9197;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc2635f67929ee5d589ee27f2572777f3ca78785cb5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9beb19849a5a342bedfc4f2f3339df5783721660b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b337c07001bbc7248ca2aa3453ee556d1bbc5f0c8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ea445572cc32290f559543d7712ce47a09e220c06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h173e3d7605e0e8d0eaaa4423f1a5f3939ca24ba40d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hff8e469c395239113c569688f3d623240320d8d124;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb77ea6f02b6d938a61033231b06476dea267b05892;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1062b8201b19bd5b52979efa02fc25fcad2df87fa7b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ef0ecfbc4c0dac7b90746df6f983eb09874f6d00fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1773295e92dbc41062844a508a45cede6a61e001a60;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1701d74e488e89843963e10a3975c93291f6d6e2679;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h699d60015f5f6a72367d69b3e5cfd3063db282888c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd1b3200e315f4d1152fee33fd49034de0514c6c7c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19eb10a8964b5a72be135fbf35ec7e298a36bf1491;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f116f473045903ad55bf963d740bebe668a21f96d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b45810e8295071ea83a9fb485af77cfbdc001f9751;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2aee67e14f53459bb18f7be12c042e188a5ddb30be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h167d5a388d10fc3ec50182773b9d4a86f75966307fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4f1dbb6552b8af6074313fe3165e098e9458aefe30;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee1da3ed79dac1fc40ab08747d0329e0c004b9772;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82235249c16e2c2cdc6548ce02e1825a1417938933;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0c1db605ee19dbc56a5326041671216aa4bf72f36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a2c336b8d1382b387cebec555418d7875c1990ea6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a7964f4c960c2029e2553630eace9145ee5cfebd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h312688bc142ced71dc344ce529b448f8f4fee6698d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5203a8382400973660534458318673794c109bdc85;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7f955443b5f0391f5e72f82ea58f7f752415e7cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15c80bc6b3f791a270a1aacfd3b771c0a9daf99be7a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb0ebfb60dc4e9bf4b4ba68edd3b9cb00e74d56a54;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7705516519fb91da3b2e9340483debef80cccc0e62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h655063bca2449afc561fd7d3dca09c53fe578e1e36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f57f142032e07c8e54f5f1c73f5752c4498ac5849d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h428843e4e45a555d7ccb3765e82e98f3ad44f0fee6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h500cece7e82c37f5825d22f74d85b5b5c821f4dfcc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b860cfdef18efb48a0bb9c6b49b4af6c78bf7d6f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3159b9ca05c9d84dd01381e277857c7de773f1df37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3d4380f0d7c2e4ff18b4727757a64664bac54af2d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c4319e5dc5a450db80cc7d58cb0b3230840453bda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3b71b02b3d90faef32f5002b61797bb96e5dc8737;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126b9ed6077062eea285d663140e5c2e2fa01944039;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d75f6b192d1a715ced2e5ab45d4f314acfc44c68ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb76ceccfab01dc9ca2f9f35d1b3e1371b205d7deee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h343b610a0cf64241594403e9ade14ed29699da72d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0f778bea6fd9785c8d59c6b7ed2ed411c9528b22b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d2352f4410af4af3176fbffe3330955cbb499332;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1718ea7e1ac50385e4d692bfddd9ab22cc04cb692a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h69b7d5a3571c3d04d2f1a577d8caaae66063359601;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7309d2b4724e657b791f043ba2418f433e6114a9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h427d2b2cf378dab3bb4f766836ce83d21f233bb16b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11334e4053619ee183db3f341ad13d57d046c774518;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cfdff0fdfd387ea59b316a7f76623be93c28b28f31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h70e4f50e4a53669fbebb26ab59943d7d44bb7e11e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7591fde2bd9fcd6a3ee7eccc7c5c34d91af2dc0803;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5e198ecd2a7b10bb1e8b2f998967cf6c8a805f84d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5ecce518e499fccce6227a05f9a618d153bbcab633;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3e5332e649b732d2f7bfe56312238ba0e3f82479d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h27322eb22794f7251d5522f496af79b9edb6428fed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1745d8dd8b0417e5d32f93d06854d60827a9b5eb28e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae1768872d63b1195c3b7197d524d194b2f9daa08b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39f85f779c430e8eb8988f4c2c2d925ac1bcfce850;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5257cbd5bd3851fb23eb2816db147d8f7b85d1786c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e9625d1e1543135eaaffc51060e4d557b5971cb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51e4e631506737c489378dd205467526dfb375485d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7ee9d137209f0c92529519fb98668f9a5da725088;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h58d31e497d3642cf2cf1defe7e559b7d9710d5fac1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h71ba18be6cfd3fee25ce925b1f31134fca03f23fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c439a1075dfc4f85647b8c41d7052267ad298a703;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7ec3a455ac5dafcff947abbae4342d57d49279ce90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18448efd4cfbd2a0d25c2f860fdd8db28ba0b9a3642;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc177e99b747362224e8b854e664180f5d9e52fd430;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12aa1a58ad8038a183a56f33c9258a8cd635911fd9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb60e0142e53a5489e2c4c14d6da6223eac963b1907;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hedad38795b58385c22a00e57eaced81de79b573193;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbec073fab9f360900744bc1417d579cce9f566682e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6d35d8dbb2fc18ade541c396efa0d81a2a0b9c5531;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e92978cf228af3e20e9198560fb0230ad264578d3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8478910a03d8aad06cce10e9722fea6732dcbb0c89;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heafdf2edcb4918bd25c8d5cc74f4326651e9361b2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h164b1f03e32d3a4ddca79168e00d1039139a2c3fe4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16563108006d32e528cd7e5b1cb8d7724b9cb062b2c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea9c41e13c3231fa23dbe8001787dca3814d4697ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ca3fa6751f98062c350e6cf0fba1a8d0a8d23526c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cc831acc01311abff6b8bf75a784367c88192a8b80;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e247cb35b584821acd6ec20fd8da79c3ff00eae0b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e77d27519414a5bf4236dfdb08e4ae0ea39cc66fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h131f78d2b0fa483a2596d8d53666d407d7261c0ac2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1356a960313c962faf66491173917e975361a02e490;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14861a85793656a0df2a3bd408acf2a816f3d9f43e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75cd4d50e6b3bb0aee66b24fad629e1c52416360a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fcebab829afaf54cab6760f74e419542539617677d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1ae7c55bc69df16127299b60704d1633b6abc4247;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1631ca9aea012c864b24834ec983f0f01bba58a7afc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117c57e47aad27bf623a68272f1611bea671e57364;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1144dc5f834f5783167e043c4ee93d6c446f37a8572;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h390adc3d0d9597e2d93a46b41310954c6f897fb07d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1c93f7cce2e208da8ce6d610a0e10e8cf85cf9965;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h582fc6d0056479fe2ddd659fcc3a0744af3b0e56d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140a745ea73b82d8e3ec937fb1bbe8da389ba3f27c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d67af3b5afd3bb8bbc223fc0ed9c471f48263dcde;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5864e159b3b7f34b35bbb046995d58be195ce4cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c72340e48a64bf4c0248e1caac8ed3b5054ed78ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h96891cb95b9475d2bb345fc15c1ef2fd9ee6048e2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11093b88f67fd8cc59deb100045892e0eb3aa19f595;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd97fc36554c8b233339c7a7469babdb0fe19cdc37b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6d7363f8236c92d507d18c0a12acbfbdb5563e83c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h987ee8a9f69749d2895e26d006ede6fd3790cbb055;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h380f6f85f36857a093c6377e7ac4c1e06ec6065b0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d6d0d00caf5bf973e077a8658b6604db24a032985;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb403708f0a10e1a15634d31eacce97dde36bd0b3c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hecf49c6e8b0baf6b7c88b0c7611fe2db26d788bbe6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb82ba99e2b6301df006d1e5388dbc388cdc0b642d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f28dd6470b6f8ce3997839faaf23df6eed9bee1e09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h76fdc5d032b836873f278bd197c42f59fa45f5d72e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ccd984e8b9e773e1f682316e65b9c43dae25ee8fd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he90143e11df5821a6770d6271401664712cd59f2ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ac67f2426d7630cebaaa02219aa43e0cfb3d35846;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c71c15ea133cc68b0924ccfc6148e7034dc2d6380c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81bf1fba80a4942e360f5adf9a54064ea7b39a2e0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd3c8010bc8404718469532eafcc15dfc0897d8991;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6907f91d4faf72bcd2a97c22632844513ffe4dcb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc556c3165510c7be008c5222769f0823ac9f9b729c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dbbac641a84fd2ad7ea76e318a4b8ac2ad798f6e79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ffa633ffabfa39e84ca394962ebd179f78bfa7d1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a5e8ebeb10e72f2a25c6e7c12fd0ac19b9c3d2cf48;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1248c3f8b4c7f05877a10801451f3c8b47862a01841;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ff9f43ebce5620f5302774e5e698432dcadbb9b523;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1baed884bc78f3276ea19dc56e7d2fe20e9e6b0f864;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf925d27b9e7ae7ee8c61b4a1668aa8506ec400fca5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha6325ae02457e56db9eb9c027bf53d706fb92a8e52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef23d68a37e463c3b6511e1b39d2c3476a291e3bdf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8aab0a69e1c0b9b68f78d76e0fb54c847a67aa490;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15eca4521b1c2ac3d4c92b31b47d47929a000da4fad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1575b8745212c97bda19d7d90826232d3c9be917167;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12bb66236796088aa2ad88d287576b60e386483e6e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aac7a77e1338a1c5052763dad8160051c7157c629;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c979f6570d155f049160ac44ae1665938639aa4fb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87df801b141864a9db27710b51cd4bbef4a67c8985;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fae5c744300ef5615d086d8adfbcee578b2ac7c952;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4827a90d9d22562ddcb94d94f322d2c58f0c906b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9aa509810f9ed299276ae41e0c3ce27bd9d0147248;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e18d69bfac5b96d0bf8d020856b801e62410514407;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10dca86f6b89eeb5551316de4c3c1fc114fd84b28eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb564f84591866a8dcb200e3ff9a58d765dc595e245;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63e141bd28fa9d508fb245cea5035628ab5f5def81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44dfea4e7194f880d288d04d965abb7b107b907ab0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9257b0260380437f893ff2e154371473506c0f3dd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1135fc4916fc11bc88c3495c4e7773631ece2a94364;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cfa1dad11388651864b08c16edbc5e99e0f1b735f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb3f21e6b2c2e9c2733b1d8128f670a8bfb9d101c3f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1228706ca58e478e27add647e26a5b0065dda4604ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b58aa2b5dcb1bbb6dcbe105c3d3addab576d58c90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1c900b954e54cd00bac679e83a924685b3742425d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135005ea4dca28cb6d642345aec51a5358940035321;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12101ff043a712c8265bb3b11d548da4d1be5569dcc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d5c9651da9bbe5b788a438ba78bec9d0464a80fc1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d847e940087730fe1e18c0c5477209991d1e660aa8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1253ae0cd4217483aed3cdf14472b7ee507cc90eee3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7313414489b24a30d133f9bdf35ab912011321a470;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdda48b0a24e2e53598757ffb62050889ee2803c2e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfaec06c133729b14f597155786050abef468ee05e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he68fde2035fff24382688ae3cc254eac40eb2687ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6168e9216a84b567fbbc81afd34ae1d94071c0f343;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf26da9052ba3678b5b6cc91274ca0a59094401999;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hefa2a98256ee8d0cfdb7532731bf43c3383a71c05e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13dae36ff8f7fc4e42ccee7dd3d187110cf0d999e86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1036d09cec9fff27734e3b742439f93e18dcfe04935;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda9722a46c7ac419c9a99c75a70afb6be51f457895;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19880b706e99cdecd87669506c88e6dc40499079510;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8ead21cc6e1238ee93b837bc010a19b566842f3aa1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb38d03b12db78008fac6026266c361da0604299993;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h319abf1fb21bd692adb46731dd6d090bee4e07b47d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3787b023c84f0953cf6d9024031c5340e980e42013;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c93ff5f0ce96660ed4ee01f3c53b1ebd901af05894;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h802d15375015c8a002873dd54d6e083d21d7a4ae32;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb323682b437478a66b54cea30a862a54014f83d58c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafd58510928615d36d6008442e63150ffda7530cee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16069040a7cb2cc228e07694ee390d324ef4c52ab37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d3ea1772d907a51bcdf7b93adf9e475747511992b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5be68a8d3224e93c0d61099cd69bda9df2d09e02b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he07da7741ad264499f579f2adb99e7f004666ddfc1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbbe31d49d925db1a199ab778a3b844bf7300caadab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f2cf2aeac0231e03e919f9f5999805d11a59e0f4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19dcc8a19427a46aeafa15230ec00a3d9d08b7c305;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d225c5b82d9798c18d1e2b4b1766c264b66216e49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d1ebf0eef4228d7c8a3ee960a91714873ef493430;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d10147891248831dbf18c6ac49e6f3ed237c0b995;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10dd97c85bafca6506430487b2ae60fd5ce2a97a7e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb38f373c7cab42308550c164f4e0c12a268f4067fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h77f04ad052f1f14fa26f439ba5f882e14872babbc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc5488eead19cf591cb200f8e17df276ee08270be75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12d5f0ecbd3e01db8ad1264faebaf17b562fb4aa8be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3f5d7cbfd182aaade01fd79e20358c9d506a1eed8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8139e74a1600f40606860de3e20b614d13940dc3e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb01eeb7b5f33a6c13cb55a75f595731c20c84d48cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13170c55f2abbb34c61e545bd02c1b658b898fc0d9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c0f68b70f5d73bda6d3f239b0357d1aab0e23f952;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7342a34f2b69be17365ad8ea83aa466226891abce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f0a7a57e73cb6969403ee587e1b128fb9adb1b29ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1462ca87356b63fbcc76a8f801fa791305a82c7be78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12464db9f672c1c2eb5ef880cdeceed9739fcf97106;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h124807381c8a72a908faf2848b78933cdb91002abea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h480f4355580d2bf876be7103ebf674c10bfe327544;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13643e4b247a328461a92641d73424f65208f9207bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15762240404a11bc65d65bc5fe6c1432031e0f647f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16acf5bc6e3f0bff6d4c9ef62f8700a19bfaafcec6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h35320587161845327f351643c0c66e53db98aba3b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haf0b87dd757eeabd11ef9b8acf3a43320595378b00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h454112662b666b9b4e8177e0951f7834d11779d90b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118515823bbaa3bc4e4dd30f05a3e35593b21974993;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6a50c6e174b9d21cd012de871970a9334a9c8e147;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ad78e38f01c198a57ebd1e9d28cb24b6f4e3f151c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19d65d7c257dc08fb1f45673b4c2a918fbb8587ac06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12423033ea04bcc4e8060e89b9cb4b1800af72aa708;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa670c9cbac328e081ed690e83a246984d818bed57;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97b73c5041036b4f5fc7c662423c617ccaaa5a2f47;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e88c0e5d141a2dff855d1941eaff6b581a07c58e2d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1afe66a04db312ff2cea3fdae2e3dbbcc3009858988;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd9d86850987c98393b68ddd09488c2f17b51fd9c09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87c4a4da325aa1036c6bfa8b02b41f71a9499d2159;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d05c520e7f052b82723b6dae6fd7f37139958c38c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8cc8ecff8fd7f0fd34e4a0b03327cf8fae8d49b03e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5f2b8608dd687e0b1fdeed5c3eacfa2d764e2d473;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c48fdb205a5bf17ac3bfea7924730d342d11a595f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a09d2e6a1b3020aa49216a1132df98529477303459;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140b3f3098f6d2f0ff732660a457580c6e47505b808;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h71295ae93d5feb0e3a72673f9b7c39556ec7100361;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h159d8356bc6c249ccec369dd7e48354aa1ae99eec38;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfae5fed06121159ab22af19a7d4f8d7826515986b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1294ae5c3b3c69f10217d682d68007a86b257684828;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f00b3beac043b3c901aa3bf48ac44b4e9bec0f4457;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10a6a20fa4c08cc0ec90375bead7ea88fb434d62fe8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ab3fcce0ac71486bf77ef2134a2cdcde0eaf26f73d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h96ea79b8bd97509acfbff135e34f6f335029a6a762;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c6022a56e9b3114a00fb96a415bc795e3eb05b7669;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6affa40c4107a8f7be631cd54ed87bd2badb412c28;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbfbd6357f0838332bc5d8d0c97db4fb4a0af2c74b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c39f2f55a1934acc68faff86dcec5a1f125d17137d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110652977beafbcc34bc1949b27ce877fc2cfd557d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1164e59ada1df7ae641c988a0a94ce5e721553c0e2c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h61bc7604bed8d2aeafba4f9f9abc7af43396d9077f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h863f368bea2f32a52908438381ecc88631906d2d10;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106f047ce3ca885d8e016d080dc643c0d1f84da0b40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h408737807bac873dd10e72a83e5f61674d7f9e48b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h929aed23d215f2adaad37b0a486e789fe9145f722f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10419a369a2dec70c7c71910d7a5b4fb3873efa3a15;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2fffb7e12bc0f9557af0f069ad190586d8fd23f87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c18e459e0279ca13f0c84dfb22ea1349e9ebe74f4e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14ad8c1f3988237d5a06a875938156ce998ede547a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he7212d7d7d1552fc963fd5e740d1a16396ba482b8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ccdb333a8c13ebb4e15e9dd189ff8423ae6701c1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12070b732d2dc0669eb4e1d256761a318e833eca958;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1375917dad3f6f433703d1ee1db2f0739cd5ab3427e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193267a64536a561b2e21a0f7eb28d9404199328f03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ba03ba440ecab76e8a28e592a9f5e9678129be412;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h527b46191f61a2562e9c3ee7ccf5f2ed69acfb67a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h44910dfd95c9d999053da02d66de40a78f08e423f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a554717dd09440a65ae0af07ce8b6adf7f63c04c27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c39dc7a3286a54b95de513361ef164cc2b06f27206;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8eef59bdedff6a1d87d12776e6118ec6c0a31baf96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf795171523ec058acca1ad658a81c28e6cc3b79a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd603673b0123f6ca158fc0f1079f5f04206ea9cce2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4df2433640f847f6882dd64e0983d6327d7feb3009;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22ea99fc498f7507bd4074f230df7d316365075d0b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d79b3a9bc577081164c867a2da2b0ab21ca19480f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2fe3f807dcaeecfade89ceda6828e478e372f055d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a5f11c7749cce045305727f75392415f56298402b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd214f5e1aecb9c31be1b7395c29743d4879afe8ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd792e64b0189355a1b916dccc24517841fa9a0e92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14288ded0e531c30c840467c07d875310f8603cc2d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf37a45d3d6a6aea245a62d342fccae60c82d0179c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h146a6e0386a778d28bfa8eee2df0026e2705bbb4245;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9687030755234231443f841cbf6567fb7cde8f55ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h168acb514e2024b2087bb310deb015d4a7aa5078f35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdea9d910a284fbb42a07aa8c89797324f82c887c87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63308fdf6eb63ff5bf52ff47be04ce883139962f9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a6ccb3797e6ed89c6f9287474cf086312b7ea57bcd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10315ad359f5e0aec6f170d6b0b13f56a011468f8e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17de10fe64c94661cd1c7c13dface0a620a795c83ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h94c319ba4945823406c922caed972243891cbda8dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d044a6c62c186853e42f07c35fca5716202efcc9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12651e7672f5a438d1448054b486c41dc5044d26377;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a4ac73ab4ca379d321f42d2289f4657db9d9aafeaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b5b389e48f474dac08dfc2ccb78a505158ee536377;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c01875533912502ad0372d80f27190e6b5c2ded000;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a20728a2ff4e54e750549ba824483d3c48a7f797c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d49b4caa907acf9e8facce5eb59d6a31797e6824c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h98aa45d9dbba7eac97f2ab6b14d787d57295d31c03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd818f857670a338d4f16d98138dc1ffc76de79f329;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1403c72cbe0911027f6fc184e3d48e716b61aab7d7a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h59f68adf5e48a24af3cd2d832519bcb594d84f6dd4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153f66e22088b1af215fd17d2cc261d711312a1fb37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c94c0f351b6e2580fea366fc2d0745107414075238;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1667d7df6c13d06f5ae1209996b750e28562c5b22a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c4ffbb2424e6062dd740816168fcafbd4f97236b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19035d16fd407058cbed4583bf8b8c72ee626f2f774;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1408c12db71e9babe5dc427e2d53a108aa57d5a71de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f0378a998063742161528e893272544052d67d3ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f58542008bd6079a4aac1d0f88ded726baabe41487;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17282d8cc05ea2d39c6a8a0924105f54ad1735860f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h59ff016540c56af45c7ef544a089c785d98a623b17;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc716afcc121d7eb7c71ceb4f3181f16532ac4d63f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f59b13bf1cf102379b8fcccb0b4e9c114bbedfac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd312aea14d10e42d287b5da7f2f64ef8e60bef482;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h185de27ab5804a26cc65ec540932f23188f89948910;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0ad02ef8dffb4d139e0af60ec1ab729be45aad6f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6edd36f9493e176175bcab437d7d25dfe379cf718;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed850d01cdaa3b634fecc0baf75bdf6e25f9ec6798;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1541aabf075b8a0beba9754c029baac3756d077b1cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ab686f6d2ed8a39e48540ee9e3e585c94f9da474c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1faddcdf2ce173c0ddbf061472787d853c93c2f44f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h111540bb256f612a94122db40d41a6731ec3a1dde27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3dc6147be3e82897de71781128dcc39ea1ae79c06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1595f47e42137ccdd3d993f01de405b517d6416cffb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h76ef7eaf0ce22118a788e7a82cbfd928514d864b4e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f472ff2f29f6f71f13b49663f8773bf7dfcbd2525;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb53cfc331c1419fea24903aa35adfaec1816c22db5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10055c43b1cfe43f7887424d615234be558c3d6ac4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0dae062c5f5b562775bf03187e4d9168fe9520d30;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h104aa65ad0fe0855cbc84df2cff97fd8491d86d8970;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d3bca7d60f54187f5d48dd4c878926583c511565;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c63089be2b39a0c150a7e22371fb4fd6538d6e5c5b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8561d62f9a4bbf1d4e2f157e83ae238d77a0744021;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a0d8d54784d712a262ad7cdba6d4ca403856cab51;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hada75fbc34d3c8a90f238ab998fd59a5f70c14a48f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d2e3af47619ccc5232541ca6e576d5c2af3948421;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h381893eb10bbdc147d332ae335a221dd495930f06d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c264753a8ce9df7b6dedca8bb7721c017361a380d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d7dc1f60aec4643d770bc1fb0b6db644e068f1fd9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b42af7653611f7a45f43b4002ed43cbe536cd04f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cfccabc0003d05b1202d94341590bd1a7d75fe9a6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c1ffeca23dfef8a47de9acea524e2667ed942d6bba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1690b055c875ccfba82960c7c27d3ef620a9f5e4699;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h72274a82ae6725050631d1817b1c222ad9cfadff92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h70dbe8a307da3707ff019647f8201a7f0d59bb0e24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h40b6b48c22d35b931ded9ff5c96eada50007ae24b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1148c7a9e2b59fe681e06e535dececc0aca4bda99a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he696a00c874c4fd989c3ee8ae440b076d4385cf253;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6f282476f9727fe55c9a472c8ab62daf8877bd5fe9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1390c85d7e14d5c71f16d96425d2750847367908a3c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf184760f3a7dce15173fdc027b0a79d6fdd69a5cfd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ec2acd6b1e64af8a329a46dd08b6e0325f94e8d0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a06ff25aa95771eb3c6da03d2dc66d872415de0ff6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd66784a02e16e6635c7f99211b7edb8aae78db07f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a0e7b47cdca393aebcf1ab2ac970063db3749e44c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbac7d49ba0fee9216ecf55b0e9d38a039ce8caf183;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ee8b0ce856b9be7384f7aebd907920d938682c44a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17890d37c31c760d3f95ee86855d1e0ae67111c1a63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he73487507cf1a968ceed770a791528931636cd21d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a00d6d2b047eacb8e5c9e2b87efa8cac2debc8c68a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3720dd569bb0ea6f0598e467668383688e87c55618;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3d6855064ea3590faa1aef49ac612136555776e0c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1267e124cd3f5a05e798a91a1b1b1ba3f3ba1a5bafc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3ab20da56be5f64dfa435c5b2a6c24d24379510604;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e386bc6049b89f2e33a7c527f76e980c2085bcdd62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cd5c605ef20287038aad3f7cbdf9676089d57ece43;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ac618e6396a02beef769421752304af596acbc79e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1020b0135962f8568af3cb8d659d0d375ec1b2abf9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e158fdc6f0a1fc2de4b17e71423c9616b7e19b506;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf33cd39cd4839d3e24f70284cd20a0206d4de94e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4dc6211215c651ad89b5dc238b77938149e0521f27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb9162df2efafd9827125690fe11b635c461ec7b0d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198a56c1ce4621a674de523fce4f24882e5bfa19cb0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e3922d0c48deb997068a9c15f95d451190a6ccbda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he7146ca52a2b75548cc9952ccc06408dd5e3d716a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cae724cfa244a9a1e514aff2e8ada74906f129c065;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1c31ae53311a9b4162a7e294ad85823e408cfba42;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b3f0356989dceb90c7cd92e9d8ac59315de7a9c118;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3033934efb24c95faa8d841d31fb695fa1f2daf0ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf7d58976d6f033af46bea23abd588ef0de0c41ea5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ea4bb5e3b4a54793ad595400d04d31f1e2245d056d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hede4cb4ba8ff36fe8bc0310975af3575078b3d73d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75354bf1807b9bc9ec5e5a753ceedef2e5adee16b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9af529178797f0b28e6d0986b2c020fb8cef33387a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h35d5c0c1e224daeb1a8df2c0cb451dac022f91910b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8c216e1e67c9c7ca7d820d8dbc2613be418a5d8c63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hab684e0a96ef59de670c405f78175e09cde19878bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he447b3f9d1c8932ee0fd4fb3f6561f6692d5501a29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd41d75da32678009ed0dd9dfad77422a5cd4e6d4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10766df530564c426955b8c5d9d7877d0210080575b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a650d858f5da4cad636af058ccb97760ce07bd25db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b60d756f3d0bbcaade2e53ba955d0b57e6dd26c8f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3f6119f05ca8da8a3900d9b3c4c8f0268ea28b997d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h69c6b4930c5d881e3280646d7e99f4cec36cfda79f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce3c13784e842a7f5f22f3edef8c0ea37dfc94e323;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1da3661468ad66143fe8c3173175b63674749db2ee2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h181da2c0b178627aab50ddfa73c10305e49b64495cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0bafcd11f5126c3c4584c0a4ece1464d4faa11fd2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e899bbde5440465d279b06688af24eb7164f827d88;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51b6179795353eac5d8a062928c900f87e4ed18d6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe655352e1a0da16620052f7e538136a03cbffd2dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc97ee48cafdb8fc5de5309b7164ee01892f85786f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15fc9beec167ed8a392bfff05ff27648c1c6673009c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d7b21f0ce73ee3c0ac789a43569050c8d17e5a25e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12608659c2774109a1c89a3f99caae3ea2478cb2d0b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he763ffffb6ee2c9894871bb6e96f15ef2d6a1beb7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h99a5f384a271211d6ea7f2e07d178573ac7b658bae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ecedd769a97aa3753cd5455a1c2831de97a6f6d21;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b04373fdf823d39b50e975f5e55e7ed057def25b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3dde6897ab5cf6e336d130454a50e8c7f28a8a482;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1838e32ef5b6a69ade25b0ed4dae5d662ed19112afb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h91ad35034a6b3d58230896868e52ad2d341c7d1341;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8cdfa46613850d75adbb4760141a48cdde3907fb9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h235971cce0ecbbc05e9de8fc25e55a5a86b1ac131f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h92ccf33e14160692c7f79d093a33bd252301b679aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f984bcc30b3244505510fa18942efe383d1809bb9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda08cba81184d85091c18058ca3dbd66ba98af98ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbfef3b9e46fcc22fd210e0545593ebe74994f9ef49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h668d0130728f6100e643d63722bfce491d74c3ab40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f0bd97556367f37130869c61f374c2a17d1cdcb9fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h155e9add46fc6dfa8d6c4adb038f12b17f84b217547;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4580d7c1b486f8a38502109e90bbe35c19a4b6f887;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b891e14b30bc6abfb56223261f543762a95ca32855;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1210b8e8fc93630c90d502df7f26524ce8cba7e973c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117694934dedf8d896df0621f2e0f8fecb42039c563;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h999625a6af5dd41819498e8646ccb5a078304c27d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h816148cc3de07787de4a54b3b24bfa99b7c01f4cc4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ec050430b7928b5a61c1c235ce9bd030a94d10aad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a6f11a231b7a85721432bb4b0dd5b6a206401a131;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e4e3d5cc1e50fb3d2d77d28b3234b3f275c2aa3b80;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf84f6bbc3707fcf1ba2bd09431e460b6f25162471b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h185fdf2473f3cfa16adb7a4f4e2ba75bfafd53d5580;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14dc3bdee07574a0c399a501145dc854b3ff577d6ca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h207d0f54781acb8e3c6d46ca64990c707518dbcc8b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd8e60f47f269e2914269f36e40a5b32c523baaa147;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfbd71bb71c97f2107d17ee5d91777a67bce4d311c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h634a515bcc1eb6b711cd0a799e0f618aa4c3124dff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d04ab897e9376e1eb23b9ecd2e79eae6cc7600476;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h133190a3802d419c6eec4dd9fc28733bdcf9cacb717;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e087e70cc53a360d2d94409596788d32747d3aa144;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc34c4805f9fd35593d21d361eb6879d4bf5b584293;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1976831addad1ed09c8070fb7d222979e3c9f422f02;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h125043e594b199ffd265d81aadd94539c2bd5565904;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f32910d815ff2c0458d8d6f947d2e4ad734414d0eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5cffa5611a5965693a8b54bd64066693da8e1f1619;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165f6656c3e35db759ca3c7b60d56777f2ea582342b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18573f2e4f6047f4eae0910f8276f813d342f50252e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18770abbb1ae43c1761ee0b46b2258089f32dd00d41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d6a7d2f5c9912ab3b1d2a3d68deba1cb364d81ee9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdfeed440b38797adbfe8841e60c2f92c553933801e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ec6d592df0ef2e197524e3d6b6c2e43709314305c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118928001ff119ca1410f6947e6ca4fe7a70b966299;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd19612e7e27455b4150076d5391e822bfeb11491f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3fe93e49cec8bb698bed16db64fdb25cb57a1f1f3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138e4a3339cb0b33ea66e350ddb6dcb7f5349d808bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hddda4c866abcc8e09bd2c81355c2d52889fd43bce4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6dfc15820f9b0c7a69c56289b5da2955306174bb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h424c16530330be33c9e923a571fc4b2ef27facee50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0851bb2b3176b9f0184bbdde336d720f216af79da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h331709e252396e287f734392e7727fc8d79f766f74;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14a661f667584b110b63cf02cb6b4bae803ef493014;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h32aaa69dd5251f5aa41eb05d493f3a925902cdc759;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h88355dc0193a652a9d838005f753e22f041e39efb9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17f1127473c3350986f3f6a00ed9ee23d9d631021a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ef06198450c0647ff118ee42b450795004514ef1f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4fe7a07ffa6970e0b397a6b07d68912504805c8c56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc278ef2a7a2c81b4fd6f42c38b147715ef956d4a43;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1297da4ad7be913db40607a3c81792a8e99c95120fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h609349f90e689232d0b6a2b57dbd91861c2de45f65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18667b420107e94f0fe2437a8eee527dcb145452bfd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h106e8c6079bb512c7ba36d700ef6ad4d3445ef40f00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h193f27b00e409fcdedbfa4bb95fd81084ee94deef77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f95aa5ece08d22e52114a120db7d6266f55e2c0ce3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d97e5342d8eb602e1871232ffa75ad2008319f73f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hde7fcf988f0fbb4f755ef28fcf65eb67f49ec15cd2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97afeb70a54f7a3611a4b67b16d393349e4f9d767e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h792f3586e3d309b05dcbfbea1dcd20342d015f5674;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd9f921cafa95dd08ca45478f7ef20349fcbcf059be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c0aa4e88d5a6b3382c9a09811e1335b1a395c5505;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c4cce745b608feee42f22b64df602fb9354335f193;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19dc81965df36f9195883f64cf02b30239e472b7b66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2ad393585b7ffb8bff3617cd0ba8f1bfea1360703b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12869b06317222d07c154fd97a681b969aef38efe06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e5b667bd59b3d9e81b07d81e3c0160c86d2fe082b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6e2db0f3d2fe058ae8c5458f4cf4357b27a373a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134f66373b7f144ebc355d782b3ddb9268a7e2c821d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he083551ad54ebab4cfb39c7c78c4fe80a7db596a78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1638fe670c219296460b1b2c305107a3753f1d9f32d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h446ca806f1919eb8defb4dea8233052aaa65a11924;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h36775fe56e9b58385de2cfc93ff20fed68e2043703;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1387098dd161259805b1561bfe9baf02151babfd73a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13626bd2a8cd8e011e23ffbc1a9b5543a9fc8f94167;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14eaca180d532c862293b0457b38c18824e88beeb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h38fbdc300bf96230604878f7ae07c2ff3e80b50a05;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195701258c9525e4c2ed635dab8383c7bf65b734c8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108e4071e4ca626bd8413d46937c84b2a05fb582282;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h683faa6b8c2c38f6d93388ce91169bfb9c29665627;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c78e939d5a46ddc57be1d31e0b260463966f10a24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108e2dffb318405b7374555e2cd5ef72d78d4046a50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6424727668ed9c010b7a35b935590c02ddc5617336;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb8e2706bf640da63c6f5a63d1186797e7e65494fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a393a97de38719ff5f1e5488870c29b9d352fcf3ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5baa3fa93dd5684d62af844b69432425552aeeec29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h316150026c3798e04af5e024f6a1168f51409be134;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7264a1e1630cc09eb105b71e6885deeceaa3c76f98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha0a77a6d394cc033d4dbe432f20cf495683a972506;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc1309e3ad7d9781599bdffe582c19db59ad4f674ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ae54740a928c6ba286d37cc19a3a3b5f32b727054;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135069efd4b5a0e14dc3bd2de991465bcfa01625c05;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he290f6e554d1d63965488e0a29d1f4e1664f36ede7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f76ff18f9b33a584e0fcb01fd767a582d2d4e6e292;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18deff4d2c371f2d9025bad7e01b98a565055d1efe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h484c25e7177124e775504d909b2ce833d42274a416;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ca9b39679884226c04b414aa409c146702b7c4b3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141fe2ecf91deb4ad25a5ac61b19fbbb4878b20b57b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h731bdc3b0a290d675a2ab8705d79d48202d45af4e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14f822ac433a3712a95d3e299316261d36cab9bfb94;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d113f6d50ca8fa6c05a81076035bb228018cce1fe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf342b4860091d2b41ed882e46642d6df75b99283c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bbacffca2f42b50dfc84b5c11e57d443e72ee139a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be142043ab238ac20fe294418d1d882400eba7f757;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e576f9645af7578e7fb692e1a3e25cdad02f542516;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fff576fb980a72290ceb3296c0654e230c0d7cd465;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17761c5bb2214551250dd444c044a57fa2cebac54c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h152ec9a33e72de75aa94d7b93ddcc4cfaf18e38278c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10b727b5b70badb777e4429dcb9934abed4f966384a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb4363d7311cee6c82d7ad6b34f03c304348397d08e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb8adfb3b2fc0f659ec10248d9eea571bc94057597d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha026aa70f7198bdb93e29786798eb57087882cf6bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcab90e65dda3d5cebe7083df7f316ea09effd7d44e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e8ebd5d3c0b542377e1feb3e184ed0e0dd4021f63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h182fa22eba51d03972263810874e27a4dc4fe8e010c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11c1d3d84955b82ad1b5cb812c67471fe276db60c06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14a5e7547935c76a41ac0451fe16740a182d0d3aa1d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1311fe00eccc2c3466bb431074858ba248362e984de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14018fcc5ffa1be20eb6c3aa919d73dde489b172d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15dd788eaa31240468c4fac55cd6ff13634070e3161;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8d0404472ba71ae4a9f0e77d36aeb469b9134a103f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a279ac00247489cf43254b8d5dcc9662f96f1278f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e2f8080e156312127108fb79fcd892685536b7376;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1ed0bee10946cb72fbbd186438fddd533d2bcc178;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h73e10f89d60090f1de6d38778f4c546087e28e42db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h145a6fcd545462363c16aa6d3ac1442ce4e875b9147;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b7a739575c7c336d9f3f69ee1a8380a80a597006a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17365b1d3f7b84fca9fce1fc4730ac8a7cac540b8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1347d6c14d2a409fa4f714fdb748a0b3d55f975d36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1200dc43c86ed840e99e358c6fa61eb01bf726a9790;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175db953b0dd31a7ebd211af5ab35a2296e36973833;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h72d209b43e12f38fe3967104d66acbba593fb6e212;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118893fdfbd7f97f1c876b2f7e59676fdb288540c8a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12bb3c86b986c6db17240c2e45d79e0f985f1815c1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a987dedd4943488b72330eff7d1d76d03a177366e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7cc78e65dd9b6f61d4a509a70f7cf0cb545e5cfc9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17fc2b7a7ff47c01f549a6ba41862229c14079b670e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h248cedc558f126e214e18f65a969b8e446d0df0f75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5fdf4f74020658ee4418448504aa97553f4d8f41e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f4371ae709c54131a94906b437af6da7c8a4864359;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f652f7fab89406618dcc56c61f50873c16139932fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80c29b4e34c4e4fc21bcd8b3883280708c92ae3384;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110cadb0836b8d24081f7246ee5359ac8bd8604ea65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h23187e37b1098f412cba95d7683a502e7390eab6e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb8b4062e938cca6ec637ceb04f4301730244e0a26a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5002214bef031cf2961992135781310896864e17bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h274f28e0be43d617e24c952669185749d20e2bac7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1913b4edadd7116f040543b3ffb79a4aa142b399d4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15d4353d3de1c108c233a8be561faad60a43e2ff098;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc4c205a166687ba215bf0e673b17c611620fe9ec00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h129f7457d2bc79c95b4dce19b14c77bd924ed6eed27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a72e70bc231d6a9c615b4b5cc1e44a0c4db5eac38;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f2de0a6f8f3d02d6ad1850f653b8341758f26979e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6d46990e9015ca9794184f21d20e804c0c289f9b3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2fcf1880e9298d589105064a3f23aeafee03f9d465;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c48c1ea8e2f7d67315f4364e852d13dec41a2ffa5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h115a5d15dbd0f3185b07548b911355b257f881a386c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f40e62841eef5ac59a19797a0fee356a26b236bb1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af0695b0cefe8bca1b47e56f344d7944d5c41afaa4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd0ab68f198a1fa7e48538874ea8a578ca8330c1dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda88615a6f8e25660920b6f4e373030a84d2e1a298;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb0009dde87f4b9478c38be0c7883674ea6e0a6b2a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15996eb9aff968fc994e4551e6999ac638cc3148628;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1048299a38bcfbb27879600ce12a8fbd0d6a53ad131;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'had558ca766023e7d9ef4b84b3dd910639b18fafb0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81ebfe6c3b90fa9671b468651e91ec3a5d0cf2060a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148fc209cd1e7b2bd4f68fd906ba43685047900f933;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11040d89acc8731d30acacef8e87b7b16cf94a49131;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57651a2ecb801d12bc43ae27cd9ff9f6c802e974dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h90d8b2ef83ce5c4fbc0a4285d237d67df27183533c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166b0d7e0ecf9c222f3077f33aaa577a0066126fedf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e44a420bdeadb975582872d6b8c56cc52f96db4a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h404f46284ad4b605b856ab410597befd15a00e0d94;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h180566b69f46e9397ead9c3299720d9933938a5bdb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed6322fe69f01a6837fbef0611d65b628483f16bf9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfdaa536639c1f81299c644912bd1a90985187f5463;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h225333255adc0bc7ec8e03d176bdf1e7a120e4a3fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14dd27fa3aa800ad7d3032e8d59ca325807dee8d86d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he636f3f49fb834bb77dcff7fbeeaba4c751c905f52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137b46d0403035a6a91915452a39226fecc0f71db7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12383240cb23b77a62f4df6e2cedebf32f189b5c8a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6d3e50754fb463403bea21e704a9dd7834d13cf5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2e77103f2e9ff666658ff6e947167021a05a433c47;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14be7d618dc46f3bd4edb5bcb0815fa243599231e53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb28d8c91711b7133ac77a9277f1e9826fec5e8d9f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8ce00cf909b97af14f70c190a7c823a375fe7a633;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0360e44ef83ccd9f5bf0b6b5a0e422095e0833ec5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c70d25f6e7b9068a088b27c9a7ad42bd7e8df697c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbcf3306db1d6e46c246b0d8d3a8d044e1dfb47e7bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157121a1e646d405aa992c0cdff768e215298d47fb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafff2951ea35f1e87159d5cdce0fdfe8477347d7d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h189172593a44ad79a55e368c1c00fdda2b765145090;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1051834eea053f06f2aede199d39d849e4b8119858f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha54679dd97a3d3a1ddb395c3610312f48391cf5dbc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hefcbb7e7d341ff88a96c5a5d65eec5bea6bd0ed0cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ece142af5df0f2b3647823b9a40d26accc79896488;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h209690f3c452312652855beefac56a1e97e7a3059f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f10d4c1986eb873beee6c876dc8d662c8da229b93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17588f2b91057a3a00d9b77ff3ae50790a15dcad083;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2a1c530a675c6ac19611e2ff04bb1226bad44b6ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he92caabc304b842759dfca06991ae6daeaf31b562c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f4009ac90f90977c245476ed4740e262727b7a23d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1233c79381afbf50cecdf880c3edc3ef4e070e84c35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ae381d8ad3cd3c85cb233b67008d0b3902c1f6d189;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ce83a9d324fa200feaf60453ee39dbbfac9ea5fef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d55e80697adaee5a09504d4f8335ba639d5acada5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52d04608111e5551eb1270de59dc7d0d705098b1df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ca9593c3fc45a9f56b9dd988364a369eac8ad84e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18904e2f38fa8746d7bf4e52f24a0f6cf89d64fdab5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h412c88e4ef69635a2409a590880328bdd5632bcea5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1108b9144cdad192dda38b845511348b6b8b134aed5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153def90fbda1e8b33ffbba399cd6e444202fedb5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9d9f49ab32814967dae48e78b44ff376b56b468dbd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf79d944664e009778c56dd8310aeb209cf18f1c361;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc317219430a41d24027a9c38dcdaed987894cce459;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ac84ad21f59b224fa6fc78de565524bc5426ecbbe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf919cf1e553546cf6011201aac63e665624fb44e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1202fec54576baadd579a38a455dc02adafbfe2ed17;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132496ef1f73fc0f3339b9ca414055bf8074dce5fce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13faf722dd4c5d431feca97235d2a6ab24ff91dc454;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c953aedcab9499058ed6dee3e1e05745bdf7bdfde4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c5eda7a0c7c3c1475f99b8e47efe70d60d4a7d12b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ad2262be20a790a3c48140ac189ac12cdc3928ad3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc1790f3fd7ca0a771a230752e00fd193ee7d1920d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffeaf69813971be5358b880bd6cdf15a4a803c72a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113f5ea6840ff5194cc8628837b621d057baf48d0e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c2214baddd5345d92973374d785843f387b95264b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4511d5fd13feac8e269cf8b91a491a821a3d027141;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heaafd42fb7c6e0ecc197f70505d0895cf5872c183d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8a25dbc03e776a0ce04b8e86750121bbcdfb2a76a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h875cc345252662842ef4bc619548c62d6e7069ad22;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa0f6e5068bfb5326426696d401fbab6048d21b423;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18fffe44351ecf4fb9697855f88814b8a392762f699;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a949cee90d1a6807a8fe4aec8cb9e61718c5527fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a534157ae8db1ab873331d8b4caabe804e44c954ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h260656344a54a1b12cb45eb0aeaf3716f346761005;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h173e11d3e8fce609ed2ac672798e288684a39040b62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h105cd3f85b9a7dcbfbfe18e6c625fe2a78948c7108a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h285679f1ba06cd457305d13019188737ebe5a7904b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfffe32ad2b87461319624712f9d87982fd9ea2131c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha5dccea544d78b969d2d5abe528ff96603b653049;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11ad5cc3a9902a445214936ddc026efb93b983fd633;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198d4e4b9b9316d2cc76ef083fa72e16d842ba861a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h23526badaf8d1239e2607fa2e956c530545768e4b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfa0654e1aa98b06f48922102e4951710c26a6e03ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141fe806c1a69bf83b3dbee21fc80a51361e6f953c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha90285da01f0bc1842736a0833d77e36458e5b24e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cfb325aa68e29d25e5a427e7d8c57718e1e93c0f00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hef8f74ca20b5b51ea956457595a906ddcfa7d88fb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f83b1d844e040e71be8d934611f3f6add2c0ccedae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e67376df13265193023753212e1bcefe5be1eb5c4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3b10aab37e13cb213266e10f8d659be6ca1ffc59e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdff94a1191c1fedec43e3e54016905620fb6e0d721;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10faa25d13cc999064254b84aa61493a65d0798b746;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6f636c8b557828c8d322a790a4fc2bfe912729055;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169bfedb4ab44a1cec3733a2735f6b13d9042ad1b3e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h170ea69bee8d0e8a0090793a3fc3e9419324e81fd62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14ca547cc8ec082a17f9e77f5efe8e0662278de55de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbfa7532ec3440bf4c2ac2e72232f120f482aa009ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea8050f2261289b5055709ac2f4ffa0dfb9bd6c397;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0dd806a286b76915de49d023afff26ebdb013d998;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h682db1f615b4d23d20c705b9c3bb7fa89d39a54ed7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heaffa3eab3290181a67e07d26eabbb2544cbf4c926;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h186f2fb92fc92702fe39558d33de622dba08012a4ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c95a1ca73b99353e55b0aad6be9a26de813cd288;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7f9b2c714927e638608e71c4e98777ef91a9473ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3d0462b0e308e69b64ca9dd5d1759a71f41e930a02;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d3299b43589e1e2fe60afb04966e8427db9791e45b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h153e7104317f9d16f54e1699437cac302192314e5f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1277bef43a85919567177dc5919c14bd2183cd7ec26;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11855e5d03b1a4579ac2de4fa7846502245c531a4dc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192936d9844fc8705f4a630837033c40aa211a4950c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11bc0a4990346518c3e5404f425c46028018566cf2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108296f11ce60d8a0d0894ace7054825a99bfb1ef53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc9aa21fb56917ac409b9a129ca599a988edc7b9c8f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc6360b6f0ad80b9a749654db3a9d5ca01fb0a21605;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b7597f290c1900789ad9c3fd255c95b9850f183ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89183f08d6802044ff22c9f2027df64a3e528003a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h155587078f78fee48709856ea111e38761033664dcc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ed6605550e1b14c0fb3cc4c344287e3d0bfe036c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a0e46b8874dbf9126bdbf385f11453c2e08df0add;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0d8d824e011a1a6a41131ba177b7d53332eb8948;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16122b64a2774017a658658bb97f902d99e6ea81afc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17066c8e6c2e6e19a9750b996701d37dc2d33b5eba1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1ce7f7c255d02af89fe85c313f0250bccbbdc30f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h160d103ae0206e4f6d686fcf6050c43b4319ba43ce3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2fc7f5c24879a2e706c0c94988e23d4d79b3e004b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137eb9e0e5f58e47200ed5a283692823a176bed50a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h45c40438de9029c4e89944c88c59aa00b94cb4c6ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h219f5887866fa418af5c68a49dabfa1016d6dac915;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197f49d9d2d8e450dfa6db2ee93b14b7aa69df21b7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147262b67ac2d2259a565ae59ca53c83a73bb06dd6b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h60166920c3a9c72539f10ac3db36b2465e4de6e11b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf1bcda07ef04a1d5f933a7b076c7301ae64d984190;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bccae02b4338711979d86e77aaf8371e8120f8cb98;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h180a06cf1e8e4acef1bb01efbb1e2122e55d3f668eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ee948d8ec9e037c060be2e6996fcf17c47e230e53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4cf800000068a9e2c543040e6f6d79bb490dffac00;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h88a27584a7b0984adefb0b84b77fb6cc65596e0aa9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h37c7e2d644e769afd20d87cccbc3f4bdb8b3a24817;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hffbfb0151b40919376d177090a81fb3ef2af08105f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dfae1374f7948a32d24d6eaf7a2d51777dc30de586;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b6cebf6bb8bdcfc326372098777c14504042f41c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h935e0cef9fcc2284b9c6681e400a3186e0707773c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dbfeeb60ff10d3c8414290b2efca112782c43b7287;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h179eb376db1ce39b56ed9251b57fd0fbc804dd6153c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h70d4a1cd798feacbdef5cf223a7cace861bc6db2b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc303d9eb9148954ce8741742cd619b126fd0bdd0f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf5c4e9baefb98d512b985d1ecf5b9c3ff2e5211813;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h772d35b3156585cc34048a037ebba5303f86e5917c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h894eea6631d590878ad6912a1518f287a70ced5d01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hccb2ed97b2c02130d40c673ec22b3570b68feec912;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6181c4ae38261fc1942560b0cd5e0289a3ef4780a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cf973f5965ebde51473281a0f3e18a90b751e39ce4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b8cd8912315c523e3ff68b835b01c0ac8141b944d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h481d12878153009d85017edbbeb40c7761f49d2635;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11af6b84f46c13c39678c6853bb7bfeba4d7cb4e564;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16fdf447b59b62a1e405d50a075d9d17c2e18e418c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf6200b4bcd2bbe39290e6433c84602eecc0f8b1ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1903191187fb4ec8310b9cd742f6bd5e3752fd6d3ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141fbe266727e9198112d3fbc420330de99ea2919b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3ba84fbb7a2728b0f36ed2f92937ea2c1fb0f07b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1211daed30bb43be2cce7ff61ecd1239f01dde2176b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ca71943adadbf25df6ce8d9f1150c0c8168967999;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c03f382b89c424038aecd72f65c497603cc756f65c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h71421869e3b7de68620e237e64726293545f761395;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12456d7f339271196b090989400bbb219f637a21165;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19394e3e47d3b72a9579f6d7299dda262d935d81ea0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9da36822eac81b47473b2ef3608245da912b43926;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h341334353c60625186ead81e1c60cd98f06d699528;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h71ff7e97acd4a0c7c14e26ee91292936a073b0beea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h159df9b88108b46bc7c9f0dd5930c1c45290904f507;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h151401bb96110bac25ca36b44e1b1a8234da89ba91;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14f5db7f192db3d9a2e5a27b12274f70ebc0b2e2d08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9c3e4d2522043ea10f1b363065a870d0a52815ad7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16803c7a077962d1da70ad8c4e54826bec41339c647;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf7c0017b15f887b0caef0f8b7565acc7866a5e740;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a3eee0cd164804da3e0da2fd1660b693bfcb301c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb31a9955e785feab019fdcc17e4f4c08682e7c5b93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h297edee8620452dd9c1320c97d94cd7a7debba2277;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbda883ac7156c828f51169e3d1ed5b49cd7221048d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c3ccfd8f7533254d0e3091c0304a77c5cd96034e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h124af4d35bc6a31f177759c93c4672b074076a7f01c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4941359d1101603ea9e8fc6fdea6b007c92c84d7a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126e0cc35efc8ac4cbf21989e47c8dd17f6e627b625;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18486e65d7e3371af4221e609482b7f1a2b7fcf545;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e9c04b95ae21eb30e6a8965b6785569a0935fe236;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ad3002a738d892aed36beb7da52590c6a4cf3d6d25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h881523ca3ced5d5731c427abfa0af9c7a0ff9872a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h51c411bf2875dfcbb17c5fd4ee5d7263e5d9523afd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5a962229d1c9310882e5ed20df9d0ccaa213129aec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4089e80fb91eef434aba5987c0e06e641512bc0b27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9602ba04047301a92af97d14feacbf40a5f8530a9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha531b414ee21fd0da49df4c2fb18bf043ac585e94e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb03bb8286e5fe4e38e1559e06d1dac3bd3c2a65178;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13c87b1584505a03ed5ca14931feec2dca85ae362d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5880b5115132a0e9c851c73dff5502786492e8ebdf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1522b436797e2d7b64b82dc0bc4b6a8d68fb2f0f48d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81284c537369733efd70d7003f0e549ec69eea6dd1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b5e036a4e83842124fa79cfdeab9e8d53bca2d3777;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1849a418234859a0019808350de8ac2cfa78dcd85a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h581c5e859416b51aece28d7abd01cba24c446b41e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7fe948b857ff4b03a4a1f7633dd13652d3d2a624cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7015fabea1f47700f0694c0e3535dd88c1fa4d6530;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfa7e86e2db481f4027c2fb7cdb54ecbaf30a548e46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h64c76c3638e128c3f2fe4562004dd9d25e9939ba91;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he27f3252d286f27badcadc7dac9ecc0913ab5920b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1daf94bed919d7148357fe2cb5db606784ca2eb0823;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd2d32076b6bb2ef0d3b551d33049767d00a9f9230a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d42e056a63d810a9bd13abdce817deb9ab0070546c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hca0b547a1010b54575e3c43fd8dac7dbe6478299c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e409c33998c1d9349920f9c761f4ecba6921c2b27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha0f3a2157c28a7e8aabe133a9463dcf1ac872b7cce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1342e87a1852b8acc778865074c947e84e87f621543;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ad7d5733c916350df70f96ac9360185181aad707cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd8748994681064279e7ad599a6d4dc4bdd81d0f57;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a316d43421a96073e43e676ac89a0d99786b8f4784;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82d9f38a60151fd20179d33d4196a2d4ebb5c00c2d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1619bc5de55a5e170eb0b4d9690cf3e466d7357d26b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h468842bb75b520b736ae9de1644db3a9e53deef69d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he75f07f89d4a3060d6ff4138f634474209dea4d021;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1237e7bf84b9b7c2ea7e3943dd37a1f4c056cf4e676;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h160c3a4faa398b6de6ed0b148d873147e80a1e34947;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1079d6aa6d657a6a9805c17d59a8f73694de31c37d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b48942111a81529f2737047868779a2b93400d48b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8e79380a47136fba8ef5e011a12da0acc2bed7f492;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d2af477e98e76e429e39ebe5f9c6ca2396088b1ad;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5b6d6e1303b698f2ccc06907cc908b56ca70ce08e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he94fb574b1e5e771f477744b1c1a1b33296c2fbdc7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19c1b0bc8f8edc00ffabb0a035bd2857c815a696a71;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1ec8f7af7957ec1e773feacef7e3221dab09ebe0d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h43d069619d7873876018153e7fddc1baadec84d2c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a2d16bf52fa8bac809eab95ef8c068b5132a132429;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b92f239d28896f1b54bfb0220961418d86a63b8c93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57c53aeb3ac1c87a5807769f2aee08b44ac4b377b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c8e223115344226a4a42f15996d1dcd9b6ab3d391f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63ce535f0b211aed2209e5b70aa22356b3b4afe187;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c6d08d0211975d11ff26e7edff5653342288842af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac98fd020326ee7689df3b6fb022e7a8ce8b8ba07a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17ebedc30a91a8fc152a9052dca091f0eb16b22c858;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h158abb3ea8195f5110c28f8d75f5b7d44f374f47f7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14bdf2e98a47eb6f1ac6d1288846a4bdcac6d35aeda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1173ff3ae42178c6ef684fddeb5a1568db73ba254ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d642b20760494ed579c551bd1fd21f5694b87c42df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h127d10b808781b3d46fe91e92fe3af0b026bfdd83ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf250cc6d30142bc50c75c6027a449ab3f10a31cb4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7644d16af1a29ffb323b25f0b5f1ff830640f08ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2981ad5664494bde86b108bf0215099e18bc8372ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174bbddac5cdbd924121bdeebc85a6d786aa04fd500;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4dd841d97128af7bdc1335c31b74230d3b59a55b80;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3c9208a0744c693f93c39bf86930a3f6a25d15913;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57bb1f2bd9a69e45b2faef8a9bd9906388e4baead0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h923ebd96dad99cad13735d20e857742aa63dcef577;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha635381db5eb2c2d39afc51c1f88b11cf661d82155;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b9c5e1525ddc3f218f7d6d555440d31e76c9573f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2be5af32101f9ed4b82e99c637e716e1a3a417b8de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18e5e26f038d2d6b4d364fdda54031334bc724f73b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147852fc46154d29ffdcb57a495dde6c54b993f269a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1312a148ffdfab923a5f53f9f656228d5b2c8f0242b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1344a2f45fea2a4a53a064c9974bd69ad4567fbab72;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf47fde1415942a6fca3ae1ecc3a9ad91c1fba811da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b21ae4efb38381e8a24a65e15eb98035fb66c6e4c6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3fb2f8b52404cde0d86003d6b2327db47470ef859;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4057934fad09d954bce01bf203529ca116d2a563e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140cac5c75cf2f3a50851dcc2818a4544526f54041b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcda303b0faba16bc2da8cae661d091d7753cb2f71e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e0589518e79d023c885b1e8f535912eb72d8bf93f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcf6ebcee497b03a2f49a3e2530a5ec5afe21955906;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f461590ed04473d775586de73a6d8600a2daf2cc16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e7d148d56b5f8a59b822e62bfe85cf67e52674b4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3f380f2005ea70062361a8222f208137918035c95d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d0e24a32066e59fea7335c6e17d3895843eb064feb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f8d121608c93650aa79a52e2ea74474c6a10b779de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac01919532a4291300897ce50d29e68266a4787d5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6ae9010f2062ef6c2df72bb102bdd06be5c4db117;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3555df645a521c4243839722d5fcb00cf0a910a63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he686823b1399a2d8505e1520ba4490167344bd6510;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1115ec4e19f9532820c076a391bb83862f71e22b5d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5125f077e4e2c7570b830c21db89155efa101498cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e625fbf3361189ea1eaf36ab8d7b977ea7e4296c29;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a45cdb6dcf7a4230746abe81e195771aa2c60a213;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb30992718b8cf6b3a7f77294dd512638cc9776fc6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c52497af0eeae4f8e50d9e2a64f26b3a85743186cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h189189d5f8aaf69b2c25c4893147a9d31eec1052f79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11e72055c53e217055ed865f333496b2a1485cee420;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a7914245b82eb7005a5926be48145c115d3efd62f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd19860c56d5f8ed3a4e59e86acff3153e6cd23aa6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39950ace1a850da0287aefa35356b14d61d85f21fb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13e0105441ae96aa832870b364a2151ca41dbc2b60c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ba1adfc591d42651000cab802d854ad812bef1abf6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a1818ee8308458bd34e812133e38886ef01f6484c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a0bbaf0700e126cc56fd9223724fe6475716ec90d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h107d300381bedbf333501369b441191e56a80c424c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f791416c0916cee83a85b8e83e66d62e061c476db4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10838b61b8087f010eaa57a40c7f3a8245213683401;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8151f434674099e2516b439e806066d26201ca6222;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed3254676746caf7263254529b77a953bc4497da5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195f59d510f2f8173d79247c931cc6b082b03028e5a;
        #1
        $finish();
    end
endmodule
