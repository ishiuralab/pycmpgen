module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19);
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    compressor_CLA16_16 compressor_CLA16_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19));
    initial begin
        src0 <= 16'h0;
        src1 <= 16'h0;
        src2 <= 16'h0;
        src3 <= 16'h0;
        src4 <= 16'h0;
        src5 <= 16'h0;
        src6 <= 16'h0;
        src7 <= 16'h0;
        src8 <= 16'h0;
        src9 <= 16'h0;
        src10 <= 16'h0;
        src11 <= 16'h0;
        src12 <= 16'h0;
        src13 <= 16'h0;
        src14 <= 16'h0;
        src15 <= 16'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA16_16(
    input [15:0]src0,
    input [15:0]src1,
    input [15:0]src2,
    input [15:0]src3,
    input [15:0]src4,
    input [15:0]src5,
    input [15:0]src6,
    input [15:0]src7,
    input [15:0]src8,
    input [15:0]src9,
    input [15:0]src10,
    input [15:0]src11,
    input [15:0]src12,
    input [15:0]src13,
    input [15:0]src14,
    input [15:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [0:0] comp_out19;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [15:0] src0,
      input wire [15:0] src1,
      input wire [15:0] src2,
      input wire [15:0] src3,
      input wire [15:0] src4,
      input wire [15:0] src5,
      input wire [15:0] src6,
      input wire [15:0] src7,
      input wire [15:0] src8,
      input wire [15:0] src9,
      input wire [15:0] src10,
      input wire [15:0] src11,
      input wire [15:0] src12,
      input wire [15:0] src13,
      input wire [15:0] src14,
      input wire [15:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [0:0] dst19);

   wire [15:0] stage0_0;
   wire [15:0] stage0_1;
   wire [15:0] stage0_2;
   wire [15:0] stage0_3;
   wire [15:0] stage0_4;
   wire [15:0] stage0_5;
   wire [15:0] stage0_6;
   wire [15:0] stage0_7;
   wire [15:0] stage0_8;
   wire [15:0] stage0_9;
   wire [15:0] stage0_10;
   wire [15:0] stage0_11;
   wire [15:0] stage0_12;
   wire [15:0] stage0_13;
   wire [15:0] stage0_14;
   wire [15:0] stage0_15;
   wire [11:0] stage1_0;
   wire [8:0] stage1_1;
   wire [11:0] stage1_2;
   wire [8:0] stage1_3;
   wire [5:0] stage1_4;
   wire [5:0] stage1_5;
   wire [5:0] stage1_6;
   wire [13:0] stage1_7;
   wire [5:0] stage1_8;
   wire [9:0] stage1_9;
   wire [5:0] stage1_10;
   wire [8:0] stage1_11;
   wire [6:0] stage1_12;
   wire [6:0] stage1_13;
   wire [12:0] stage1_14;
   wire [7:0] stage1_15;
   wire [2:0] stage1_16;
   wire [1:0] stage1_17;
   wire [1:0] stage2_0;
   wire [5:0] stage2_1;
   wire [2:0] stage2_2;
   wire [5:0] stage2_3;
   wire [3:0] stage2_4;
   wire [2:0] stage2_5;
   wire [1:0] stage2_6;
   wire [4:0] stage2_7;
   wire [3:0] stage2_8;
   wire [6:0] stage2_9;
   wire [1:0] stage2_10;
   wire [5:0] stage2_11;
   wire [4:0] stage2_12;
   wire [1:0] stage2_13;
   wire [3:0] stage2_14;
   wire [3:0] stage2_15;
   wire [3:0] stage2_16;
   wire [1:0] stage2_17;
   wire [1:0] stage2_18;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [0:0] stage3_2;
   wire [1:0] stage3_3;
   wire [1:0] stage3_4;
   wire [1:0] stage3_5;
   wire [1:0] stage3_6;
   wire [1:0] stage3_7;
   wire [1:0] stage3_8;
   wire [1:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [1:0] stage3_13;
   wire [1:0] stage3_14;
   wire [1:0] stage3_15;
   wire [1:0] stage3_16;
   wire [1:0] stage3_17;
   wire [1:0] stage3_18;
   wire [0:0] stage3_19;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage3_0;
   assign dst1 = stage3_1;
   assign dst2 = stage3_2;
   assign dst3 = stage3_3;
   assign dst4 = stage3_4;
   assign dst5 = stage3_5;
   assign dst6 = stage3_6;
   assign dst7 = stage3_7;
   assign dst8 = stage3_8;
   assign dst9 = stage3_9;
   assign dst10 = stage3_10;
   assign dst11 = stage3_11;
   assign dst12 = stage3_12;
   assign dst13 = stage3_13;
   assign dst14 = stage3_14;
   assign dst15 = stage3_15;
   assign dst16 = stage3_16;
   assign dst17 = stage3_17;
   assign dst18 = stage3_18;
   assign dst19 = stage3_19;

   gpc135_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc606_5 gpc1 (
      {stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3], stage0_3[4], stage0_3[5]},
      {stage1_5[0],stage1_4[0],stage1_3[1],stage1_2[1],stage1_1[1]}
   );
   gpc606_5 gpc2 (
      {stage0_2[1], stage0_2[2], stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[1],stage1_4[1],stage1_3[2],stage1_2[2]}
   );
   gpc615_5 gpc3 (
      {stage0_3[6], stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10]},
      {stage0_4[6]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[2],stage1_4[2],stage1_3[3]}
   );
   gpc1343_5 gpc4 (
      {stage0_4[7], stage0_4[8], stage0_4[9]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9]},
      {stage0_6[0], stage0_6[1], stage0_6[2]},
      {stage0_7[0]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[3],stage1_4[3]}
   );
   gpc615_5 gpc5 (
      {stage0_4[10], stage0_4[11], stage0_4[12], stage0_4[13], stage0_4[14]},
      {stage0_5[10]},
      {stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6], stage0_6[7], stage0_6[8]},
      {stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[4],stage1_4[4]}
   );
   gpc1325_5 gpc6 (
      {stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15]},
      {stage0_6[9], stage0_6[10]},
      {stage0_7[1], stage0_7[2], stage0_7[3]},
      {stage0_8[0]},
      {stage1_9[0],stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[5]}
   );
   gpc615_5 gpc7 (
      {stage0_6[11], stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15]},
      {stage0_7[4]},
      {stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5], stage0_8[6]},
      {stage1_10[0],stage1_9[1],stage1_8[3],stage1_7[4],stage1_6[5]}
   );
   gpc1343_5 gpc8 (
      {stage0_7[5], stage0_7[6], stage0_7[7]},
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10]},
      {stage0_9[0], stage0_9[1], stage0_9[2]},
      {stage0_10[0]},
      {stage1_11[0],stage1_10[1],stage1_9[2],stage1_8[4],stage1_7[5]}
   );
   gpc1415_5 gpc9 (
      {stage0_8[11], stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15]},
      {stage0_9[3]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4]},
      {stage0_11[0]},
      {stage1_12[0],stage1_11[1],stage1_10[2],stage1_9[3],stage1_8[5]}
   );
   gpc2135_5 gpc10 (
      {stage0_9[4], stage0_9[5], stage0_9[6], stage0_9[7], stage0_9[8]},
      {stage0_10[5], stage0_10[6], stage0_10[7]},
      {stage0_11[1]},
      {stage0_12[0], stage0_12[1]},
      {stage1_13[0],stage1_12[1],stage1_11[2],stage1_10[3],stage1_9[4]}
   );
   gpc623_5 gpc11 (
      {stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage0_10[8], stage0_10[9]},
      {stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7]},
      {stage1_13[1],stage1_12[2],stage1_11[3],stage1_10[4],stage1_9[5]}
   );
   gpc606_5 gpc12 (
      {stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15]},
      {stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5], stage0_12[6], stage0_12[7]},
      {stage1_14[0],stage1_13[2],stage1_12[3],stage1_11[4],stage1_10[5]}
   );
   gpc615_5 gpc13 (
      {stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12]},
      {stage0_12[8]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[1],stage1_13[3],stage1_12[4],stage1_11[5]}
   );
   gpc606_5 gpc14 (
      {stage0_12[9], stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13], stage0_12[14]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[2],stage1_13[4],stage1_12[5]}
   );
   gpc615_5 gpc15 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10]},
      {stage0_14[6]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[1],stage1_15[2],stage1_14[3],stage1_13[5]}
   );
   gpc615_5 gpc16 (
      {stage0_13[11], stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15]},
      {stage0_14[7]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[2],stage1_15[3],stage1_14[4],stage1_13[6]}
   );
   gpc1_1 gpc17 (
      {stage0_0[5]},
      {stage1_0[1]}
   );
   gpc1_1 gpc18 (
      {stage0_0[6]},
      {stage1_0[2]}
   );
   gpc1_1 gpc19 (
      {stage0_0[7]},
      {stage1_0[3]}
   );
   gpc1_1 gpc20 (
      {stage0_0[8]},
      {stage1_0[4]}
   );
   gpc1_1 gpc21 (
      {stage0_0[9]},
      {stage1_0[5]}
   );
   gpc1_1 gpc22 (
      {stage0_0[10]},
      {stage1_0[6]}
   );
   gpc1_1 gpc23 (
      {stage0_0[11]},
      {stage1_0[7]}
   );
   gpc1_1 gpc24 (
      {stage0_0[12]},
      {stage1_0[8]}
   );
   gpc1_1 gpc25 (
      {stage0_0[13]},
      {stage1_0[9]}
   );
   gpc1_1 gpc26 (
      {stage0_0[14]},
      {stage1_0[10]}
   );
   gpc1_1 gpc27 (
      {stage0_0[15]},
      {stage1_0[11]}
   );
   gpc1_1 gpc28 (
      {stage0_1[9]},
      {stage1_1[2]}
   );
   gpc1_1 gpc29 (
      {stage0_1[10]},
      {stage1_1[3]}
   );
   gpc1_1 gpc30 (
      {stage0_1[11]},
      {stage1_1[4]}
   );
   gpc1_1 gpc31 (
      {stage0_1[12]},
      {stage1_1[5]}
   );
   gpc1_1 gpc32 (
      {stage0_1[13]},
      {stage1_1[6]}
   );
   gpc1_1 gpc33 (
      {stage0_1[14]},
      {stage1_1[7]}
   );
   gpc1_1 gpc34 (
      {stage0_1[15]},
      {stage1_1[8]}
   );
   gpc1_1 gpc35 (
      {stage0_2[7]},
      {stage1_2[3]}
   );
   gpc1_1 gpc36 (
      {stage0_2[8]},
      {stage1_2[4]}
   );
   gpc1_1 gpc37 (
      {stage0_2[9]},
      {stage1_2[5]}
   );
   gpc1_1 gpc38 (
      {stage0_2[10]},
      {stage1_2[6]}
   );
   gpc1_1 gpc39 (
      {stage0_2[11]},
      {stage1_2[7]}
   );
   gpc1_1 gpc40 (
      {stage0_2[12]},
      {stage1_2[8]}
   );
   gpc1_1 gpc41 (
      {stage0_2[13]},
      {stage1_2[9]}
   );
   gpc1_1 gpc42 (
      {stage0_2[14]},
      {stage1_2[10]}
   );
   gpc1_1 gpc43 (
      {stage0_2[15]},
      {stage1_2[11]}
   );
   gpc1_1 gpc44 (
      {stage0_3[11]},
      {stage1_3[4]}
   );
   gpc1_1 gpc45 (
      {stage0_3[12]},
      {stage1_3[5]}
   );
   gpc1_1 gpc46 (
      {stage0_3[13]},
      {stage1_3[6]}
   );
   gpc1_1 gpc47 (
      {stage0_3[14]},
      {stage1_3[7]}
   );
   gpc1_1 gpc48 (
      {stage0_3[15]},
      {stage1_3[8]}
   );
   gpc1_1 gpc49 (
      {stage0_4[15]},
      {stage1_4[5]}
   );
   gpc1_1 gpc50 (
      {stage0_7[8]},
      {stage1_7[6]}
   );
   gpc1_1 gpc51 (
      {stage0_7[9]},
      {stage1_7[7]}
   );
   gpc1_1 gpc52 (
      {stage0_7[10]},
      {stage1_7[8]}
   );
   gpc1_1 gpc53 (
      {stage0_7[11]},
      {stage1_7[9]}
   );
   gpc1_1 gpc54 (
      {stage0_7[12]},
      {stage1_7[10]}
   );
   gpc1_1 gpc55 (
      {stage0_7[13]},
      {stage1_7[11]}
   );
   gpc1_1 gpc56 (
      {stage0_7[14]},
      {stage1_7[12]}
   );
   gpc1_1 gpc57 (
      {stage0_7[15]},
      {stage1_7[13]}
   );
   gpc1_1 gpc58 (
      {stage0_9[12]},
      {stage1_9[6]}
   );
   gpc1_1 gpc59 (
      {stage0_9[13]},
      {stage1_9[7]}
   );
   gpc1_1 gpc60 (
      {stage0_9[14]},
      {stage1_9[8]}
   );
   gpc1_1 gpc61 (
      {stage0_9[15]},
      {stage1_9[9]}
   );
   gpc1_1 gpc62 (
      {stage0_11[13]},
      {stage1_11[6]}
   );
   gpc1_1 gpc63 (
      {stage0_11[14]},
      {stage1_11[7]}
   );
   gpc1_1 gpc64 (
      {stage0_11[15]},
      {stage1_11[8]}
   );
   gpc1_1 gpc65 (
      {stage0_12[15]},
      {stage1_12[6]}
   );
   gpc1_1 gpc66 (
      {stage0_14[8]},
      {stage1_14[5]}
   );
   gpc1_1 gpc67 (
      {stage0_14[9]},
      {stage1_14[6]}
   );
   gpc1_1 gpc68 (
      {stage0_14[10]},
      {stage1_14[7]}
   );
   gpc1_1 gpc69 (
      {stage0_14[11]},
      {stage1_14[8]}
   );
   gpc1_1 gpc70 (
      {stage0_14[12]},
      {stage1_14[9]}
   );
   gpc1_1 gpc71 (
      {stage0_14[13]},
      {stage1_14[10]}
   );
   gpc1_1 gpc72 (
      {stage0_14[14]},
      {stage1_14[11]}
   );
   gpc1_1 gpc73 (
      {stage0_14[15]},
      {stage1_14[12]}
   );
   gpc1_1 gpc74 (
      {stage0_15[12]},
      {stage1_15[4]}
   );
   gpc1_1 gpc75 (
      {stage0_15[13]},
      {stage1_15[5]}
   );
   gpc1_1 gpc76 (
      {stage0_15[14]},
      {stage1_15[6]}
   );
   gpc1_1 gpc77 (
      {stage0_15[15]},
      {stage1_15[7]}
   );
   gpc606_5 gpc78 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc79 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc606_5 gpc80 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc81 (
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[1],stage2_4[3]}
   );
   gpc606_5 gpc82 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[1],stage2_6[1],stage2_5[2]}
   );
   gpc606_5 gpc83 (
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[2]}
   );
   gpc606_5 gpc84 (
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[1],stage2_9[2],stage2_8[3]}
   );
   gpc606_5 gpc85 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[0],stage2_13[0],stage2_12[1],stage2_11[2]}
   );
   gpc615_5 gpc86 (
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4]},
      {stage1_13[6]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[1],stage2_14[1],stage2_13[1],stage2_12[2]}
   );
   gpc2135_5 gpc87 (
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10]},
      {stage1_15[0], stage1_15[1], stage1_15[2]},
      {stage1_16[0]},
      {stage1_17[0], stage1_17[1]},
      {stage2_18[0],stage2_17[0],stage2_16[1],stage2_15[2],stage2_14[2]}
   );
   gpc1163_5 gpc88 (
      {stage1_14[11], stage1_14[12], 1'b0},
      {stage1_15[3], stage1_15[4], stage1_15[5], stage1_15[6], stage1_15[7], 1'b0},
      {stage1_16[1]},
      {1'b0},
      {stage2_18[1],stage2_17[1],stage2_16[2],stage2_15[3],stage2_14[3]}
   );
   gpc1_1 gpc89 (
      {stage1_1[6]},
      {stage2_1[3]}
   );
   gpc1_1 gpc90 (
      {stage1_1[7]},
      {stage2_1[4]}
   );
   gpc1_1 gpc91 (
      {stage1_1[8]},
      {stage2_1[5]}
   );
   gpc1_1 gpc92 (
      {stage1_3[6]},
      {stage2_3[3]}
   );
   gpc1_1 gpc93 (
      {stage1_3[7]},
      {stage2_3[4]}
   );
   gpc1_1 gpc94 (
      {stage1_3[8]},
      {stage2_3[5]}
   );
   gpc1_1 gpc95 (
      {stage1_7[12]},
      {stage2_7[3]}
   );
   gpc1_1 gpc96 (
      {stage1_7[13]},
      {stage2_7[4]}
   );
   gpc1_1 gpc97 (
      {stage1_9[6]},
      {stage2_9[3]}
   );
   gpc1_1 gpc98 (
      {stage1_9[7]},
      {stage2_9[4]}
   );
   gpc1_1 gpc99 (
      {stage1_9[8]},
      {stage2_9[5]}
   );
   gpc1_1 gpc100 (
      {stage1_9[9]},
      {stage2_9[6]}
   );
   gpc1_1 gpc101 (
      {stage1_11[6]},
      {stage2_11[3]}
   );
   gpc1_1 gpc102 (
      {stage1_11[7]},
      {stage2_11[4]}
   );
   gpc1_1 gpc103 (
      {stage1_11[8]},
      {stage2_11[5]}
   );
   gpc1_1 gpc104 (
      {stage1_12[5]},
      {stage2_12[3]}
   );
   gpc1_1 gpc105 (
      {stage1_12[6]},
      {stage2_12[4]}
   );
   gpc1_1 gpc106 (
      {stage1_16[2]},
      {stage2_16[3]}
   );
   gpc2135_5 gpc107 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4]},
      {stage2_2[0], stage2_2[1], stage2_2[2]},
      {stage2_3[0]},
      {stage2_4[0], stage2_4[1]},
      {stage3_5[0],stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0]}
   );
   gpc1325_5 gpc108 (
      {stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage2_4[2], stage2_4[3]},
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[1],stage3_4[1],stage3_3[1]}
   );
   gpc2135_5 gpc109 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4]},
      {stage2_8[0], stage2_8[1], stage2_8[2]},
      {stage2_9[0]},
      {stage2_10[0], stage2_10[1]},
      {stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[1]}
   );
   gpc606_5 gpc110 (
      {stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[0],stage3_11[1],stage3_10[1],stage3_9[1]}
   );
   gpc1325_5 gpc111 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4]},
      {stage2_13[0], stage2_13[1]},
      {stage2_14[0], stage2_14[1], stage2_14[2]},
      {stage2_15[0]},
      {stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[1],stage3_12[1]}
   );
   gpc1163_5 gpc112 (
      {stage2_15[1], stage2_15[2], stage2_15[3]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], 1'b0, 1'b0},
      {stage2_17[0]},
      {stage2_18[0]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[1]}
   );
   gpc1_1 gpc113 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc114 (
      {stage2_0[1]},
      {stage3_0[1]}
   );
   gpc1_1 gpc115 (
      {stage2_1[5]},
      {stage3_1[1]}
   );
   gpc1_1 gpc116 (
      {stage2_6[1]},
      {stage3_6[1]}
   );
   gpc1_1 gpc117 (
      {stage2_8[3]},
      {stage3_8[1]}
   );
   gpc1_1 gpc118 (
      {stage2_14[3]},
      {stage3_14[1]}
   );
   gpc1_1 gpc119 (
      {stage2_17[1]},
      {stage3_17[1]}
   );
   gpc1_1 gpc120 (
      {stage2_18[1]},
      {stage3_18[1]}
   );
endmodule

module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor_CLA16_16 compressor_CLA16_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56036159923f7b1287bf6a8d50d67e9168f98753c5f36e0d71b9554b1e4ec1b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14f9ae9a5e71ad670aa309fcb7418cf5a3906a18b261af23de8738bb9131cc8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h783fa3160ef20ec3ba91af7aa32e8535c1b589405e78c07a2857489d5df62a6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc0df7d35a4fc20110a61193b6af9df312a989bd4d4eda3313bb6ed10f2632db4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31857f3dae9033b9923888c3094e4f6331a7bc43a863534cf9d24e0572ce03de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff3b059a7b4c7c7dda298ab9fe299cf224b64d7cd26d2c30d6c32a7735e77eb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9c7703a2f568f02b0b91ddd0030002d59594e855592d4f22aba7d9806a1af5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4636432146a208d66940def137b4a3cee28b06c2acc28bca1a4475cab514cc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc65ca8eb40eae56e695984b396e68214c8235cd46833abc2b58400427972e164;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82e6a96eac3dc67b1cb639606c10fe487550c0189ebb66dd8bf4f63b75311405;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b891bda00f15d00923c9342430548d433d6623d26bec405344c3e7a2a381c05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9679743e664827df33ce73b2fbc5b6fef1f1b41a9e1ca604441d04260f8f5263;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcba5e465aadbd627d733fdb11a728782831d180f2eea3f30be7edc2fae9c06c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41d6a15f92a6e9cbb84909ae3cf484d174240a82907faefe260d1f6ea783ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba51ff9068df97304edbec8b7f11eb350b99006d56a4d3c2f7deca3edc4a2036;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h805caba32cf8506bd916b145d6e45ac72d1d889b4da6cf4802af5eea82930048;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bec5602f00d7ec644db180aa97561476c213048854ca949ae80a619ef61a765;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3965b1835904c1988cac4640e435f854dc70c6e2af087b3c93de6f5b08f1fd39;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb02cf6ee4b700020397955daec2c2166dc0dfc72f7d9af92d768c3c76b158b7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a136b81045b1feb5a53cdac336db3a910161e0771eb8b58e6b9bcf9a7b48c6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9866fce58ed91926701f176cf5738c411c4f4e8c54613848d49ba33e68c65a91;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha7df60820b30669e7e7670723ca11a0c595249e83212ace18e08d51e151a476b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92606f626635fc4f7f41f5af34d8b76ef39b603572b22764d2f3e628d8a6c1b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea89f3612b1520ec82f81c7c09095ecc57f894348cd4ee8419b27ccd54cb7fe7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ad02fbfbbb53310e1f22c734833325f2cc77a158639498fe4e97a6d047ec557;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had17cbb3d38144ac0caead70d04c5a22b3c9427c80e3d8f6950ffd1cd86a6d39;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5dda41e458be06e271953c9051b37bb73105dfbbf3d4dfb066dd0e814c72a665;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ceba9c63e51f889ba8d5caf310b3b65aef39cb64a9ef438e3bdd3220552ce10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1051c1ac0b5a1a16edb391a1a81cfa28bdd0c42d32366717136707f55de9a6b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6c3fe25fef50b9dd24b006e3b16f83d04cb5305957fe79d4f3f5c2c71bd9aa0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb1ba26a19dd791ee3eb61c70034ae0748105f7ed2d94aa812b8fa7ac80d1d66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7ee05d1922dae922a5238f814340b52baa1f017e70c0dba205b5a1a909c173c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8ff5c99b10471779f193977a86eb236112aede8e8e7626c5f4484cd1b2f64f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf7f06a7d756e82e4c4207b552836c3dd3529415acdbddf929ea546d300246d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff08f93bb4bd2f18be32fbd4bc4646be4bcc0faa690f8ae840f4c0b4b5e16026;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c38c439488bc91dd395e11deda3fc552253e99284212085d6f4c3f765b87c82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbdd23e0108eb6fd5f80ad8d8ee7f0725c3d000fd0c7ce59f5c27693a36900201;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec9d506ad33baeacd1aec82281541ff71418125ac47cdebf1a00873a2393c117;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b2c3f1ec334a35ce077c739477956799c060d3d2eb11b29ecb41fe3cfc753c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef3f83af4113306652719058d636a0e530f76e95c10ab6a0cbaf828c5a09c9ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ea6b29a2cc0c61d7a39caab259a3f167c9e8a5d8fde853122fb8202929843a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97e3e202f4c1ba98208558b54c70e60b82ec99e14cf695b71f17cfbc5cf5b0bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5dcfb4d80ce18064717e10d5b367c70fb3e41108c39422542d7118a38a286915;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf3d02c98f4ccd0bf166a3ce23a3a178cca0b6939812178df9186f10eee2e8964;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31aa1900573248737ec0782f7b3811fb19d8e9c3f93952b5f424d9bb24f1653e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9d16a603024519a4e903bdc986ac91557edc8f4f1ba44432027bb7fe9dbf128;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba66ee377eaf886aa0b2e2b6ebbbe453c064edcad86609301cb931bc56dc8d6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96370db80fc4860c26880d8367a50ff5fa8932bb8cae88503445f8e4633869e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h327da47eafbcfbf07e9339066c1eb3835e66bde8405dabc5ac12d1f940c79884;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9f6be8a2ca4ddec57b8b8280e792eea6620ee733c50f1272f69abfff00148eb6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73f2e6c2bf7f65d61f5f2528a601b01bda47bdfba3639162ce00ee6515fee656;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he64f8282f1a11e986026f76b6ffce17857219b33b6bc1ca465ec499ce5b5311;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11dec3bdffa820ef506df65fae1d66d301913c172ec189ba288e7f962fbe634;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h51af50898f565e76f38c8cfb052d85ff0f7ddc8ced5d97197f6ce5292a870c01;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1341228a433a872f0cb28574f03c164fca0f0395c61dcb4c581c0e5a1181affd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h331adb63afbf77a06c92eff9f9a7deffff262a15baff358e356dff7d29050c24;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5eebb1fe8c937b8317765b1925579174935d68273feaf69e1107c785fb07a556;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e4bdb3de20c1f5d95fbb7dd2fe0b18aef12d88e2db0108108990ae6f4a35360;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8e6059e9b056ccce2510dfd76fc63644ab37aacf27f8dc9805512cb638a0d72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7b2eefd12beee64d044703a47342b9fbc2047d42f9de22820fc8f93cfaa6c18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h484825e1d8d300d9dce59327dcf4790559dfda4bd72438440afa8ef092f44568;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h134b418a7a70dae328081c85d00e80f3c755a2095746f3612ef28cfd6c61a431;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6385daed90ad998d571d19bc8e157542166d0c2fcf4d1754bf76c7d3ba3394e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b35353136b787cd0cc086f07aed8c92df2937592dae1030ba48a89cdab0ec6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d1d58f701ca0b01cfd1dcc21f21811e04901b8f515db2dd6b9d06622d076c17;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14a3e4006468871be0ecaac3237548e71166e68d060d16d4c1ab5305352628c3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1be773ec8bdf73f31f4e5f2e38e9eb497cd3ed60e923bf2dc7c3569c6c3bbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha078fc054bede275578f2b0df3ba2ba5bf1dd8c6cc9a3f55b57db8d0fc6386bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae9e3c373c76496ede2798560dedb2ff7428687d2032a26a7136e1399339194b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha429f7b9e79bbbf01cfddb751fd9349ab57222b613ee8d218fab3727fb20f53f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf457d8a7c157445d397fcf26cc02797c30c0e3c9986e7d931a166649d44edd9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32f986d8f5c4fd78f6007571eae063d8845e07fba498199700540d67da964fde;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefc47c2d2ead8336ca82e63ce4bdd1f7a7b25c636c2edd470f16312057f55cef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h26463a18fe7ed3defec4faa3414f070654df24a8b4e7fd34759512a3876d627;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12e13ebf26ec4efe1c47c068c9d21b2eec0101e1bf0d831e97cb4519464b201f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a486bce39a72dbd1956e93354d5ef7b37713bb22d39da8e03699200c32a9ce7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h95597064a9e5c51e8012d792a07f0f29f96707f4c10b11d43e326036cc31051f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h562f63e8c8bf30d7df9ed73821c2b5783f22e2912d57a7281388b0453230438f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43890841e0f4b6e6c05a7cfdc3f62530bfc2535d00f7d8d1150d2d8b624c3149;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24a359f34e76501cfa722d67c77c7da58dc09a790aba0b053bb138fdcef4b45f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6656b3faaf16111e458d8ad6b11c9b73d6e82517a2a80bb4392dedcf6f1bbe37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90359e882c40526785aea3ed3add346f8656abf5b68607abf6313876b4b1f507;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e196c6024306edfe89180aec01ed278a464591922988692b09890809c8d549;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2bd4c2c7879fb431bd7d17a60d7415340b2e51c2a71643e9d2297c42e0d7e7c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9255e9f7e6517bfdc4c9848b7e7c16f4f63fa976239f04046cd791d5ea09897c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h227f7793c55268e2c68104d0579be3c88662bec5240a747404f24e0970e8cfd5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8ef15d19a281379f8fae0b2ffcf5b85257781491e2c07d70dfeeb08d734b94b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49d2bba0d9c1b8e76e30f784eb72c9045736a4e96a161b51f5bbf88a11a848d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67dd0647240931f757c66b8be7db6d073a62de2d31d80766ba30a19272f09750;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68be173c512cfd6ff89937946708b2b0ea772d4897a3104c945d6bf253e8f0c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc2cda15d349476135881e12e4806626a312d19e7dca7512441840c5ae1ef72e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ef4ced0c7888f00ff3503d73d088d5cc37ba12acf726105e938f2c866cbf09f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbaa4b6640fad5fc9a4d2cf07ffb64cc97ea2b86265105ccbb1322b85287d6eb5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37b81d0928e225e6288538ac65320607046abd621e28504932f47728bf0967d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3f30ef94e60b53b89e3bde906682bc58e64565eb8967d5ae0a2a46598297111;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4870de85759f7a3a5c2adaacfe6b24689a3cfc656343f8e6142d7bd038a55582;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc18c5b8c5ac18c4a1dcb434b32578ec94b7ae54af6f9ca7891938369822dd800;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4b3ee5dd2ee72db4d86e7cbb6d218d41e920eb1c47b4a65a85d7921ca1e141c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d0c1d9132b00da71cd88c95abf9001ee1c2bd70d0c28229e197a8594a2761a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefcdac26130427f05f19ef9676d77b7ee8cd0acba7f82e02ef549ab2fa324b50;
        #1
        $finish();
    end
endmodule
