module testbench();
    reg [30:0] src0;
    reg [30:0] src1;
    reg [30:0] src2;
    reg [30:0] src3;
    reg [30:0] src4;
    reg [30:0] src5;
    reg [30:0] src6;
    reg [30:0] src7;
    reg [30:0] src8;
    reg [30:0] src9;
    reg [30:0] src10;
    reg [30:0] src11;
    reg [30:0] src12;
    reg [30:0] src13;
    reg [30:0] src14;
    reg [30:0] src15;
    reg [30:0] src16;
    reg [30:0] src17;
    reg [30:0] src18;
    reg [30:0] src19;
    reg [30:0] src20;
    reg [30:0] src21;
    reg [30:0] src22;
    reg [30:0] src23;
    reg [30:0] src24;
    reg [30:0] src25;
    reg [30:0] src26;
    reg [30:0] src27;
    reg [30:0] src28;
    reg [30:0] src29;
    reg [30:0] src30;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e9b6151cef05f141481b79013d626eeeea3c1e213e454b2b5541d9d685148134671ff0aff6aa7354eba1d47f4aed8e0a21a5b0d535fcdb1dcbd6d96ba7100072951a8c8d233d7dfbf7d55a4b9f4c06b3275d1f2c4b65dbd2a3dea165bcb3d68dadb0836f8f0a41fe36907d6c3ba657c14c810382baf4f95;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178ab93211c79edfd22950b8c39e646b10754126565e17005bbb094fda66109d1292f416a7eadaf566d07e9f02de1fed3ddaa57db0033a98a8e2c242bdc5fe27e2396fde9bda70501ea6aa659f4331903c421b525bb496dc302f4222de45032addf2924f0f39ecd70184ba96cd5e7d6ba48ebad559af7c3f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac38910c217a3f53403103cb2c60a487f56feb71ec9e3c9c69ab996127fed44d292067512a0d31c42d8a55d243a0fa2225fbf6088b49114df932496b0fd9021489f22679995c39430bfed2f244568bf1aee24069f9df3ffe0712f7960001b023f60074dc87ad474264641f53236c9b949a878c0903c62657;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c683844f866847abfd678b692df530d6706cd080521de3e2ab7f5052435a8362f8aea83c8faca5090c09d3098c81b4eee31eba7b6fa9c48f0460d286505b085d33dcb2fd8f0ace82c3817d312474a9fb6c4e4408a242dbc0ead8bca936de2e322295b244072b7d4fdf98cd76e89099b1895cbfce8bb9dd6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14fef0800ee735fa9e48940e636638170bcd80c90db3aac9692f4db7f00812fa2c0ad7fadaa8983a4e8798ca1ff9d30c67af7fc1d7a1534f15348f180c98bd25c630fb21718b6d1f902f419450462052338d9e8c70bbe4b3f70960ed962cebbc1cf111e3208636217c3550921f8a23cf8183147df4d9591e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4650addee63489066338207815d021b42f7eb370c457e0b20b64bf916aea896b90e7ad8cc34131437c0debd9654ae9c14023691ea5473cfcf959c4e246a2e3f18d8ee2c45bbbb4801a97849e5b2e5f074181276cd3ceb1ef88d21250d8d4f34359507bf8d377f8bc60eff0dbcf0f1a8033143de21a90b9c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7c2c3caf7ca6086c8af98adc0f341bfa978142dc44b2b8bc78df2e48cd8f50a3830ff91fda3f9cfbf448e16cf404901eb9696a137849e5c758904c5f477bf7d5633661046d8d3c9ba8b5acc61450884ec6212ffcb68053f95345c832d5714bfd51f5d689733802d3d542eb10bbc7e6fb1c5d3758a9cc11e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa8bf6bf8507af2d95ee031157dd6fe4e39759716e86321adf51eec2e1dc9a05675ced1484ca3a1d5579c27d5e64ab9b0ea73508c12ea085678a21b97a259a749829a0fc5d059b0ee91b2b10332f38c728a42978b55f57e84c4b00f10e3432d4c8d6b87fec12d86b6b784e31b78ad7c0e8eaad4aa28ce03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba593c5462c618f55c89cfdaabd8825161898b5a560f1b7c1ea2ff6533a2008054588172922e6b672ae8d44cfcf8903f3e0d1b10660baaaf873d79510e4e5c1d437c69cb739631446c76d8017e5e86e8d4a7c9e0f1fdc1e98d61560a75e6bcc14204034d9e66318a8a24b556ecbcc24c86475fd9c4c0a398;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c7314b5a036d664130c2b3d8ce39e9de676a597e5d36aa60061e42134890058e690e6657192ce31d6f23b750517a20f9181d378b4a984e6f44d3e136c4737f4bcbea98ac7e1a1ab15734dd835c6d7c59e9b79bee6666db12387be03cde68672b29992198e87050a8260beccbb7629e95d2d5e76afeac4e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ca2d531760215054ac8382eab30aeb3b91f276ab20f589f3cf5b0da545ad5a3b9ab434998974acc579a6689573aa5967464057139a96d8f1955c15f6af580afa3eafca404a63bfdb224408de71cb540d3d8c61372685153dadf5614f8fc661fc5a9da652d19069cb6f5493b175a2e8d1a64ac5c0a017549;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha87bbe14107446206c2cafaa6b1ea11ec3e0a19cf69fb845e7451ffa03b008eee60c6fc85db87ebe6f3687191e974415c66adbd9f2e2d71c707d2410b354dd802bd1599b01723ee2dd38da025396035000421b4b7f16c1b8f8baf6f05585e474999b31aeee88a6389d2c820642678762a1958c87ec315765;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he856e0d893cc0fb67dc7cc4feb4eaca7891201b0c4a753458cf1b0b3b7a16eec36d64fbe15e2dd6e87e1f9e3d321fdf1a2f445db2335227aeb88c261ab7c0addb2dcacbd42dcf21f7c75cf46ab405cb443dfdba3efd3e4700b8fe0ab16eda9cd654b49b3c4b63e4f7ce734f445f87d8405606bdffbfd047f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6407ea9ae9556c0259ff2f287471df16ff260c51375f7441e8158fab715560068662b50aee56c912d0c24d8dbf96ec1c1607fb89f3bd6b69b499ce4b4f789f309bcfa4c843a3a32b1cca06ed5b4f279fd388be82d0992291a197f5e8bc6f4438c42cfcbbfbb5c50258853f46131ee780d568b0e80bbca7e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb820b83e09a4762e4a1e377c5e6408847653fc46008d8031a4f888ff2af27674afd2f3ab15829c921724071a392286ec7a55778434c9d4173bbb69ac3d9eaaf3a612ae467f2088fda052ccc47db5098750803f9151be875d6dcdfa280c6679606fe80b57960cd0fa0487f267dd00159849a1cb57d9b0ff7d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee822fbfe0f42a223821083215de9ee29825dd303207e68483981142c4191986617e45a2a1f3a91f15e900d5ec0d2d133956d063febde1e287ab357e01c849769987f38358cea5c979f31bb46a3a4c0e579f39781e65d6b0dac4b881a9f78cb70d61239051bd97d1315642420557c30e026ce57458ba926c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h24de3315f80dc47a76b5b916a5a634502b987dadf0aaacede06424637baf52682fb9f98098f1ab0df143214ad9bd6d09d59c7a59689b84a0863700fd1b627b3771e3046192dc6e4170fd3fff7836291c3b9731614e0c76d78652d4b2e8161b90b5c57f3206ffe0221d12a4aa569ef64af3a91b01b9c6112;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3bce812ac8619043af55312d103bf1a4215fd1998380a167b213f67d4aa6cdfa7d2320e50e4532bac9a4e0dae4a50ce138d39eb35dcff82fe7005674c7dca73098c89899a9bda37ec6af69f2fa6a4bb6221149f05ccfb86520f72e13a38343de2d88ac84b704ec47c5cddcbd83ba1f3525cf0f8d122ef588;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aba3180a9c42473792a9b4449a6984c993025e8025cfef15831f159655377503dcebbe72957c6b04a317f88b8b7d70f35cafcf9d361c099992a1fad6370a27311f41ef466960ddf7ecc900d962545537f6ba9672174b6b9e1444d9f6a46479bc3985d22b89f7af67d805720b78ba14a62ecce593d9b1da14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h140e122c90cd66c2d6f1dcc42b5dc37c93a22cf79be5aab1f87bb9e27a8c50f826a22742b46f7ebd64a1fd04977ffcb5662e08e1dddf054a4be169bf08b0c7e0d08236b3c608125f891485cbbad9c8cfc16ce650a190faf94ee9b9897d1696f9211b7dbcbbcf9887d0cda59657c10dfc871210de3ef4d9475;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4f834ca068ca170af0221aef479470af1677a9a2f30c1f2c82a6f99d098412e69f8b21bb35df951472ab5284554f0faea196523007c7020252168ff1781d1ab93cc018404e560a20b18fbb5ec5c3c3011cb09fc2a1a6322f766d09b1e29140ad3379392349fe7215d61163c6d7f1655962d5ae94a4ad3044;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ec0e39fce00f7de1245c73a6ace96b0bd3df8026d61087ccd2504227b2c9567f23c25e55b220b762e9cef845abbb512fcb0e603fe06e0e78da906ca625e3e3fb44927981efbd45253cb021a2fa9d9cd1f32c472e6455b4c42740b18aba065f681e51a57be51c468bc0eba86a550672bfba6fbc0bdaf335f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfbedf0c48f64bf90b6b355af0849a79a2cc5103d5c752566671a481a915c4f558ea3875aa450cc4b874fb701adca08e21eccb251a19d84f6a1135e3a8a835a3a078e1ec1a4e4dc2f723262992697f6e81b6f8f9dd516268c7d5796dfe036641d8377209b45bc2388c944ebd83836c69b5c39585cb13f18bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h87a9525df21096172bd0a7ca5cd46fb8bf4dde52caf6c41d9bb23724be01198595650cd5a84bf3317613d45a463b8ad41ddd1abb80f353206babeb678c52779bff725fe673a0107c470ccc26de35050d0ff6082d20633973d9862fbedd5695b45d21091c4a8d6271ceac87421b9f86e3932687da7ba50b48;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b810a4b283b9cd960afafa51feeb830e8a4359fa6d3cdeb50b3bc52066cbd5e38b12d56b814f30f8ed741f24cb115ee28cbdb3fdccdb7e10d5c388b6fcf6406c66b330a3edaa91a4ae8aee4ad2b96dd6e4227d4f0249d7d8d73ab4a3d6de30c615baf881c52e16263921717dda6a4e827c45ea72916e5a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe727fa73b5896cd00c81cea0538ddd20f5a9d928fb346fcdb6ce2c04f42fbea26a1e202fbff9b8e21c444addcdb65370765d28ef4588a2a5e6c32493f1029bb49b50d920e58e399acbf50290c01a51a248b2d46d3e6141ed67b4925066150fa72a706b30ecd1004f0ec25c9ed060a1fc8f75890795d8df3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3ccc1e1bf831c3f4602004e323f198d6dd8b55b0fb739abe91ff7b761766557305bec4fb01b34cb2dd61faf319160b0c8f6815c824d6faf0e3894fb939ad452a91d824145e61904ab070f49726273f672445f533ffdcb182d7ae6697caa8a5a4cb8638ca0251d5c0c45d760e924f32e1c6dd3fac89d399e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd3e2eb61b4003f06c4c02a35f0bb281b46a6a3befd2922c0429a9904107069e94693af75fec5d71bf8439ed4576cb63cb90ed73494395be7e12df3e71709dbed9d5266ad5ba6d951983dff9a04c612e31f38085c4ef5210a3ee365c0796aab17741205c7cc061088f2095b009289dcd324de823fec828c47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb44a550e5e9899ff6a5e7e6ff6c5fdb958b8d434a84491ae4c2c592a4b571dca84cb0ca90e5260742c60cc3a33c0a07d41add8e23849037264988090ccf4a8901dd1cab68b465a5d8a0b54f4905e1866c2c3cb94f3d992cbdb348f03ef2f036d0be774804858995357c2f6febd845903c3c0c22d452c0d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd541d8bc4c6c0df6cdc3ddf1d11e76b0582b1dbf292f101e9ce8341e997ff68f69fb6c5776b6b1822c9132e36551fac64c692768a0ca88ef89ac5aabe05fb9c24ad7e7a7948b40e6125e81d674da72b3f6e3104ed125b017909ebd1ed157e1f9b12e94099965b0e08b36fdc7122a3b54c622df07853f95eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h21034d6df7e86674948fe3ae88bd6767df675dd283de6a7ca03daf52d0dc02286505b58b2e56d99c807b2803234d1d928c1f958f9312950bc964d5c49800c0bc0bd6fe6f5d43cfcf2de02656fefbff6a71680d00caebe444c89e83f5ba509ddfd8d806703684dc9c49c61742a87bcc4d95174be3431f1573;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167c0f01496b13bdcf228434f2a4cc8a821d082bf0cbba04c9dd32b1479ed645dcb5887ec46eb752631f86e20e91c02977156642ef9ebed2314c8acb95e13bb04dbfe03c2049c9714bee378f773348198c398e0497ffa46345c0ca664f3f4eb58bd2dbf514f5e61d598435080c4892487efce22be067ba69c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h131a24c63fe77a5b13a664e72d14c72e020fd8fc832aa6624082bcb612a0296054446fbb402120995d3d8f4f8ecf826393d6a30ae0fe69ea51d49092678f6e343596837b5a2a4fef0d16e42c0f668d944adfb85eafd4ab624ff5172cd83f541137e320bd7bdd17405f781932c6fd3b6193c7e079f85b9c83b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h337ce3407d037990eae8bdc63487c1f3028e97ef57d7b1d6981a1bf9f083856c4430a1da1c37964a493299ee9b71e89c20df256fd410ac99feed44363c7216e10d30197ccbb8b9659c7530bde6eb5ba7904e15c01caf01508753f815705eb5e5ce63e7c3a479ab5c8ff982a547ff1ca003724ffa86354c63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h183adabe884380e1a70078d8e867509e7eb583717c94d88363f9afd9b58f08c11ac07db8818ec4bcfc4bc1b985279367f9d3126b88ecd644730be5e2fbdfba38debd66b19e57e93a21201b3aba0d9ed9e10ad22b495d891dd3fcdd305b720632f80e74e4fd903a51acc4d8c7cc695f526c6ecdabac833a4a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e461ca9276076c2989357434133bd754e51bb2ba51c02c61a3901589fe97f86695751d38f376adf5252f127d1ed5f228fce709b9dd931758a2c689bc19faaf55e035cf18cd1ca454c2070145641d1af765e77cd27e4f450d621aa808bcf1ee1f21e5e4e97ad02955d77ea454b96a9a0239bad09b7c20b13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82b3ad70a29172866ac3ac8e88147cc399058ae431cdf5a917aafc83f718c580af228c0175667a79b0d39a99c5c69742d4b0501c9d20ee799f434330aea274bac5b8403f90dbd1c0322afaca8aa9100e2164ab201f4e25cd28fae6112eb6b3d721b9cd2a2ea06bab264691587e45736075e970b9abdd5896;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b68e28133173a2193fd9eb706624f02c7de408e6200910bfc55851b3e543569da73228b965f6750f7301f4b18690618fc479a75f5f8984e35bd7694302560fd70c9df2e5bf59321cb929b933f9ba128f5996bf801406a4e0b5c6ef3ae10c91c57566b67145166551f218b2e02c0f147301d1bbf5aa0d09f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149a9d286857fb13ddd9aecb6fbc2e9a0d5b2367cc168b4f2c77385143eea421672988246c834cc7b6dd0e97056ed75a9e7191bb1917c8adb8226a5153062a710069d7771953ba32317f7962131f6d30e2e8e6f6bf7a0212722e383c6d4f9d0e5830a2b5e5f352c2cad1de11b623bccb38f1d47c5105f09c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3b12e112c49a6175c46752999d3843f205ab8ea4cd0403cacef3368bb822e663a192326f0aaa62bb4834ff1d15a19b05893ebb89f19f5dd780f2d3a39439c4566a11b373c8f0df0dfd013fd95a4f8fd1ac64acf6ef302b32534dcde9def66bf9c08cbc8f48d5c2a3ddd1d63f6a4de152477e4225e9179a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h87ee96a958e89e6f3d9b51d2d17492cd4f65141e639edd85bc3e9b1fae8ac7c3bdff7aabed56b89faedf49fe3e4a77b6cca6d3934a2b9f10d04fa37346fd48311fb5e359359a18289e1c4e77a4c22160ff7d9107a5d825701e7072fbed5cbdbbbf22efef3f0cd1cdfbbc8c6f71c26387044154ec633d4732;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c1d3257e27dfbc9aa2be68515c384e624ebd28759619fe49c446919f69266fa9bd466fd29a2317c79acd94b5a93c5f72e10d586071f31463f6d8a4a705f36ff130bc62cd15f90851a083596df9e2e9f005eefca71d518d46c97414ac130e927a88f0da2f11de708c9dbd9232c13612e7591401d6425b432;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec593c44dbc7e054a8ecaba5dada6d74e341e7bda9b4256732a571192b25278b766f33035a4fef0a0866d78cac3c878dea6692dff5df197e27e3ddadc3609139e2de0f54bc3782858cf2df337959ac8731f3d2ebb39d5b53dae3b85603c9625b1d0cdbf9b88023420911f92dcea1a8a5b3612455dc75506;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1af9ab37fffe60caf5b10e2b9b2dc3d586c52163f3a452b0d7d2a9b36e59898e667a4ca13a55796b6c521843ef47bab2285f477259a163c1748c35832f3d0083e51c5e11e50374cf9410b5c85c40c797bdc9d6ba55439fe5099ebb5c218b60777598f0c4e4ec5cdd92d4c49076b9ea457cd001033cfd0e2b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d210e813375c5289a0302534562b7afdf18eab87c8d8d69c8769cd9461c98045e82d394be7ff44b64c62a2b3798f5c15c091cd37a3113b68186d7ac5a172e1a372b72d13d47fc1bcf8d042e5816079e165b07f7293b63f1ae23a735cf13c91d75cb9dc42d07629583e72aec75a665a19d041eac1767941b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138d78f1a9da6c798ddcd9d1920e3b2fd3ad98c33131fd49a4051b6c848c06fefe69d04ef59438da1dcc6ad0d04568a2560deb8b5249056008b86ee5cc6487b2e4fd1c7b02f6b553554ab55b15489ddc04bc74aaf8b1b9c7231056bf05e1be4977d97ee117281efee8f9719451207c7a527b7dcf5d660570;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1260cb5f39d2d38d46ead9d4b45f6b4298a363b478dbce65a1dff50eab90cd0c325aa62553a120d36b683434f20b296dee66d07a14edae25be337aa09edc54fb1f9b674cc2dc08f6315aa66774032493256b216b5e07bc3408de1e0cdb9912eb168fc1f95bc01dff8b6ccbf1d112e95648bd41658b79a5f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127cbe4d1d68adf94ede55549f467b03d84774d938c25b0e8fe08ee592d1f872c0a7f1b1116242c2605b0bd9022424890a4b9d6a3a2844c70351eebe59d1c5434ae685bc1c5f5e7d8cbe8ed25a91814769256c96660203bdf783bb6ec122f80b632b9172a87baca394c75e69d5d6d368aef82d7e18c8886c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee695868f710ef04fa21b99c7f57d9c0ae4194a5ca34a98c7b848e6437ce4584e5e02077f3112a47e2d2afe7d106eb6b81de38b57f706f419a688b598afbd5ad205aaca5aca0ce1e43f703014665ffcbf6e5962ce353a0285d912fcceb41ce0ee24804e5cd6e88500aee90394c05c41320935b793aedfb1c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf04da3abfc5925ef9ad5fee9a10c1da10cf69613c4940fdbbd9e61f3f0151c1933072c1d7585dffae618af2e022a3304ab08b95f5af9c100878ad978e69f6a00b6dcefe5edeb852c628c289faf1374131bd113d5ea8effd9ac1051f2a3edb9568f319c4348cb289e0433a2ddb912b1f46d52791d1099083;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ddae0a611d4045a19e65aa677ef7ebc375eee7556a2afc455cff5659b890a013655a054b59eac2e51289838c137e26a8443f7075ce212aeb657edaff713b91c4c787961bd76f904854e0f04a6e42dd363d3294e7942512f0a59e4aadb34169057d1a65a8f3835719e7167ffbddda602555690e97d4ade9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b271e397a3b3587d5589424c22d3ce0a899c83c1beeaa226a27425771a219be1069311afb4cd8f6e431c2072300b872204caf143fbac9e69d52464ba29383305a5b1cb8c95aec3c6338067a478b7b7029371ac666046b5267a1fa3d12784aea36e583076efc9437e92169be2fdf9d0fa58d5f72c671f0a20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16675d09822834262142bc0544ea356132fc84ab8d74d66e31834d9e099e4af424770360189890b11468fcf7cb9dce0326f865c8e041feebb9501727fd76f4faecd80b392f175590346ec51860b36b814a49ffae2e68455695c88217925fb3da2e725162cc7c39d264fa0caf74a0c25b013515b42433c68a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b954ab0c1cf0057a013d0a38b75c45d8c3c3a08abca8dc1c56cd55a86c42a77f86dc7eee9eb453fc7883313af35cc0b9eedaeb119422b4b8a6091c69ed7baf6f0c04fb770263b1471729cb270bb25b04e566d437612b623e4b5f155bec8223c4e57898edd883d88dca49c2bcc9af646067e698c2b80a197;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb429856d4e1a3ecd68b5831d8fad69a0e4e032eed193bcffa91770918d855e992569508dbcd84a8792fbdc99ee762f981d143dd2f363dc0680efb9af935e50038bae475ac48dd260a36e5286f8a29dd210c693a1de2e11e4662a9f0a0575b1e24a46242cf6c7059c5c2d03f33b5aa03a2bcec0772ff77852;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha56e72579282116b65c2426dc785c72ffc24126a89cf64ad0a757553999bd1a8b189d99b7e2a0425d49f9374fc50f31015fb7a677dad7323378e6422efc0a8fa99b84914216c62ff75827f9a45270a9099e0bacc112cd35f4ba09534632412f4ace7f449c60cc5a091aecc3bbe614ff013471409afb39215;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151dd109524c1e451a9238a520c723bb73853045c0d482d85c674148dda3209e1642de73b629e7aadddb1a8dcc289e36ae2a50bac1d523776dc4ac5f6a2ee62a9d57a849e3be180309ed09e0099ffc6aa49078218f4d7ff1ecf5adba0dc7a4b25bbdfddddab6ed28dac5f09f929fd9f1d915bdf536e2abd8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb188fa5ce7a96d6a5ff31c5cd122272911d69ecc48c946e3e26f45020e94c599a5c5330b0637e491c285ff4dfc212cf61e040306ab01bcfc3239d880623314dbfb942bd716ff30284030d38864f66153319dcc0072fbd2bf7f338c58a861b21e5552c528824fe9927dbb93244727561e226364a93e8e6b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2886d429c2c7c69d3f43cb70729d004dc86524cdf750960fd29f980b9e4a99adcf469d597bcc9dd57672f33874102cefbef5da697a77b43945aa2965d724c1ec097acf18735dbd5b13fd8790f7614329dec93e2c53c822ced648dcf5061aeafa366edbff7702ffb1b7178cfe8bc3e8ca18ff5b89b43559f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfdf9d8a1bc5aa9631d0027b84796131024be5e454dfe494d712098747c06dc401ba4d7d0ce3696d67b3ace50380fd1847d62d61a138ba51d6d06fe6439a2ecceb010c0f278ff76eac20fabb7f9e6f748f2751e89f2982496dce31ceca9cd2bb2d5eb13822ade2ebf94b7bc50e0b80ee4dfceaf7fd7c0fb30;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1098dc5e74b59c65f66c4b5dc3b94a3fc8a24f22ab26ba72af7b6b13e75c1be79c2789ff08a403f7a9cf7920276c2cb9b7e00ee2d4dfcc5ad52aa952983bc2bc772405da445bbc8172b8d155e28826bfea58fa411fd503eb87c4c6d1f65228514087f19dcda50a13cc954d4cd35254756381dc9e9620bd3f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd43b5d82fb501eca948eacbdfd72f82852a4cb9c51cefaf553e39fec59c769cf36b2378fc7e66e58c1f9094250c2b71d7b6ef5628d6b355e6aa9bfcc504051d8820e758489107fb82504f78b0acce528a1e518d4f9f9878fbd04c5185337294369f41f2e731e98254f135c758030816b5d3babeccadbed46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h846b7fb25f263889ff077690d338c7bda18028f87af53b031316f3c8447700419a27a09a403050dcb807a075862353a0f6258368eb66088db64f268d9d0b30e0024bf01a5784c69ae0b7ba2b3c73d4531fe24fe5351edb91b1d39fcc5cf7231057c0051fad873846804dc7811a06f5e2976169612d8f05f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1513558cbce567e58d2e733b736054bf81f2e2676681cd50bb049082f449bdc4748434c8481043c0bb873fda674d29e5e17f40fcacc090538853e40eb2e620dee66219699c67932b943f1ab40ce4b98186c0a7645c9da3daf2223db69738686436d2a2e80db340532440aafcfb89f7b7877ccf347d7e50e90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156c74748c937da7bc1a443a712e10a98cdda48af678af4967d03b29a90aec26121eb00284fb2ccc8525a3d9994a0a8abdb893a8d6c4a4caabe9cae5c439b25a99b407e87266f4daa809441cb9054e6d4d934add5abd73d5e70b5345cdcafff0714489c3480e488878eddbee345b0318407e91e2724012299;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h87a02327b5e0aa74b6ad5cede9679aeb9e59253daf3e2ff31e14f8741b93551c8b63a638804edac08b9636fff3993efc7bd7a8b7da9f861cf084b3a318182bd6eff3a7e80076dafbb0a12add3a0fabee4c32f4bbba07a950f37689f7974abe953de8a2bd8bc1ec4b20449a3ebb89cfc2ef587b8178fdc9d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha74d4e837b01c5edb64ac5b1c586a7395553af0e75e1e8ca0253a96b09a6a2b0a873b65f47180af6fc092f3b8aeb3265195d62c3f84315f0bbfd943dd5ef89497ae597805d2d644482668d1665a3048bbffb90cc329aabf361061b914e9c8e16fbd55cd7a2679602c9659dfd51a7730bbdf1487179511c63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12c59809e5b10aa2f4d62992e508a3d11352ac06678bb7c1ad7d530a86a4b96d45f3d1fc69656e78764be55ab2064c37da1ea2055468e2691c14280693209fec9829c18310bbb0eb896637e18d534912bc5f5f0a619d9b5ba9a16170e56958df1ba4466ef78acc17b40a3886c85c413a5db18ca695ff0f78a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1458a00fd27a85e5e888b521d8752bc4e9f9631697c330189aaa15566468939a0aad07053367a71c46361ad7fb421cf00cece974133e4499c5b5f5130d86ea01ca9ce7c734f0b258154fb7970bad76ca16aca9f6321cbafd01abae370d1c536b9309ba7e3158bfa8d83dfc471f328008875f16f5278c8b8fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h414510de77328af23c1cbbee38363d77f906d73508a709a8c4649c889db05e52827a6ac69ed3af5220c42a5ec6a3f60ba2d7bc165d6fa4fc9295ab4f11292e62c3b192a0ad21e34d13d38d76d8af887bfc385932df4f01761a778700977afee707e848a2164337c25e3ea8f995efc21da782a32c9b4264a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf119275b5bf4d66063e19560b9a81e7f043c003938c6e0ddcb8f780642798bf332371f4a47fd495f41a8f6e466d51e545c5683dc06bb8a114001bb6117da501655bf11d1a72e1a14a5a5457fc988aa7036e12f798253c91835fcc03b65d981520adbad7a893fe20c6daa4eb316c1a604ba05c78884b6fe74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc871527dd42c48dc4a5207b9b75414febd5f63ca2fb20e70cdea118de5f801074fa936612d44c5cda2da150c3cc125647e0dac1f447dcfe3d119caa20f1cf19e5fcfbe3a07eb981e5a06b53fc2fe03d572233863c5ebf71a5341430a0d2bc4fe218a2b41f267bc4895156856951391ac53ef4ad518721fed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dad0660a48e3aa6907cb28447b3b66e2fc7e4b8f73603f06bde4e4cb4f7c870f942005c2427780da7ff553196a6c67cc7699a1b70fdad0599684ccf5039b8a6522694d4f5d6c64ccd9c51f8faca9feff29821a880dd2b79990c3347797513f0facf17fae0348713fb8bd428f707074d596e34c1457509bcf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1595820e306b8e830af2dadf2c6ec99e5887e0020d399b7e7a03ebbcbf8daeffae720407acc658b39378fee67a5eb93400f17d3f7267a682eae801830bfdeac74ae4661935967e57e06033c07468569d42b213f6c48c678a17209af7f7cce0c9dd579ea9fbf2bcee3250f7d974eba13adf75c8fd9bad5098;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2fc2bb9b74089484211673342ece6690fd154dfd3d5712e7836e82c683b5d6b2b9203650272f13e7277088ebcc55b3c99a7bed83e4023f57a15767f8ff1f1c8307974a317179d619246eca53833801667ac2a58ce2c547d7d60e754b42363e69bac474bead9daeb5a4f4ea75db9b671dfd9487f64f37c96;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118a9871538794051667e2920c27f1158ae7532cd70680c047f40a2d4672d8fb14a41937f438bafb7e9a805b12e9d2208d92b1ceaaf7c7f545f484cb0b3adcaeb6f9ebffb0fdc8dd93752cac2ca0b08733122c7ff8ad74d7d38cf8521fc31826de532974207f0fd48b403c64b90707dc997f5c62a27fdcfd5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he521b4f8e203b95889a704117cf661e6f9b2134719f211cbee41cab22deab3adc4643e3e409e00af276c75544c55c36e7672a070825fe5f90c230942b52f34073f91aede58913ae9b7fc5ef1c3372cecbc9dc2a52fb4a69676c34833785e1d2f2fd362c37ffe306ff5625265f8e34eade04518aae42bb1a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5b5dce7c1a2eb39af0a6701cdc022037138ea4d3f6ccf02cf6c5b332dd09de34087028b137125cf688ae7aa6f0b1dadd1ab55a855860a910eb3e0bb87d561a75b5012e9e2fa5851783acb82af0787ecdd7e294c290fd5a09279d1199e833d713bdceada5fb2bcc63aff439a49492d5423d09514c0be7b2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h148a47dfd3e9640625878257d9b3e6b9d359e7d19b468d3cbb41c06ef599ff8353d24eb479236429c058771fba78c43f77735dfaab0b5fd28243dc94af9679f96a104487894b9edb740097d03c4fa2ac11cde10a0d0384cbc8d70fdab5a9179c897b7703ff93517b31342b671851b240bf068983a2fb9e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf10db0e8c160bd4ccb5a482edcbe1e6e6ef51f400d82872e28029b49610b3ad6ace570a6caf8bd91227e3a7463c5138845abbf2927da17b7dcbff68eaa444ce9d6601d2d375abd97d56f7745f37b53b647d3650282a8a4261dd7173caa98a1e8d9259716366fb113180f22c2239c56674cdfc5a2c89086b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8dc486664b1888d811d512b300c2462cb4657fbed96726e042719ea7a6e7732f0326e06665228ac57e90fce4d1d58d7cfb40791e3f48261976761f25ec487d3202644078b8ca513c2e03d1cf16c983ba023951bd5c0741d0c9d89dd210d957d075851d9a240245d87e9bea83f93eeb39a1c7a2478dc7a880;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b9ececeaf1e63b295b791753f47676e42eaf0d9e27de9fa64e18818c868929009411a4ff9753c180b9fbba91bc562d58a7661efb06bae7e7a1add31fdf51d1ddee01279d3b452cce605fb030dccec14b1b33e7b91c8f047f9550be53e674b310a173f9c28705ec1ae7653b6c995b04d70ac967d07a2b847;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fdf368c94badbf229b7a094c97724a9bf8747afe5f338f247c1b6bb4992ea947fbc5451dc326d156c52b9819a7ec78aa65773b304024b1291acd894f349a756d6f8f723a829ff0bfc186c7d65f8f8fe462544595ea359e137e94c710502379bf5c98a199016a57a9447092c9dd97875ff26599cc021925b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a7d5578ab506cad4ca3acb116ed37ca475d3759e013cdef1e79c73207b1573577ee6b1d5cc8fddfdbc37eaf8a61e79324999778934110e88bd2c06d0bcdef08f899e127cbc0a29f3e73d3e077d504bb47886a1e14c8e9a0d016de3bfa8324e08fe8dd355f6520113b3b663223ffbe4f4026fe927112f58da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h682c07226568bc47f68c9121962e233627bf3860fce96926c251ec64e259aa4669d1aa16fc4e6ffce1c745a650caa634816d6e6afbd53b6bfb75eb32c2314350b70d0623e89dea380b78a8c5879640177cc1ce7e99e004e2bff40c18f43f3e62fe3d1f10771050050b70f1c7d2415b41f40081d8f69dce61;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ed36ec5c836c009cf9fc91681d02d6383d4aa0294dbdf9c912d4629e5af608414a998b83a4efb0c6400706cdc838797d74a0d8ef9e7ccf02fe51694e5e5ab08472c60e3f2c9542120b9442e2e1464f5ed591cac284eb089f20f738a394109c99d2d984606c08fabfaf05d9d9fbc966f9ddd93eb89c710bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h354fee268ac7cca1bdf533ad50c0102e84030c356ca967c89b739a75dc8d329736b97728925cd302c769c00b6f4f214cc924ddd9592ecacff30b722f95d08cc26d5fa9ce124c1469dea5a22ee0ac8429c174186ec0b1d7c992fa6bc412ea69a4f4c4f2982d11bf29b96cb81941c207699fc6826ab4a5008d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9310feaeaf56120ef8adb9e50366fa696eb9f20bddc227345225e2d5e36ae9ebaacb1aee059ae4aa53658a73ed422cfb8bdd7469f58393c17aa4b1a3b3bbba319ee23ab916be73284c69f9cd8c7920cbbec5900bd8f2505e2a410caee2610c62e895d2d816a6e9d54c1ba55d7b8c0133d850b16d0fc9133e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102b0771465ad6c1d8df231f8ae67e708f2e175453bc4a9db0d115b901881268124b4c3d929b75fa82782f866734cf910b6962c286b829f07c61ed21ad0a20e7a14be55e145af935a9826f1b3e7a2d04a4b477aa7384f0f780a42f93e4801299e47b010560aebbbea22621eec8c8227fa2d4c9b27d20dcc1e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88c9eece566a0c47ae65ac56f606e6f8e679f31d5bcaebc50fb7700125b95ae595b193b3a49862e5b7bef5dba4fab9e777da72af90e5cc04b0b7dbaaa802c04593eb448738853716d780185a765f56c13f74147d4246a57b4c195f66cb5fefe4f4efedb84a04985e82e88347854f6a58a52c2437cc0d6db3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ed783010674cf31082b2fd33132a5dc8594730769a4994e00a3f9d796a2b804867a4683b45e70d3615a40a3e78e39ff94e33aa149d5cb7ff421cd7331fb448690a30b43140276bedbd484418d85ae566492156dae591ced1f16501d65b1765db4096662775c6c436c8ee1b2203fa091a9244eac0c2c1faf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b168a86f4340c8d8f32e4887d117abb1b85cd81041620e13fdf820f16c81276919c6da447bdf65c34b59c780fc90528abb09d397d0b3279ef4d60041933f57bf2d4893a36628ade3e2de0f4c6b69dcd5a7b6605252aae5a56246a04de714c439c973529c1097080c8b5338401af1ec4706eabfee54a3ec0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bde032aca2416923838943b187ab46c502c739ac3eb7629403096de03ab16f351046c1372133f6bf14ae22a12f394fb47dc5d9809352e03340bccbcb2663a1dfa8bb74652ebeacc0662907e4767d905029f1f621251dc0398e24e07b1e824cf4e6361895b6129b37c711cb818d5193a35b152eca5612e0dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1736064669fdce0fb6f6f43ee17fdbddf69d18a3a98fb3f8c498b3a15078acbd71ecc542fd1c0cdfeec39d9359f81e0e6e9a6b86f4c48a384aca2ece8727d25e10e7fb5c1b052bf3a6225eb1017d10d19eb3812f43723d1eee8da49e0996b5d119106cd6e89fa60aafba251e14403f36ef407f4e7e27425ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da1f8073e65cd48e555c76ecdcfc85a671346914074f00c26ce5c2863807387b7055f129e5b9f1f0a3a5a7a6f932031215d20bcb08729f749f5cb60911f725b3d0b3cdd7f31c9deb300434c8c778f08d480301ef9e340a21509c4e3129b9378ab1a0c187caee6af42962c13a7a32753e1ff4aae625096cb6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h143230711b006ef64dfc4732820a0d9b6bcdc6e85b8fcc5e35ae9b59f344827b21591cd571ad51c299ccdb2b8496b43bf71ce56062f56ee18a55fe20d0f93bb363ba8960421156d224f31a896eac128172fc0ccae5fdf7b70ff7d55a09c19a58c2db68e368e90c27d5f99040603fa434cfa1faef22075e4bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b4f2e8816d6e6eb98874fba34d2110a09579350debab003915561406865de5a02690fd42ee11f1772e51b165082a7e8fc037a85f4ecbf5c71139ec44133ef38d944efc9f1632fe1379378aa624d58098c8389b3347cfa4387a07798bde648d7e6bbf88e0df0773aafcebe7c0c4c83be65ab511003194924;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf50f7ed0a45fd4175e862685f830c52308a9636e0b046d35fe7061d0595de8f082655769082abda2f2670340ea83f6cf0b0c915cdcc544ab5dcd31825d1adc878a16a8e4c3dcc3c8722701de46e96d150124e04b87af9ecbeb52c247336aafeb6047de4d9e2cb6ad4dcd6f86727e11660ae2fc5ca4ef8d81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e5e7b4b3b82dca567976d0b8a0c990f1ae18ae1dfc9bccdc8fd04dde4ec7eeb5e4c420441aa52b32b8cf865aa673bd4475e888cc7e193a2aa197080c37c7b6d0c9d5f4aa8c890fceeef7f0ccb2990520145cca40dfdaeab0c656aef3ac159257e9b6b989ecaabad406f7be9b7636a3456fca80cc1a49bc59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5aed3b1ee17c31ba6e45aade56ef52664c558408dc688ed8e2e56a7475ccae32ae225bb75a247dd50fb29c43d0f32ef3985339d3380516195eb7c00efbf380d9b432598ff1d990b4b9699ad24c4f7d08f242559208abb972c394be7bb417a7e5351b708123beb55b306889063c8d5be7555977c2fa7750a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de54467a73e7e9a92b0d5fabd482d1788635506391037979637fe9cca54164510ccf8c38ac730ff5aaabde734e6beccdb66b1200a7c92ade7e8689704606bfb02c1b0060d60f4e95f02d8aa38494bd2bd2b546071e4d4e60fd16ab293caa4a83e32d960dcea0cf9e08b8e97cf2009a820b254c2f69214bdc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c8427b124af15735910c699d2a3e5bff548b3c3b23fd09a0d69e58b36cf1a7bf749bb971595c04a32b7baac071396d517ddfcf706677e5a8e00f159042aa689f5c2a33be93d8f10426ddd82aa3606e9c82f444d5f77c8c90240562f76dacb183d7f0ca66384b1f640234ab67ce12564a4308747d30244b6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd2d369c3bdda0060904416504752b484a01bd81cfc7caf0c91a0f57ba4742f0090db75e5b544b1d921c2fff475d0036cf1b07b477be2723240b9b608557b542f46d0c3ef3db456b7fa6fb714734a61ec92bdc920e959a619a62878e71d5cf1f668f72b8d62666941bf1fe6b1365ead3a700d8a141b0c7066;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc6a868f061d70decb75617923fc38ec923bede2685a6f980e7c6528fd76a7e2cd917170976d9af86f96d8a528506d5187f4faf966652db51bab7455fb14c566d50f7a4e77211399aa3193c71bc8d7405430ca8ee4374756208570c7c668d949a7c2c2d38bafcd58ed2cd7e7fe0d8f46123b16559f096b47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b050bc16854125f1e88c4fe66383b0b19fd7fb80902be629e7532713ebf5ed7e42dfa33b5334cd752e3adba09f0a1dd828b13a0b6a298b82f82315684b3f18dbd49cccc6ea1597f6feaf4b4553835567e93f8a7c43dd49e17364b4432d4bf27bdd4222c7d59e6fbb852e5b202bd711b74831e9056a856025;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h308e4302785607f3f2f250006c9188a4435a47a7da89efff14a09e85da288bdb6c457d6142bd584192afba9efaad77cfacee01df441075a24ab72a5dd43aae07595226c7024c0c997d396c794e9aff0ac936a9e39b8d2d5b642987b1648e58592460368f052b50e96b1dda9d48f6e08583eae485f4e34535;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a9bc4a2b18adfbc0cd692310b37352a92a054741708c2b1227b4c89552fde696bebeec6c0ce6ba2bd5dc8bfe91e814d1d5b2b6bccb679d4ff87f96b5a27ff626e55501aeb7a2046fe0eb12167a557c64660eb7af7245b8ae5d4b357ee1e95442b98d3ea0321b38ea491fb17da7ce804503dfb168f44059a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h99fe47c4b12a224fec967b7f1d1178518dac22ca8b3e50dd688de61271042437f3873bd49f40125f531e91307f18fe1498b7cb651ae899480edafb6c962a3b09a7a926b8ffca452ff5d420f43501e8775c4a823ec2a2fbc6c62705dd1f24da68363410de8544ea8808910cbf09647d0f6ac87807c644ddaa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc5b6cc16daf7438c132b0254506f2ebf43ba0962029b0ebbb494250e99e0566fb2e45f84e2d4d6cbcc319fede5d8441e086adeebe8845da24035765aad6c43020140008abdecdd948f65a8ec1fd3d90520b7c65f0f78f832e1a1649f4406025daa09cd918ce04cbebe9ff6fb506c2cd51948e6dea2b0eff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h121a9bcafd0bfd809fc8d24578f22836a5b8f7cf202ea89116086d48dc20dcafe9778a0bd27a1c3210846bf2071ef1a60c31469d1b604053d28e0f96158288bc4147a867eb66fe5d526a5cfae2d20d70a792721e5995edc99321800136a68c2b327610105558127a044f61d142d3a7a37f4fea77b0d8cfa38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf4a2a82a4721bc8c76e30f23e914df4f2dc406f758e19590b53de18fbb74b6263ee68213ed93a5fc4b6f251f98644fef6d07c20b3059870486ae8b2bab46e098d9fa799f6ae42b42cce32a099debec984f9dbedc063194eff0b57ec4f77111f43028ff404848283149815260e5f2c43cb0ff7048195836ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h813f6418b62025c4df361e03435b595e7b47b1ba63cd6496142cbda30b3baa0cda2a5a60f52f0e24bf2b14a3057b175be0062989106e3872b09e63ab7332e7c7ee472b3036482cfe228edb1682f97dbd321d75529040666a1d76c1cb36de32ffdb3ca56d2abb5960d0041abbfd0a4b5326e0c82cf1b9c2a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a3953d7ca3c32a7e1767dd1ce4e858c90dda926d5d6107d9eeea4073683a479dd793d9d4fbeab37a91b9d6ef85adc21699743b39ca30ef87615bf21d2a850d48dc6ce5b6ec64b58f7474e9e01f75ca2a4be4ba8c6f14a84a44d18de3cbb912a9382dd99ac772ef0186132d91055dfb5f5c41dc051068470;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h189cd07b75166fc7a40e2fe270881f3a71d27a7a27ddd022769bd5aa0fbc853f370fd99591b33f94462eb50235f8e110e89a37012d7d5d7fc03f58c72c2c01aaa846cbb11d17e971661fd7e06dfc60a0142780ee966dfa8b98f3b4d3f0eda50a87d61cc001d25140e0a655fd7f8d2d5fea5c01cbb66ddac0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha26c7ddc981145f692c09c1a7a7dc9a0167c84011f6b8b9f35e797fcf985335a3301271e78291302aeaf76e8d60ba61319b3cf4ac68ea71bca93d764d87551a0f087762594fcc72cd88a39f133cb3c734a35acc6f96bf04d8b2ebfd39af01f8d2343ab0e367aa2a0cb36479b14f491064e1e30347b54a6e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154587ce8590f248304e538206afb9d6c3e05229ebcc487009b681d1f7f4c68eba76e0a97d2677491e425bd57302ed26823a434f319c3830f81f06d979151ae20ef6b0e754530370cdccbf0755093750e3f368d50232535a696a586efb5414b23b85b29da44654007a0fa0a911c650cdd3a170e0842773c1c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1094a763d6165d928a1397d1b2db613d42314405fa61b29e897aff0424d97ba45afe08da04e300ad9a8cf88ab283735d751ac22bd3dfe7c8df63556bfe641142a2481161109cc75bdad9a0882fa91916c4c300bc9a30f7452609bea5aac295f328caba8814f17c375be90cde92987b80403b7f02a6a218a23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168d7ac6ef82852632ccc9efdcd57604a57040897976754b1c934ecae0536cdefde096cf7677d1199127407093ee0479774333e67a40e30c091dab2ce2b156e4aa95240c310ddb5aeebe85d4f741d88b2c69323c5b7f0693b0a4d48ac0304c49e6588cc4a586826fe7df164ed50772940c9bc219327a7b3c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h648f654b65cad03784b50ad3b6c10f0b5eb24f683c4ec102282bd3ae0540f929ebe5103bf73e664c6ee484198d08b4df242a00b72381a14fe8b3239ad7f0b6a6c17b57e888325a91e443b099125ffebd192f96007e3ee116783ee9a392c67f39fbe5d124ddd2d7be6bb6202cba72b536fc1e4723d8812caf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19d58ff1c0cef942c1dc751b30bfa2ee783c42020cb6e47cfbd5e6bacbaf6dd498e6b2b860135f1810ab76ce2d0dc86e51119971547c9cfc48b247f2e34e719270393074ceb0fc117432830cf64c1b9ea878a24b003555fcdecb59a27360a1045baf2ddd27aeb3c24424e37c69597a092486a98af2eea0c57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1fa06e6dd7700118f8763678120d2916b177eae306856829eb175f9fd9cdada54408f814a6d476cb326a6892577e02fa47f197b34af7089f6b79e5aa9c23fabb3cf1374579aeaed3e02df1abdf21115e3353f36ee19e015e28594d25f65005ec11130c68b8081e681adfb0192839b9b6a857e5f432ba2bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h408578cf258f8391644fb2b2de658ae1e889dc68012bf424bec1f7b582b488bc5617f65d8086f8dd19b1bd78f7b863d958167711a7a226d7fc5e47f164d2d3ddce8223d052a9f0cfc59c520e1908687bb5abc24d10b6e91cc3d3d17f3c2a2c84d77cc8183d47607fc930854266962b89779b54f231d0b9ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb865948ee2b3b836f4d3c4f75ea9bfce79a30b59909d0ed24e41e6c3711e0dd29c865aa2ab100acc6159db7373419f90b16377ea10508dcebb87da2dee9a843e0e33cfac5683cf4fbcad70995913d21c427ba339a451359e7a31f2d70b50a8a65b8ade776c0bccf487ef6342d4475c409797969ea1d6e30f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e78bc9f76c953ab5b29da2fc49a9f14788ebbb57acf5717353ed45cc9b671e8c400c00237197cae2e979fe3aee851459e25e13185d805336725cb1ceccbfdde92d9a556560c35976371aa80823a194c28815933d6f3edbb4410c25e90f360e92acf4ed5465114495bc389fb4a5490405f87a65a1ba74432;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a6582108a1d5bbb5e9b5778af3022a70d3e1a1ac75844b098a1593cdb255b76a28cb698112a0859648f9ef2e823e7913f07203a4a251f5459acb2383297a33bfddd6288420a9af8a38139ccf6dc9a0549ecb9875b0a206ef66b337cfc9a06ee179f8421e793083c9001fa63558b83f658110b7d4ea44a3c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c0103c7947edbc83a0d5e4308b3d6152557bcf6d7b7b41d819b663502ed6387f87611540fb0b9f3f44bf4177ea34a989565c2c269ee9026a31e4f29efdcbc23f1ea148b3af805dc2875a8fb55beb2300f20370ba226ec8e5e187376b288c877bd9b6e51fa2b5cdc0d9f9fae6261ea0a8f2b09760934a3799;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a71b6404705c334aa16d671e3eba09efa93754753f21e8a1a895d3fb95a9a393dee57b8779502212a1ec56ddcb146ea8dccc3b8929c8db872bba162c201c51a1d6f919d3fbdb4358eef933c4ec0f73cb8071c03a2f19d08a0c1358223bfaf61706848bc4b227b4a39347eb36261b55ee14631e8bf695504a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc218a925bf45b2dd6879bc67d30c0ec2814c386bb3a6f441cef5437faf4bd09b81c345e374683df222ea0a07386f772d3c3a0eee3314cab1d18c36ec233574eca27b0394cd1a390770d7ec2aa8a7d7c3216959af3438a9ffcc2963f5272044623fd5863bdd43096df7c16979fbb31a76363cd88e699670aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h657d4405140895551d93de5b00a594d7a58bd127e68532d4a171e24adbfc681f7a0171b4715c4a943a9d2aa454fbb1c1a908ece13673002773a5aa5a02b8b8f6dc73bc468743d0ef5cb8e9d586f29f4810d8a2aa2d7c33155df52823205e272ed905835da68f0d2de097ef7db5eac6e99377de812b67e8ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11cb026ad910ce462ee9fdff3123303557260c5ed8009b9dbad8cf2e2c547401c08e140a18298016dd8ef643e10362c62f87e2b06c7a8f023433732a6676d7590b18a82cd05b913e5bb18284f3c9107802ff2ad62ecd8636c13445861b22f63b72973aefbc4a2c10ddc0c4cde29a6d2bc881486d8c7cd0e16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1df284902546715c54350a74eb8ccc784eff617243705123def30320fc6d9ac5fdecfb869bc5dcc8945c34662630d0f92aebdc91f64b9a7bbeea13e92a982d5cba7fb422e82c5f99cbe9f1db9e5cf38067a5659cfb6bd2c00704d6c3f0e24475ad933b4aef5d75ba2b92a377c9c49c4dd9ba8a14aa3138b73;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1173fba0d67e2b581f6a9967b89a2b7b1b730a737e6f3378ec750671b527ec66087ad5525f7faef41739d7708628d8ffad9237f0f7b25156a7df937b0a2b0b0d8099b767d95802cd161a6c596ea0e04046e6a97f1112938c464d67ad39326f1fd5b54cfe6026fb2abff20829fa1ee8e1ad8eec83f47455095;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b94c98d845f22d83e410c21e8d61680632ac47a56de1c97f7f8a3cf3b97a80f9a92b2441bb9176d804b2415aa07116f537950bfa8b31aebd26e39e8ee86a7087540588a13eeea8baad4927796c5336bd51cbb3cab25a44f54decdd931bf6c8c7fa59973fa8c0f693d6f047ac10993675bd5bd4d9b78bfad7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5fcdc28dfe6f1fd7ca01290175e1f8921f125f9a63cf895575da457c2d48f5029193e9e0a445b39dfe78c216ac3108f385edb15e00e7dd3170f5d6ad56b56c21eb8d98a2a204495ca2a318ca7044f70e3f60b6b85a7d24b1329480c55f38fce929d6e3e86cd7d60ad912c90f0f506f541534f3ac60b07c4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1464d5a7137c2e682ab1277c09f023fa46407ea0a96379c67922c4c48b935ea2c31269b735d6a65f585e08ce9d3309c348a61b3e6715db76c668a9300015b66aff68aa8d53194aea0723b7624a84b891ff3aaa3a4ca7c5546b2174028ba9292e4dce6ad53a3e5173877edd7dffc016c82b61fc352a17c12cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4caf096ebc49f30e5af42976191f37bb3668560e3d70de0d856f2771d72de93cda522dd3135cba9c0cdb2875baea34706c92b99c58629d256d4682740bddb3a838904ddd0fd215f428f2b72f851091b901badb9e994bbb8f6d05f4930bf5d7b4e0fec74329673f083b3b5dec9c2e0030f517ce47f47e3c16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15588ec5a84ade00159135c922d1990db0ffac7f3de065854f1cf59b58c4fb2bec99dc2cb2916cff3aefd7bdfc1eadcb2f4f1b582f79c34225259462ef2848d48b159f2cf888941638bca2606a7cf4bdf7a00707c5f9f83c31daf23d5fd07fe544d643b33f80cad3469443ecd0593f6ae7fd45baa2eef0507;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h136cd78540c1cc2e45f67552d000a75406b9eb5f54cc634ac8090127f4daab5e4a00f12dabca79df710263712d498bd7a2244cb531e053dfc21a19a360621417474cb616863fb57736be6ad08138f04bb3665978d707c93cf2690411d109752276f378f6c4902d8dcdb20ca1da35e1c8b25877a9319c5a3f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a654208c101de16866509cd6a6634d73ce9f2780edf3f1835c0489219b8de0fc92211472fab2be3b079ff8ab585f270090ce54f475bf038a90d24ce3fe77b6bd15affcb12facb90f2c87a1023098c58c471e1a3b63b0bc450c22109027ce9ffe53c4c2a398375d30441e7067b6a7d2ab65f6f22a91faead;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c64e9056e159debfa2d6f1f553a764398146c9ec116bbd9c8d9d49e4639b881ca070654458d176e66dd1d96d71efe5eb400b1a2d4872b3805ad5ea8aaae3af9f487872f3ca303a391ef1694249b9b7fcdccf03b6b49fa0d931e86b8588c94e2d13f6458a32316256a2d96b6ecda45923dbd21945015a313;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafddf3bae2201a67d92153213aec6d8f7ec60674d6b7650d26cd5eb28ef153442b1edffa5b31021701bf4fbc789bfa134951262c3bc8c020115e132f93c6094b059ef21e508f9be3075ddf661e62f038dd14295903939a48b74205b1cdc7325fbfadb1888a9261ce732da9ce72b9bf1502a8b5e2874a32c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8c9fd06000a391092dd2fb6b7cbb70ef0d7f0f8546ef222c183386d397f7c69bbfc1e3a708f6ffd7ac37edceb7fe65d461a7931ca8fc2718ff0849d716bad5a83a302a9e427b289c7f79bb718ae299f41afb5c184c463e70d864b59b32405698212c4075cbd84f738a716788230321b58e550b640cd427b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef6db58fbadf09c86236257c6eb82932d43f01e447ec866b9f29a4cbc10af744729ae276f15c4f5cae0d464fffa2cb36d36f4b6250e5a2d1a6081c3bf2b282f043ff59c406407b84b4554630fde203177f2495b5e511685be8128a44dc0e10328e7bced9b36bb2a8ec972dba474c11c02617cafc37b83bed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haff5f8767344aa6bad614aa0491c1c430e3efbe1ec057e0d6a0ca4d5c1e37e42f1fa2a583895d6f03ba0853d952ebb8142c058fb4d0fffbabc19e95e2410eaeeb305e4f433d6608c72c762ff67d87f5f8d053b9af8c98cc6743c5648449d6669ed339f52b7c974ddd5dfff24186fc09f7f35d4b49d2647f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13bd2bd01be27fe9df1f0e8c1a50717d1847966c0cb7ec7d2be5d18d8cd34a74f99fe96d6565ef5cc986f9d7be5dde38490c880b296aeb99a7e9ffaae266c080aae708dfc6c561c74195eff87d5928ebf3da901ecc00d244ef1b4bc86f085e0bc1148e1e265c698b9949a86dc44ac86a750882c379d19f091;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88716da502c14de192bc2e17fcd9ca8891c544c36ada2d9048915838082bb7b670388b879e4735894f454fff15244fde5a049e47a9a3ce830b95135b97761df3eb9c0bcb0e594ef40e1effa13ba15aab8f0b08d5b2f03a7dfe96a1b7f297296a2c65aac656eac5910475249ba6c27b56f967da5bb995c68d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6fc973e89f6ae9ed5512695fa57e6bcacbf58a1a07cacc1e9256eae2911f94c3d20beaa434dc7ad166b83a6b1e865d784cc574c0ae0a4c9a020bb5ef5bda52cffc96432b8c6b87bcd84e4399b30eb7c6b858f0c6ab2675e2b82af71005fc3c3f1d463ae2b97a77a1bd90153d2665f995ca46d2781eb3986;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f9839e9369281732c550014562009c7480ea433ee405fdb5f8d1f695001f16616ea7dfbd3c371d2c31ebbae6b45d0bf4e34c5a8ce248ceb2f2b4c937a021c5a0536b0e7add7b19993d02657947430a07733ba86ddc14695dc29a650a7e0432658b2f2db8fc1741e950b97824f6f6e4fc83bd9adba155471;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172939c3f0ee6e4358c48c2faee60c798f3defbd146622cd5591b288b52ff0e3f6368444aa187d757f9e922e093800a5dad9d103f5865f543d85247d80693a7eae1960c44dd946cb3c079c9b5921e4ba7490ef7e6bd5619f9d4a381f68e11cc84b46d61d9c4d8e03db9d4b7d4434c06407216c20fe33db123;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h338c59c51fe3d356f3be4dba685596bcee7b47e96576082b8a3c9dddd14450fd8110a973ce5937027ce5d6a4a86c5c89dc4a8aa3c8dad8f314beaac8574ba072a86a6f2c0f2946967648358123a5e201354d75b816b2de1e00990ff4ee20fbb5078e09ffc1d255083609dab98ad6b19c80e3377a5ec4e70e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5d6f8cdc2ea898c8947a46d1594a1da180177c68d031e9af6db8c3de7993646e27ac415531dbde9439c415e064f48b0d7746ddc608d39f71534e6dee6824fed730641345578090c076d3420b377dbdabcabcfc3df99558b6b1ebb8caeba6950385e611959d25bd7b0beccf27af36d26e890ae10407f330e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b2a3d9e0049e6606c4d91b422bf1380089c8ec0ed3bed48f25dcea1864be823470172bc3865dedab554209dbdb8756b34e8bf805e599a4fabad16aa14e1b61153062b31610395b9434c6abf0ac6fd63e9a9c8e24b61279c4a8e5e07438470af11a767e4702f225ae8bcc4efbef2ce24d2d77db5729a5fa8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132d07e61d3359430d15c922027ad0949f54cd8356bab2a1787a12033f5b4fd815cf8ce94a5d1b1dcbaac34182dc2974f4c1c8d1411a75a2d0e3570618164988452991ff983791534126b7df73c56a71f5b9f37e4fa0a831e52a2adadb23a31578802da7275af59b34757dc619b26b5d937e85dbb25f074d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda46112f00499a2bf58b4af6f5c8d0c3ccfdfe8c1e06ac1805285b789d5fe9c98351fc96d85d4c996d556b6edff917972e2388febf9db7e58cdb8ef129c7223d3811048492894659dff94edff622da288d9772b4f12470090e4ed2892f0d0c5e551e7ce56a67c5bf4493408340527ea85797f1d97283e78a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac04f2a4e15471f94b22ea9b83ee31edfd7aea902add071bda381790e6d302787aa59b4ef05c974d570da258cbc5e5377908baf3066cf65543a7a11fdc8200467957b3d3a6bbbfe2292c1bd1037db50f9a091393192ee98e33bef06528e63e636284a84bdb5e01aa8ef6e4bd15917f97c1abfe2703e2221b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa520b7242a83063f01e8baa7dc3119772ecf98301409f18be36a17e1f31174d8e5061e8c099e5c22f0a1a90763b9aff71c23bdec9ce5c514c4a46882c46ad56f8326368300920f9622fec65b132ef5c272066123a422fb2eba7b3dc2f2918d11d153bad54e8bb8961bd3b3ff7ec00a5e0e716334a08d847;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10ee136033b1a0ba58b0694f809c9b5df4c59291a4ed125e4381f9e2a989498003b86a80b49e138b297155b856dea1c9fef1c4f18d82951000632bce954b89249e83675d802ecff20b0f9ad9a6ecea323a02b4b6fde5c2af969b468e7f1dea62984222f29c21cbdb9308ebca4a06a079020ad2a5fc7f78470;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18af43bbb9c8644d79ec37840bd39d1cc5758529c45d2ed3938743f8519a50bc590ebb166684c75c9d3b02748f9c23335d13e407efc7566ab2df3fa2d1cfe6acf37cf8dd035d45e55d865eb12551c7cce93e66c738f4512b543b62f03d7029a1701da59da1d34e36331209f141b7cdcde9b8372abcf06751a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h69f1afd6424b6e7bc696227d4e10afe44d86cd9f6cd6c909cda12ad33905347dcd0822d927acf6871b5397f174e781ac1c86be889a3917b56d7a2c91d5264e19459d41b80fb39138c77090d26ee604ba9f8cbfeda08d4c35074d93afcd63405c299d3d1676349ffb168313cfeee7bbaf054c745c922a8d92;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67c48a88238d7e7a91fe8ef2ba7dd63b90a6bebaecafca28b0a51e42ef5aba1c1ac3e2586567658331c79ba33f020bb36f96b76c40851e43d86c94ede715ae5b4d990d0e167b98c1dd34fca108ff711a9d10ae0a990632d53e8f786e5fc932718e1290f915b0437aca7f6bc4d3070ac01ee26d66c67d1c9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca57ba9a625474f03ce5fd4139007142fdd817a89f35dc8bad06bce0cab614ea6c9fb0f269e4130cbbb36ed6ca060ad15ca0aa7b2dfe2b5c88c52137b6bd5a62698ea31dd1d52e55e54ac8798d4411ee95440e1fd4db38d49ab7d5f69fdd8db0b63d1d4d3d54d4f3e17d9525e81dc5bbe427026755c30c27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f2a9e1b1c74cdc8035362e8797ad00d8fc842a4fb228be5db5f8169f3749f96936378f67523a9d612ca12914109ef66132a237d5c72d342c3b9e32fa14b66b1ddbaf2cd71031d7fba761ca623e35881b0aff6136b2877988995718aa6aa96dfb47308288ebabfee51a5eb6e351680c7fbe102ba312116c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14abfc586ca2d9889cebc850136cac2500a6f5d0962cfc97c5dbe8cf01ac11eb93906f29a65b2d89115513964178bf8f3ee89a92da9e21594fab9fa0a5922716a50350aa1c1b9d11fb1fcabe0c0581f9e7f6bc65847ae72145d0ccab225aaec87da80dac8995f5844623b898ac29425e5de2978a8101ffd91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c78a0c402f46cdfbf8d00659954ad15cc681be99141ca3d6c5ebb919e27af66edbcb714f693c4339f9937e41097f1a025b0aacb79ec67d9990f9f6896c7dd00626bcf050109dde93e7b5394dd729115ff1f333757f3296508aa2394b4b8994cf3bac2a1265bdd2f62b538655a396de1d8dc57911fdc4cb14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4fb28de36d33b429e636f627298c84603196bc86aff1a28e0da8a4baabb5b583ef173f14ae59d315dfae72bff0de2722751a9b7136c26cdc2494fbfaa3ef3eace53a8ee72cdc4b636941ef64c98e984009ab0a57bfe83d66730d218b450d3d9327ede58239ca4b263a85b63fe70d2509267b4e43c9f149f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f482f08e78e3545bbb672d6556a03ffdc0296c72f2fe9e74dd01e9794c4948c8c7c04c84ad1e7166487275809f049b1e7499f2e26fb8eeb6bfd0909e7154bfc19479b45c58906f3635df224ab1e3e8ecca642cec57240958bea2078f184026c0d99c140b3382ec7b033c1e56f0de88bc77757ec99731ba7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b9d6586fd5213f380988f6ff36024a9fc39449bb07763226afa0e9f9dc641cd4d10c9393f8219ed26638d6269bf8054e7c4a84e564970cace7e991a8e0757d5b8bf6b9d8421770d015bf661742cf6d5b3ffeacea47b3bb630cc183041e529615101ad775db9b717718ab053f797c7d2ca203c381fe38104;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a6f7420338a357509775993420e2071a75532752d55cf3a90112b6046222539b2a27cdf9b1ce7fccf84f58ecc67944ce5159a25f0becac282601de50118cff4913214d91ce5c722cad19a35595258f2e353f326ec601237257b80d92bd564ebb1112524651da1775a7f1c1e28ca09dd155a2b2eb69b75df4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heffbd6644a5380fd90de81a4999a42df581aa4e5d1b4452d47dbea7d9aaf513581941ab6a68cc8a062d9703da088e8247d5e6a0fe943ce47951814f94acf93ad990956f76c128074a79f686c31a1297cdecc6c49d025baec8036ea6a217288594c212966e7b7f477b7f6cc25cab16bec0b6d5dffc003935;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79fa1a619159213ed55aad07e21cf1dc24fc1681daaba6aeb31ce71dd1ba88da154538a4d051dd8af8f0740873ad595e8740c22484dae32b4216a0fabaa5ce885cf02b7418d7bf3c350cdaa049060717fc3ad1eeabba323b6467e2f8d2beef1f59ffdeb72aea7107bbac24e937a0e3e7101388cdb18db9e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b06d8dc62371f7db187c72cdead2cd6fcc97bf3acb21f9ab6f1955871cc644c1e11ac267e105dfd142e5a29892aa1358c681bb65b58d9002c6761e2e6ac110d0c52a726b6356e086087d571551b500f9ff02a72caca77a4d4bd0f2740383b3d5f3ad4b5783bb4d36ca4fda681cc79ebe71a392f335f17d10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17440e7c9e9261185f057dc0076ca0ae9b126d0ab035268d1730ebe5f0f95d9b12e11c54b5dad12c66c2813c1f9cf88f00920b1f38efe07f8d73e5ec27a823baa1d445ff6f2ed5a86d4251eefb23cf420223e08230f04d0e6270c9528a1988448645c704e92dfc6e5c959e04ec9efa468c5b180ce4d1d0b47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f5f0132e524796de57bde6b8f99139cbeb1f9fbbc362ecbe1bb747d6ee8b62f38b3afe80c265fd44271db5e7d5f889640e49ff171af4a7f4f5bd87aecc837195e53ecb2a05bb0c2ebbfb9c7d2d8c1862411d4022bc2f1d09d2396628352e423f1de001055874c3b65c190312003715aa3b022fbbe76d4fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc0ca435c2276c839b27c5a999bd8fe76f02e4db0454e231d4216368dc794f83ea195b03bacc6d32e23a1061114da4106e37fca1bbaec91c32eb759b6c72b5a3d4fcf4b25734386e82d7cad077c404dc8d6f0d58a937336ffca6ac3ded4d10339aad6823cce341deae79ffad22865f22790c5ac11aa6e291;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2a1bb4d3188dc01b154db62d297436c5fdcaede362d7469bed27304ee341c5f49497762aa06f596ed69e70c290b0fe9eefcbc88b601818eaa997a57bd4bad00addab720abc35cc317c02ac71233067dc0b6082723d7e24c059b68a248108444dfdf30ff30952aaffef45f301aa128bfa49d93cc33081162;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7ce130fa08518cb25b37be3ae8ef13af4015f61ee493fe3164a920129a814a9e0243085596d090be95ed49ac78d6206234d837dfb1d36033be157aa33dff32a7cdfd51086d21963c27268da11c50c9093736d6a859ef7d256534c2da46bdc7de4b4fcd8caafd1cb0a0abac2859c96febc86b3bc9fc3ddb57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc666113bb5b69c8139898e017dc137334a36d2f13f40f8e11ce16ebb594f092a1e007c8a4cd6cb0c012645dc17e48718424ad54cc53ec7a458952e6f17121a7b774fef79159f972d651c9b3de907dd38536d197ef5e6b7622bed266fba241d211e0ef8cc8516dd33525588bd6c6235bccf2deac14ab57dfe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4887584e28c3f33463b1fe5f48f0b2137ca0c043929315cc36a30ad2b075d1b25cd4b6df89529fbf911bfcdd0d1e42fcf700cd4f795080ae86e0cbf95be5f726d47813042bc01d910037342bf9ab9290f380f1e9f4cfc8cbde8fa7416b8b0b33859192e064b7be896831b0565ecca814eca54b23e3354c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d8791089907ad4c323073ab8a41d8eb2926893b44c9cefecbb93ac4f725beee4ed5a778805390595d27d79b636ea9e2993f3167aa5553e39af2ce37dc379208314f89b6a03fc7ed55ccd40de3a5696d6afc4c93538538b4ad2a670069ce5a39814784c2909dd4f885e592130463cd91f8d3122d4f115073;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61df19a531762d1c4576cfa45776290dac01eaae8a79ac014708dbb13b8dddf86e62cf54df13be71c7766fe5fdbba8685de09369192a026b95b1d63e52a0385ae91ee94257daf8c094a5c8c24df5463867b1438e1e97129457f24586809ace621fe4afad351f9cacaa81e87c2cf0dea1fae71d4aa633070e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h153319a9ea40cfd09205c4d977b573fc1f90e2de46a4d4df1919b5538203f4b9a9eb98e788c7723bd6a72ef732b7fc3db56aef2a6fa1c5d77f759e15928b001cedf9024b82541b248119c4b8816b0d5d8ffdfa4a4b0238214cb061835f37e531deac731d72545286c3866e0359bc77ea141392eb824ed2fc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c651dcef3f8bd5918ca6f7ddb64170ef33c717b434f1168c9d807eee70f8cd224cede35408e0198ade7230df31e2b9927ae0813ec3d2cbbf65c6e5aa8c2a608eb16675ae9dbec930c5067726229992f63a93b868f0d5b2862e3674201bb146f93d74d47b179b61645174f8804f0c357e605f71c3a70ca2c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa8cd1e11a7dd7c66f73161a1d184ed5eb2e3d772859017f8e1e0306a438cd9fcf5a3489d55a69aa51ed4e47c2d7e0dee8eb258c3f2ee34411331a2015fe7adcf17bd16abbf47a04226f52caab2c24a329204d401cfb672c172a53032d318c79b3659877d32c663894f6709ee268beb05dd02c95937a4b5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe9e4c41f38edfe2dda11a7e1c51d9dc22d949bf4674590f067bb70a0a9f235e3b1a69ce2a9750d2912adc02b01746a83a1c92adf68b13e31e8b703d480be4dd98ff72be51a4377c3445a035de0719c2f09dad55462f06940fd34439d8aa0c9cd179ba455792c4b6e4cfd17ccf36dddde67825da5153b76f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa43b4e8e7e7f95718d0761d4aa84a85575a2685669748dd7373fe6a43943ebbec2bf004bab74f3b9be5baae5186a0f185f9be8df8c3a92e4ab99d3352867eeb37c872cd1d6d31d3104512bec86dd5ef663ea56534e374c028ca34f5c61148f4fb9942445c21f0e0d6699d8b54d692ddb1c0cec226574b85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h86d2a7827020b600255f1a130415c4b73b67936d25deab0704f033352184d35c2636d61eb25d9c00c5a4de1ecaaf0e808bcacf8239b9ff124ff85fac87c4734fb3404eb76801eccecb07d655a951a1ecffcd5cd608d31dd09f5d1806d2896765b14faf5d1d9f7ca1f27195ec9bcddcb1ee26ff9e9e4520d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c0c01ba47b79b38b9d6f2f354c2c0b85fa9d067e1e33d063ee2143a91cda3445580ac02ab3cc35f4496f36e689641ba7d4d3f4ab485e44f7714a7159abce25bd6a4e15852bf543454e4a9cf7b42c2489d3e2e8e471afe410b41e5122a31b98d9fd7e10a961447a7fb27e07cb3386b616e91610ecf447ab92;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c040cc15f68a550396a9d3a22156666a68223aaffbc1434b50e90fd0c681d89220e1bd3368d67eceea88e00bb0bf1b005ec18abd7b5afab1fe21347e0ace7e107725e88dd0385eeb98593b9ff1cd37eb0617bdceba9085a0e1be9756f881abb9c7f4dfecf6627663498ddc43549eb561fb821c481f7f5f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e63cb16ca8f183956109cc1ea7cae730ecc5c9b64972667920509e4d02a5378159463422e2721cfc114359812140052d11ff5c33cda004e38f4cd000262506177a0daa195d2667fe1a1d475fd08f95df872d5b0708310a7cc1ba50dcdb1fb6337a0f6ddc3cc28f855555fa65d4a6f76813d17440e37b3dc4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbebb2ab852b1eeb8aad6efadb1c6e2bce1bae3b77e75c4f67dfc908ee297d646a821bc8a0366b4382a961f42ed2bbdf7bb8245df313a39d0306ae199f2a3efff1d63cee0376211e84df4327c4f9b3a568cd7b11963fc07a1cbeef6c87fc301ea5b08f913bb7ac3e20fc86d153a9702cd777017bf811b4f8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84194645847aa2cef77b632df31b9359afb718269ed49b246f5a7d69647daff49c9d1ab7578827b2d6d66d77b0647bcb4795ef2b5074013bf78022693f9e6899c18eb12f8baf4c1d7a31d3732e6a6ef08ced9f2a1f72078a0b033b314383afece42e4c1bbe83bb6886e470c78aeb0ed9718068647fe38c05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf0befa1ab3baeff44ea97aca2ef0c8da9ccde7577ee49d96cce4e1c141d1d58570033477f53cda0b201b0a0aeed8e5970a3909972016c75811728a9f1ba24f30dca14823201706082fa6eced1ac22ef452ac238cdf07f0dd90671e24c1852202d9e7090c9d6fa29fef3d2e7e8ffd8d61b0a0cd29b6004cb9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb21aec721c43416c1fd8d5a5ff9a824eea4aa0bb7bf646817654e9b2f77b6633e81d3ed5f0d88669819423ae035184b4aa1fc4533f3f0862d811ff44def7f4b0ff5f683b2ee8e9311b361f8c80f595f421f70010f7c33d4e9fb59dce472e132785e8c2c22e36af2a3a553076dfc320a1bb7446c15f6de451;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ae1640586ae7601e1144a9ca7726576382389b0db7ff060ef7bea654c1ad29911ad51b956c53a77add80a69089d71e1b3128cfbb3d09eef33133b0f0b4c76cd3fa6e7cf2e2d7c5e3cd6877f5e0dbe7542fe0c8b56551ca8208b9bf2a6277202d8eff19124a00b8f218245545549a5f4a8a09f5e6806a5d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb1769b111765606f9c90048078b9c173cb72ca1701d23fc3943c9c3389fe8c6c022d377a75d70223f877abf4a58aad01e4627434128fad5a60b6c42d7849d7f70d36dc812a7dc785cc9eb3e6302d56169521647b15fa91ea2490bf4d3667e43229d83b35a4755f6668dbd127d1cbeecdf0faa1928fb8eed5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18aeaf16e2e68f7b8a43841ca562c45381f419d334d46647c96adad12ab05a0d1c21d997b6390b617c613d29aec2182a54785396db78241144b01c06248ff87d260fcb93d87e5a5896bb2b31f0f67fdae2b6acc20f6e3cd09a087d712c1b249a26d427e7736f2d2faabb1159e4afad3a65e722a059311905f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hede1774e4b98f99a792f6cbe676534aba7aaec1134972b0196349c5bcfcb82bbb13a654716c7a0c38df95dcea5bdec0b98e8fe3cfecdc8d79d57dc6bdbff82b849e0ebb6d947e328e66ee4fbf2c1f3725b82eee7241aa5b46a29e320dc7f8c967c3507b265ba90bc18d872eda9799aa56b1c1ae45869f9b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a7c3e3525927a61728ee69058839a322aae30e33ea35f40269d4bfafe5d59df3bc59a57a9f71491683890c0e02c9e88f2db611892dec61138a103252de44bf0fa7568f4abb01269153b3e4baef44f227e52737777c1b7cafca5cc00d93d92e4dfd7e6b1fa3a062dce650afe3d043e148b1c4b7c1da6b47ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c457fcac2eac24991cb52d7665f277e7bfcd761d7a508a457a34ac67c5df7e7b1bb83fa62ae87da88168fd6dd61054f8a329c701ccf0d2c4c36ef1bbaa7880df0747e6b8924edcaac3960a932ed349994067b718a6a2c335283fc151a38e2eba897bd4874fb84a8f10801cf87a532db08fb685d26324874;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb1edbfc664259177f1293d0c99d9533009c823f7e63818659c6168f00827f91f52c79279f9279b8805a3809a4f8f4eee3818547bbdf04e6b449769f0d01efa9a0cc49aca812a0b26741104bfda26b4e56ccd738359b2f87459f7351a8c6a6e34deb37577dbbf1685d25bb17b490ce00b5a68d6a566b09d33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14b1aaae8b57df45986aadeb1f895038cda078ff807f4ab0cde1c50417af899f395cc118497060f9aaeae79e8bd0a38da4ab4f2e3378fa643739b303000749ddd44b7be7dbc859e905dc34a214b3cc8a61db153366c36d282c2ca8ac648a4205ad6e9ece26d9554805c0bcf75a24fd54053c0b366b309ea3f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h431a1685de627c28efb961e7be5eb5707817d92fcdf09b6c225b40b7ff6c7680aee0b4e45d47d36e46840e955de0c259bd6ba4d9954bbde86221dadaf711d2b352012d413b40a8abb5a774b226ec691b8d4a117bb2488c29ce7273d0529812892a53f66380b126c7d3025fce770e9814bc36249d70395d5c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160161c4d08a91782ecc777531d9dc35c1c0df7b4a574c0b241ed6d526fdc2992b88a953264967b4684acd0c6d6914bc0f33dda00f651fcb7b5f2105d8c6e0025d6dfee39cb6858c3386b6e28a62dfad925f5ff22506f6afff1a9129e4ea3fed4f82649f11dd58603c1ba388e4a4588691a6b6d2e87f8a320;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ebdc2f25a231882f18a73c35135c0fe10869191c1b6036a53e76ac28125454e57fee71000b2fb09bc711a7c890056c1a1a79d0109d41bb95806186d223539b30441a31b2259b981eefb3c3ef5d8e2f255484837c974132b2f524c21b0adcc0822a69c127b5b5e98427b90dbe95807b1b9736b84a415f0ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1811ac0f66faacef6958e04f305de57cbedbd7972c5e7e429cc9d69c3dfb82541e3f4f1f45b2998d47232927524c0dd11a6fbd51d7a61b0436629a2e81cd45b0200273c9f00dff359fae6af2b36fd21fea00cb8de177f872b6c2467c6a60a99f7f2323dda22a610dc3b6558e84a2f83f202e065c4164f8741;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5f6293270c9e220b52cfbff075581b7c622ff591d7351bd78f3067332bd243dac306ba70e2ef13aeb03ed6e57ac0c2528c1dcdd6a0d40e97668feedf78c667290a34ae5347d1dcb97551ae806972da5dcd489eb853750fe85972c0d32fa19fc295e123097279de138f2e6e1373b82dc8c42fd63bf802cd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea11b6764c30aad2315b1ecc4af37f41325544bc7b947f1a4948ea273688be30086fc6c5bce539d81c746b185a69c9327b610b0738f6afc9439af1720f8d561a694e689b653b97d71bb7109e4e07fb8a4a8ef115ffd515726e1f614384e477936fd1eb2b1ca35f72e137775d99fd31786ab0d50c65162196;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hca76aa5d75d59bad148b509a88d28940f2da7b16e767f799b2d0bb7102c0fa449c4aa04a81bb2acede5aa503eb35a13e4ba9643a66858078859e284c70400f6ae2992670f3c07f26465590d8e751b05fb64159cadea18dd03f907bec72c2425021d248344680881f6bb3ddb090f937d389069f732c4a709d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2189f52f48459bbd693efeaf5aeaba9f406b63b672dd1eae0d1e663926b98cc0b8ef1251520595d654561c48c8b22f76a1e29907d336533869d202d0bc17e41373f1b44f82808d9775bcc1f8a8e72a2959bd0ae328d0b4d6bd1e5d4f0bbac780f1ab2dc06fa6d6e10594bbd781f24c8603631ec86583bc52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h341602fcc69e65ef9c8b3f556cf5894077131ed4ae0be961b0c0573d04cd09e536d262f7e3cd8a01e26c6457004475467572f44fa9562d5d9aa53a5c744e229d97d73cf1ff191e095f28c12e2e88b3427a943931737e1b5065318f4e8659f6a37d76d2645ae03f18f9fb85eed713000d6497f3b14c636152;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h888d2ccd6229148df3651880a3c3cacbf791b7a1920c19fb721efed3f708d979fdb933e67fa6af8ec48de69f65afe1e96a3cdb0fb714e19f95b030ef61040a13ffe5a85d41e462678cc76ded1413a34d75283314f1a4406a92cbbb58fd1db4c881896299af83dadd046cfb7ef8643b4e00d545b799ff43bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c39dd9173a4d0e99c6101c7c5b5014427ca01b838737d6452d3392e6bb40c7b41514fbdd52c1f44136da26c23cfe6d63f4cd1e6d8a6fbb28cffc62788c738c82dad33e0b1e2155d24dac55f18546ef3e954cc6d9cc13bbd7429de3a09b84480eaf6f777e750ecb1c5ba615239b35ef4af1a89c93a7138768;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3cbac0f9d30c1dea78e5ec66c2173be76603cd98667239c0505ad68bb2498831ca4ee06ea85e29d9bc3f4a457fa861acf9b6d1f384af288ff3df3a3fb335810a13de5276505e0f886cca16eedf6178d6f9ae6e1ae6cdf3a362621739f3497a0f6530db5113f161dae663c918b951bf40af59c2f10b35b1d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1daf62bd7b139a135f8da2a064bb9a9cf9d0dfb3d4ceaf243e808b7c41ae1c669241782ff2f30e9ffcd35167b34dc39cde1a3b7a9b27346df1aac0f82898002fc0d8235201df67eab43f0e3681e9347600e6e9aee51f3ac64d27e4500a7b386729eb1b25fcf7fcac83c2483f88666616a7bf15c6c6162b0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2b0756fbcb740a37ab4a870a40d37987b19df8bc1d9565267e03a16961ad4b4d5ce442bf81722a30cb92b75a7a4ea44e5c96288b021ae4aac75810bd40838e6f3e5040c331f36f56fcd02201bdf082abead2f6849c5319ac1b72007372b2e1d87f338f68dacc1b1a47ec009a4e2776fbfb563ab61c425e0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee61689c08f342bab24eec14f45bd9aa2dfac9d6aeaf98da5c9e59f458412d20518b04cd9bd4d0b087292c2dec0f1f25d331dc51a2d24764b789dc818f9fcea8cc61fbb8d6a3ab039570a7738a739946940cb0967036c1acfc04a37870de3dbd6e2c96a41dd03abb86e41cfce70bfa04e525ea1c09f2cb0f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h105cb2ed725d2637ff1e4a69bb640a6837d6da5070f361b3782b00fd9ded8f03b0ed891e7def4bf15a6f48b37139eca448d1150a98604046cd30c9f3c58da855d3e8c4f8373cad6c690fb92e5de5d5788baf2da73673a81eb6b17543341bd82b977ce1519f40221c2c59e6cb3849e219081e739e089bc4e2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a1f5c3b4c5a4b3f4aff9f785f83a9f0d2d7354cea3c733bbc740267930e25cf4614b1d27386f198357a9422e0c09ae8423af0202da85ef8b2e2e1e9c6ce97df39f4898a3e81c24aff71f4735cf87d12afbb4b1eace8db00cf3a1ad9b86b6e0f498f2852b8d5127c502e31e178b76ed0f054add9261423549;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h94e53c5ece224e08364aa74538324d36e94265d7b3619d535b0868bfdbea5f08411a6c1776667837fc351759c47576a8bd5265222b517b2732724f50bf41f50631738579891e348e0b226375d04b728aa25aff7eed8cf09af4e9163fa1302b2b99fceb97a28776f96e2ab87993ccc11d852a79aa503069a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a36dd08bba3774fcb38fadda24ff719a1039e80afed5b9599f6b62cf256fe8751fdafb1afd43b4f3cdf15d8ce7efab0de13a4b7d519680ddb0266f41593a271b8374eb6526c607237d35ed1ddfe13327e4b06328e39880a15b05926569bae720d8f3de88a850bd2ca2aed136a871f0d6261403eca49dcc79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15ef934ecfad871344b1d9e651a6e0576eaff3318354181ec9d03a183c3f43d25c8a3e5934a20eb3165e4b1b7404a5b7c391e77c51e071c965ed5846829b19e898d405377e134298ba383b3105c1c96edf98100de5d92b1a15f3151a7a2a87d3657722126a00aa4a531f06eff5584f442b55ba2674a742ef6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63deb7741f9f3243036ac72f9c33cb6a891db30677a31e5d152b6db35f4ccea17b9c2cfdeaf092692719e956a83a45f3c1c1f018bc1ddfde8b53a719735d72bd2a85f41741cb2382ba6526f8bab10c775df2c85efbc5daf9fd5a3217e358b7a6b8c86ecf710ff590c3d8ac39f82e93e03b1d6d427b59e007;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16309286b4939a5e303a419b22a0eb780958e76fd0e2a8b406e43dee376cfcfa21c2366da5f33efb44eec33911d2aa0579db9bf7e0c93e274024467d089ec98701498540df3430b609eba2ddf3b9a55ca5ec5e148a75c030ef205e06af51f7238bda919690db11e9dc3df2c8682d60b36067c5571a7c352e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a32ff38caaf633ef3c2fbdc1a2ad752a3b0e7bde1cdb73038ada0eb90dcdb64c9ce289d90f9fce131ebb570b7622e1c577687d86c8f159120b9d9706197956db8be799a3aacb739aca61a0a610da3c632fd2bf3d8f9ee6afacaa7e8f2d46daef90804f74b4d7021de1fb8107fca2d77fc126a4d7eb592540;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h150d9fda24c7a8a1052327756d35c56e5cad34e8c1bb13dda2c40ee3e0be76707b6b4120caeed98bb0f0dda85314056b05d9a750d67136acb452fe649d06104d87544b19370c1fd52e73c5ae78eeb1507da444e34d5fd270d73b17b830c0dbacd9e48a8ae59def7ccb7943d5e9d57d6e3cfe2bfcf5f37744f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ef57557b19d9a3f21b987bb5161b8a97a2eaa1b7dac4ce5d12449d9d91fcb7c6ae5fe308bd3eef441012506272011a65ba1fefadb391be49729708ad83aab026cc30aabfcb74f90e7f233282d0a83657f69b7f9e256e7e7daf85b6cb268d853cbb1c1223e7aea43153e9559634b53fab6793fa98b0ac1b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e68efbed9c774a7191f9cece6bd094345e6dbff35b81224236e07bee56f376671d7a52bbf20c8306d9d74282a716b9fc7c7e002a84131997fcd2ef56b408c7420087ee90927203646860ae3df6262d22be2be79b07979ddec7417d22b8905a72b79a00321210da159606993a32737941a2488a466363c720;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6771dfa6a19a90488e7574a59cf3d8819e8ed75f189fa24737422b46c4d44eff9763f93d8868dafd8a501b890365793f6161845d54304b46c984a96fb179f87c11d0a5f42d0a1021d04770ab9003d900e4867553bb4d12ee69e18d3273e61ed2c0496be09230c693e1ce108b791caf3b4f4ae81552d2b72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1227c0723f40948c5d4d511bda9857a3e10f161456fb89b6f5ab4461cd9a047d4efcf8ed0b8458b4b67735dd330e995a7e60cfbe46d6d3d490fe815cc47c59d159b0a3379284066297d342a3730a24cf49624c903d3c929e8db02e539efdfe5738d58b162cb3ae631cca8dfc29126ff49f73dab07ae5d7376;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aaabc036a96c834c7a944b49feec4bb0abae257180ce8ef09ea3357789e8ce70accaa48a1c62601b80d48e053ab83f55f6fe681e71deca095b6394f4da8bd38363bbf7c17ff090d49ef46f8985ba03618e38b2de5fcebf255fbe187d8db6faa2b309064e36cbd8cca0c97ed553618a4b428c735b6acffaa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19483c0ca2886daa7c089616f5ad617357b2876eed64c9900d33610b9ca3d454f14e9f1d2eecef4ef7627e8caa92c1b965bffb4d93be63a44ed1308a20535e93011ed501224cc2725bedd26eb95486cef87a79d3d0b4a11f48205bbeabb3a3e9f96a2083148eb3c794361d0cf53b114c13d8d49bcd1cc1508;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c063d425f51a7f3e1a7ef3957ccebef6bd36c5b54388e38e567f7f10f442108024cbb187087cc826cb74780345f018740016fad46b0bc94abb6614cf8d7ea26100fe28752d97ed6a27418a691c98ce40a29ef5ac1b808eeec6c36af9e5c3540c70654856e8727447e4f7d9218d34e0138999141635346d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haee097531f815a3bbc10de16358b7c31b47eb910cf205c2e16508423cac8ccd74cf279ac0ffdc364487a720004c21cb3bdd7760db0869570df8d8f9849c655ec434f5e91c4e37a1a8f2b3fe9c54dbe1588a5b2d3a3f2cbd2f0c4cda266ef2902db53faece09e417961eb9d52125c5a9568ec42cd97a3594b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h892376e66b6c51316ed51f3a0b21fbbc9488cf4eef29793bd65b99b010c5601da6fa4fd066ba7d4e1028865b78865807901dcdf574d3f6436b4f284b1f1fba668e37949c782ecdc1398da7387b736645121fdbc1eb3408bc3e1aac53921e8f80c7a3ca807e7ab82d903f23ea93c746151b7121574f3c4d63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13267263ff3fe824a9b8711c70a43ab95b661e9bd37ffbfbd58f86b972f73ec16114a9601d44b6c2b98495bd591e58a1758eb4e6595949dac0dd4f1a2fdd6ef021ad5fb3ea4c426a6863c09f3fd2ac2ae48724e31df7f785165a2fc0556655f47b2a3bf4a720b6160eb6eb207ebef97ba04da9fbd6426185f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae3dd1c216ed4f8033721e9c09c7fdbc82325b2ac6aca8c60eece70e3506345a2c8864fa15d745771094d7f75d4529be51b92dc09eb56b31d766a682ce584544ab75689f9d3e6e52b9eaa95a937500a81504c6d0567f3a7a7eb090c250f24014bf2a8d98a5b8762f8d58e06c1a2f0f119fbd2d85aa0bdcc8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f296ca6608e9f0bf6a026f9e2ec21f1dad1039b0b55ce13dda7bc3fa9582614e7ec19a64b5fdde7580f28b707cba21262793b6a4301f7828896ec16dc274d160a1cadc3fc05ab0f9666e87adff624eb815797f3753a77f35c82e5ab92da766a6ab928ff4a11aa5568a8c6900183d34d637e961da552ac72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f09b4791bb533a7ced554001faa82a6fec236641b2b5908b5aac5576d290e1dc97b92a48bfe25c1e70d3e1c5318501f7864730ce795bb4750f325740be0948979b4e3bbeaf34a251c7a14c50b0aa05dfa73769531d892967ff1c33f6f0d4b1f22b56a218f9c7f7731ba9e6fed9b338dbd16d543449c777a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h162695174ebf24a79e372c4a7a09148d5d9eed5c7ea635b187b2001b8553128bd061e10d7a9a8f678d6b2a85e07508a2e00f5e9477f2575e9d229ddfeb2c9e84e00164ea7a31026e26df28e7feaff805054aeab3ffbd658c2d5561e47d3163720d6e33ef7cb2dff935d96820f433288867660213f12bb8f7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf008b57d054ef455092f4fbc20c91e81b3593c1ce33322e4369b9d28c005708ca3e82990df37a71c6a5433e0f676728f82ed13de57a7969ca8e0a42e5ffce1f976ddde3746cfcf84d224e58d0211f62d2a64563ffc742410ec6fd2829918734c376339697e03c9e4a2f549fc28853c616746371899e13db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcebe2d17a8aae9c8dfd6fe0c0b9afa14ece8166e63d87f73149ae4bc9a6fee3d6df75f5add534f1cc0b77af6af59a83205f837ff2e9a0cb1d9722c97e58e635dec372cb518b5dd646ef2a8e85f922e091e76c1aeee0bc1e68a264d255c71a1ef329c20b832f38fafff67f9ef9ce55b8952c4f222d072a729;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e66251b1c1f52f61d46e259e433c5f674cca264053665ba2f20c04a854b4b14af40ddd24e938b8b2611bbaa78c92172d7cb2ec0559570a45b15a9663519e1a1292eb8ab678bcb0ecf95fd69cafea841c30cba1a0e1dfab8a7ce3e2dcda449e1afd9ea243451042ee6a44f91fafe05009929da14d24bae01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c850583d1d15a2b854da8d69008fa23f02d9bd616faa05146c5a86434d7f02c305e1a75bdd4d3a18d40717c29c310f3d3879d4e8561f7e398c57daa59c9a1fe9c7870a198ff3af49d667f6899969423d1bc470ff9e33076953782dd1b8528ca236ed853f09374dfd60955e02ed48ddcc26ddb64faaa6f83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed94af1905382cbefe409051b0e11cb8da749a8c916346006bb5c3491744434b0f25a9ba49f2d2778d875d47e08e3493c02ca70d982b19f248ffc9dd3b494faefba494a5373f632a08d3ea906d207b9aee90e081cf7e902d56f5d95e18b0a58ae9ed750b8b6005d696d727ed078cfe62d745df1b2410736d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4151ce88346da89fe6c9a6fca97f8526be5226abb23edabce681ae4c82094108033bebb2c2985e5833c34523d9c5c0d899c5b5907e160620e3481f6dd1cdadd960e974b3e561249ae32a3003db663c046e6a42e5a1e492212dcf5dfdfbf4a3b34f777f7a2929263f440972501ff29b0065d944aa9e0d8ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h882b88c8e0b3aeffa36938b724dc7da214246f40a6f6cc93001feb14402c1388b2bef73d6a86b669630d5ca2d41a3d7791da6f90cdb16fa52dbd6c59ae65565a733f7e39413333339621ae066d4d56d6c7396f1e69c95482139f51d55bf322565c7523708c392655279cf3898a335210556482a57c2960b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf8e2174214dc775d4e1b347a30e0f1bc7d9ea896f29817073f32cc87561857a5ab316a3d78a533b0d18b378b2b995a4bd637b1a26282a65da7cb7df12703d206a252e59383406c884ff3c7f8fa55d4d0ee1c67173517766ef7c137e1c6012cdc98d23a8348c7e59ac1cbbf20759e9918b99e0bd632caa910;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132d157bcf9ed581dacee3d88af3608d80b4de0fa89a0b62237cccce5343f6a1eb6be23798ba57bfa454b929448d7037b84b5410c944435cfb756ffa5e04d67b49a6591a9fe80b2b46b4fa0a68bb729f2e030b91bbf24388d79732f85cffc8f7182c39d376a89a6e4ca3e2e507c0962c4a5b1e7cc8ad31afa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc58683ee3b2ce3b953ead2423573a5f72e9ccd86d0915d4c5896af25f11ece4317b4ab21476cccf38d99915247792eeeb90e8e903059d6b6bb31d0757001e52b5043feff56789a8109ef2a39fda06bbb06cf0540077be5ada139d53fae6e654f80a070e404be5fdae26fb202d6e2c9ca41389fa994d4b016;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1f79fac79e3520b9fa673068e831bacc0e273ca0b80858edb67441e17cf7bd25a922e94df5175acb1031889d5ab32b235a8d805c0e822b7f08efb4e08c6dfdb737f573a6bf111c08db01806e6a7cd02405ab706abc35f7d3269ed03f35d13aaaa95dfbfe6962ae809594979420a39b41a241d0ef21fe7a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h228a8b71fff7f036e426629094e16bf3afc69d7c1bf117792ef3bd5a713d57bc6d7daff140bd5220357b4ca06dab8e726d4918aec11d35b003737b75ec2ae9f58b94aba1df5150f5b105a587a31a47e19a86ceadc5b7cae721ce408f7563481aa1b58601d5c8fcfe0a8e894b94fab74de5d8736bbeee8301;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47c654805c93e68b09ed67eb5ea984dbf1c5149598d6ce6c8be1d2cdb90905286d61f2c68c2e351408aaee29c8f5b11ab5a4c261d1eb6cb058d8e52275abf1d372f79ea88ea486ac27f1330ee175ea226ef18004f43ba1a45f53dfc08e5d8146205e68906e7c9de11c7c8696e14319e5fb4c1a6eba7ea49c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16cf7f0b7a508b6b8ca7e66205d932ddf9184af28f981e71d02043b79c2aa17bde4783ae570067864e60da6012939376ae0717e74c8da2f368aefbadc361ebcff3b71aaa2cf9731a866e34121a5f10851e85a4fc5d902149acb058a8d08e64f4fe9833ae7ca745ea8bc95809ccaa69772a7f6c77893bd8ca6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d9ad1ab040a7d988c4c240b694701f59c52c137813b52b6bc7069d7074aea29765a8d26cdeba9e0cbc88503e528c09c7cb6178a10567854b3d0e1dc3dfd886983923a821835b5a65b19a85abe6ce46ea88ccfd49b195db1c22835fe2a3b4ac8d78156090d733546e473d5325097157724be326b8d5b3b82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e2578109db0a61ae58b32738385bbc67ddc979fb5b6367f8705f40716d7fbd61ebbb145ca308e792f219e0cd2dfa837339c57b87683818baf08407dd034f251467b121259c45ef7b21eb1873d8fb6c1c808fcb9c6b961ed6acfb47aa7bbec8b3b8ad6fed68435c03f9949565800431601aa284fa5380b75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1233bf170e4380b1718f375a594cca5165ebd6bcb2bce31f52e8dc222fbde3a0cd3fc9761a6654cbda6252279a19d93d5a9e04a73f305f8ec4006c51630bdcdb880e57a719299b207a1b34f08cfce61f879fb49491b1752ac3b8dc5de30de18bd5bc8c4378095737b098a80781b889e9d1bf7d50dcaaa5d3c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ba9c71b716107f62c4aa822c09021d1b3ec88e31ce2fc538637a8661917ac4e43675b1ea27b5eb7d2657b6c85ca156c9c9bfd7f6f5d052bac5de537a9f6c945778376365162ffaf0a6f95fdafb7541335b815a41184df1ec7ea67dbb9a6d8e3f7f5b611fc72c376514d500f08da5e0b09d21eb9dcd7e963;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151c961b3722124c86364b0ef703b9047d999ef004d87ab509ba0e4f25d865a158770413d2e68a38dfe2f2135b081f0e1ea456cfc480306c456582c27f53ff53dfc087739e6140736f2a39c1c2fa645b9f73e13853de5e97e0944d0daf7c7e99f2882d156f16a2240f063f29477caad4d9eb714386d7c9bed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116411f296a76461cb82335cda35929880c7219c876ba7c89e81a3f4c8669bd5744febaa980a3c3366a4493d4b9d132408a01d146270ed8677ea622d7bbe5a76df2df16dc24935b275bf18766299cf463fa82906d0ed4b1de97c002472d2f20b9f0231e641f36f920b2d57450deaae9b71565c7af8ce5ff6b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63529619848a9435b6debc74a8a8cf8479297153c7dbc910ed1801969c3e8ba9e14bc63b215bf0040e816515b4d2d7ec76a9532da59b83c794e6ea156560c918a0bf07498be80403f437d6f7088e575c90eea6e16e7e3f2ae116f8c20b62dfd37dfdf8af8cebd887957e24b068396861b90e11d9e68a7580;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163fe4e23a7601ea8f53c2747f7e33435ec093a24a8d601837f22b11a72d10e15cc612a7c406dc69ba91150d8a861a0071995eb303d1965d355678db74b243fd66119190dee5b0f8fd4348d64e3dc3fc18b1a5041cfb3f84ea01e1c0834a0badb97443e46bf2228789cbe1b991b9bbab3900bc13d9f1e7780;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12db03f2b1f594202bc2c2ef1f68f51ca360464bf9794d152f3eff73e51b0ec89162b94e49e4ad3294a5fe1c32c31fb3e689252fe2f3a8c7a1d720983cd030612d995909a34faa82af1314ecbc6ba0a70e4c1074209a5f1e44793bbe3354b1da8c0e28fcfa8cade6e78889fa422a225f47a416c6e80ec3dd7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c5edcf44be62aaa029f2ebb10b9c830eed734de1d655d607551108bf7f47c7d9a1544697e8a6a7f7c1c476594b1f926730330b49034be066bbddef554425d0c9d8ed6617084cd22f52a08be5c20ccb0efccc7b943df47ae8279f6fd4436e8ba42c764b2b7a630dc661e4217676d238aa9a5398ed983ff71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e52bddc61c32307d0e9fa6b688aa6e4e5f3031ff5bdd7be98ebc55a15df0ba2b8efa8d5c4dfe136540d0de29bab448cb1060de90982fbb6e643bebbf3d2278b266fd93acba979f2b0f584810aa0873cd8bf07b80fb7ede20712893efbb53619e72ec2b20afb59475e66ff24a402397710f633a88e7fff75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de44054274f4ca5bb73cdaad3dc4180e2a95d052937ccc917d327672e17a86637dca85be7cf6de35d0d09bfcf1ca386f2728fef9f5a4762892b3f7a523279f05673dd7ecb98550f540c4dbc1c1a101ea13dc31320e643359e3c72049a8a6a2f4d8f55fc1b8cfd86088365fbadd0d6ca41f2e86aef1914ed3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd775931c48940011266d31bff5bf4e6281b3a04c9f349a5f0b84e594fe8831b2e2cf3082049c2d0422e23019bff974fcfd69d7aa9d96c5c237ee5f011b6be87f09a3c5e8289eed5fb1e6e970c0f280b2b5c81bd30c76457d584ce0531b446618c32efaf8a5b75004d3898abfd39a27ff3d9b101edd8de498;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa797a7cb1bfc7c62709063a90655942bfd2a57e62ceb344c154bb95bd571fa68fc7f66018d18bc17dbc4501710e245abe7e8d227f397338a2dbd3053f48c1dbb70a61b92878345c432d12b14fdeef4fa4f3119ddcfa69a2f918fc3bb1f894d6977f0ae1be1c92f4fd2bb4cbd88c3eeef8f6454904d772f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h247d8104737468bfd17fb6e4a9fe8ba7c8d69de649b8671e5672e492e3e14c139fc079122c83ca3e86ac1f3be5e9aedb781b5cf28281ba783e26b0ad46352f1ea5c7a49698086f945b30c0f86920c4421bd0c906112e9bf3c8e319713615bf6a3c77699d58ea59359fc69df45e8c61e05a5c55269f77a02a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f21ff94805c1dc81ca92e2028be5eaed74a529f00ff9d99427c0ca4d9998218a6dd1643a57ed8281b8f1f900ee53c244a4d3464f6ab29f6097a4edfbf59cbc512f282fc718a1f9b8f94de56357728461ffcc10d762b30c4f107258967f82f8802e7b3e93b473358537828f09ca73f4fe8f8d30a23d71cfb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h504ddad6d6d90ece55140ded433297e65f25ebc034741ec1b97f4d5d4676543a9c23c9687dd93d8eb1e774f38a74346506bada1e370e65d710dd08d4fae46fc3a45371289558e4a36a00d73b71e0734f4ad5975e90c2f991fa84911d5474bf43d356fb521f1a072a57c0753383693aa588f31946407dbca6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142a24dcc15ca34b2557f0c52ab4ef66a8dbf2a625b01aa6d004d6a21fdc5a3a156c92de6fddb9a086f604001abe93e5a794306374b1948392c901a2a5e54a827c7485bf8ac25bcaec57010c843c5a3eac2b0eb1769cf48aa98f077f25383ef121924edf5d1973a10b31c258f5100c1b3d2051a1c14ec425b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11469071f58a0b9804de29ac2dcacb4e179bdef9875fdbc933a07cf8136c567adb39540be6509b5d3e7fae17080e7f7a0eae55498beb654a14ac9041b77523a8e77f4b9d25227401548b00f7039f61ca3cc3eabfc5dbb1f94c4cbb695cd2b3a5d42f0a5e977fe4b1068419717f3a13586188a1791a95cac1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138435dcd6feebf86d32754bd0ce297eabc82704187be691b749512d5109ef9fed9d10abb8e42b433f1773364cd4dfdeafda1bf313ac54c22c9c019a3d31724cdbddf24514712fd4bec434a8745e1f1c8f453e70dba108d51fcf507d7a6c0ef0dcba73d02b087861171625145dc8c020db73821bce33fc3c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed6010c5a08773f13d10dbd1ec6a0ac86d532d3119dd765fa54bcc4c631dda24519dc50cb7f172a02909fd82b2d8e41d7d17f7c80e36ea1d46b06c55da59aa9f5f76d20b4c949d1778ffe73448202f8c79d77f9cf784994e9e64a1226f6db299b2e5e68f286f3b0187fde3503c95e73b46a97f2c762c5ed5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1797fd3ac490e9e74ac378421ea2830c4f48728da3c853b1f7865dfa378875c2b4728c25bf1f19972de1df53da3af61e155ab5cb2a373e98453a38854946110700055b57001a5c41d08a497ec55357c12bc17944357c8a92036513ecef1feac0811f2c88c01f9521919b283bd4c7e0b7fa00e56ef9261f41e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186bf6e322a77fbabd04c3d83a315bdd96be2f50e51be3dbf5715adeb08dc1d9c243ed57611afd1f37ed8a72677bdd079b7fd29ce52438d47ffe9902626cbb20241154ebe3441d473fa7546705510eb9b22c0c3cc767313f2a40682a96fc1a3d6d14c95dc257064db7ba59e042615432e266cc841bb51b095;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58515e488a4b9db5546c9a78cd3ead6c759284518faa33226bf23c291f320489d13d785e6ecc1c5677f82ff58bf9cc922d1921e868eee72c5e816fded6c88faf061a8f6881daf0b00bdae1984153d56c11fa147a0f97fac4f4a7466346bf9f0f0dfd4aea3d2c3e3bf23ef1d33b0c8edddeff2a47775e29c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb74a90fe91f8cbcfa521b563707ca20ed9039ed7f30af9a3641b7801a17de54fef26339db45c6b2e37b140896954aaa500211bbc2f939b5f6225164b26ab601188209e44471c1db35309f10d8d8e70645b136e00b737b8dfbb0f7c701bc0be4b562f5f3f6fc43790c5305bbc47467ed9855856d8c55d153e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e976441e704f13da733e031f1f306d5d17fe039011b186d4fc5c2c024e9d931303ce7ff478e441ba2eb5dfe9c72202ab0e2ef270f8146c17d487f2e84d1012a6d371fe991dac9f09eac7643413101d8770e6aed5af2896d49cfdc45a6eb4e77f6b1c4cd6eeb089db5034853ba9783f65a4a8ef4cd52b059;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba2578752e14b19ca88146e5010fba310cc31a8fde2efa74e44cf3f491e09fc8dccaeccf295d76004d48cc8192a76c1ba86fa15c1fc4abe52032805f9131c9c5b64a66e83a1cbbe27ea1b3fdb01d9c89367ad710b4bc0f23c9255c7bc714aa00b6ef7afd278800a21c6937da9966c682aebb70e77d10a37c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113517756c5edb455f67b43938c783991006ff4f4ad688ea02075318831ba498bcf09464cebb6aedd1018a9b85f341fedbf7726a6005a38513e49c0f5dbfa1f27c0c2e7e2bf325dad31ad4ea8c6bf2cfaab9f5d424ec449ae6d3103748c515cc2082717cad1f82be21b78f4217122f1a6f22e4eb1c402c75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ec768ea0aee78be87c0501b58c6eb207cd3b6bbdd65b3f10f265d0b2abe0bde565b69046dfc7818463a05366f76cf1570506cc9099151d8dbb2f2b8ba63bce2efa372fd4a9889eee7615f9ea99b59830d56d30622079a474a611ad71ee5e9989d70913365aaf5e4b99d996033cf53b8c28d9f64c5d1bcad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa6518a16744742c04bccf9759e26cf88fbb63ce957f99ff3df804e5845ddd7c95334d1765e3b270c7b6356cceaf225dbac6390594e680611a2a9dd3ceafa6fe8baeaa05128d3cb0aa661d85655250f3a93d539173357884d15f6ce027756132be733a4948423108bf74aa278529b69708b2cc284620b9fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d8994d8749ff7e75006fa1b5a0bd8d0d8e447db7d00b7f505a5b0bd7007f7cdf797fd257d928fa51fe7cdbf4f4d862a0ea45696936aa874ee5cf2014882526c43425fd2eda2e64e0f38031088f104d0888e3726c3929b9bb360ed600a03f6a38e593df93d484df746507d905ae433072d7461e3b7bf0f94;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a75778e26c471c8fdbe9d531daeb732c2ca09a9cd465cf1fbca9fd48891c670ba29a7e77691c9630d4790a065b6b6912d1dc18291644306bb984de447bec3647dcafe1c9820ee5ab8fa0eea54be756d7ee5d3520d80ea4d2717422e07df78871012db8d544859f1b7d16a524fb0023d9f6c10b06120a1842;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b46d15c6d3d96ae04e422206acf5cace583422f5df0df45ff562722e7a0a11eae16572579d884e2efdf5f99e65509fcd2f920670f9376ba7abbeaecc5be53ee11fa20e48c9afc05ebc810d3067bb4a14f9d7232ecb062a464c7c46cca949582cf9fe40bf48f49ba84afb0e9b4bc781771941b34fc5c33a20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee83445677ef00ea0f4672a5ef4c53ade288ebf78e2392b640e3c76c850f51ed118aa9edd456e03da2000ed36fcf9d12bad628ad95a1832de6240d177d5ae8121e5ec4b055f87f88081d4e0491f8f34b546fc327e60786f989722a9b98201506f32821d8cfa35276058e6da77bb15f93547c56e1e2b53f9d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h602ab20602b2599e138b8c69928a9580aa90124441f43139ad5b7e010d75f89ecbcb64ed70735c7d610a096cdb285c6c52ce6ac8624af185089478b15b641d5e5724972bfe5e509936362093b01ada5d0520e04179e701bf507bffb776eb0e8f2a5afb9dce70e56ea2c2c870452445d41039b657736b794e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h161b015e542a2914e1fbb4a4335849cb004354ab43d1ddd83d5cec5aac2335a49a0bb87d3986d26216bb4262fe93cedbe5ff9652fcdc4d22f7713886efb4da6c8f1b055bfaad848984fe0567cf67b14781a6334269ecc146eeca0adf47638c106346f3e2d0a193480ca5fc0646cfa8452038477b8e104b0ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8df6950ad30b8e4c745674ccb0f4844c57f0c15846c49c89a27beb3389214d24f4c36bdeb9b23be0de91de4723c2b1caf39ef63415e9a264f56474c10f3c6da67cc025061da17262b1e163c7cb4c75c229324a660d0c59d67c9c9857b0abe6053ffb46b868db20ed55090add8e7addf992a0996b66e97d3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfade547f3f7f8ed4e4d277036a0ee6e8f59ea76c6001e20409613298160ecbe9b06cd92ae4ff9992940199afb8967b8ca568f46207624c42f02d068ac22e3918fbfb2d09ebac0edea2f55c7b0f8a59c1d99c85d01619b318da00a9241a3202f2821c2ef36bc8a2f1900d9e46f9aa37b47fc372a634c7211a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcaccddf32cac486a086d76b53bb9c3591e154df0e69944a24e4ac1c0b878b07e7452bfb849e432a0baa97d452255e3a73b72067d1716e242195f6e0297729bca3a8d451e003372609bc3f46929b7033ec6834c560198cf95ebc92dd3884a5dd6e830688c6362577b64f6593f183e499a7947b4662015b8a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96000f65ad30c1ce3348f5f2d09622b4ba7b0df24ce2ec6694d12de5b3f8cc3c3c80b0f175d988288e949018f2d56ac57ebd261a238a1e0353e04e51342b74bea43fb80e56a8c87d6416f624383de56778a793e678122d4d600e86583e9ae00470884443a36d1c00224c422059a3f4638288c46464de69ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11dfaaaad9514ab465787cd7fe2ca3e49f546095c5ad83eeec4c49a0a7abe483359e5fc7d7b34bae2245d35bd4b681e761189faac51ac000dcdcf875d0539a8890e523bbe7f06c892fd7be5473ff6da6faf9acbe25a93e32c4dd4927824be407ad00cc05e25cdcf0730573989bf5f9e5be325f5d348649466;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2a067fe5bc858af7557ef3b84e500b4345d28ded5b278d42cf9bfc2c894d1da932d8f5f4d057d1612b68e0f3d8ca8e38cc4b44ba292fc47c7e4ca2046ac6cc52851e80ca3bd591bc16ece2ffce7e857b1840bdfcca10fdef6db22eb99f958ce03905d957622a3f9abaa38b36ca1f9667600636ae2d8f199;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h123c13eb6f202c67e9baed96793c3370cbeace158b5008eb27a0de7b228773ff645dced4f4342b0feccc1c8a90ff60baa2d0f4272e6181c0251b2b1031d2eaaf916cf19b35fb68bc7b263cb03680f9dc42504b2da4e64e80fa16f5359b65ad10f42d26036c14c76edd298e6de3c3201be39346c54d76de752;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f8243698609d6d43e2f1c59f6ef635ca22daf649317ce8dc6bb3f75128eff5a53b77418470517effc5bdbb124f6c8d7935fe2257dda9421b08cfc5cb681a5ce2ad0d1ad22b5227cf7e448e9e274238e8001acf54cf8db2ff035c78ca024817909725befb934adc8f5b67772e1ec7cbf4db23ca55e79f7dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf6ab4d74ee3c056358bb0ad84c597aef6505b4070cd62e6338db0b6e29fe0724c60a2184d58c66453e28512c8835b0e390bf4adb310e28d9841f2727e4d8961fe64dadf0af7c6482e04292adadec80a40f56bc1217a9ebf8e5e1e0bac20174deb76ff6da9544f581ffcfda29702a902c0612aa0e5b0d23b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h120188493eb85798019ad82761d5564a746e0f7200c80e02bbb109b01786b99e3ee08064cfbc99758a0696d3bb1c36460b23caa73b04d4e0581af1a05d6e7d7fe5393783a29fae0cf222729089994bdc8cb30766d0237df7fc334813d02d0d6e04d5c5b364efbc711e6bbbda84a9e6d7a507fd4a37313d97b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102f7e1d591016c5fecb8159d70cccaffe9b2ff6588957e4a8467951aaddaf75b9136b2b89ac2680f0b438a0f64626860afd5ffe7eb27022ff91fd46fc4fb154876b514fa029212364af5867310116363a81fd963454d99417a708bfed95e113272658c695dc4dbd65c616d02de10abc9e8396dda874fbc58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa6b0009bba0a9dac0b526cd4ab1d79b12353af7b5121d865bd618da044636c1c3c7a4dcc49b14a24136b8de0495c632b4ab4e83b0ecf896c6ac07240ee58f5787b226d84f0e4c599174ff3f115c06f1dcb457712e6bbb5e0460bd46ae9225eb8f31317026fcf65f418552e4db16dc59f59b5fe8fbed077;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e8a3484e29001488529e98350ff8bb24d0642f6ab5e45f9401fca49988fca1319ce1e54f28f730eaccc0d497d9a02ffa21054f41c3a557fba2ce9fdc48236f0655fbd8000d9552a630de378a8877a4f12344e1a2b3d320383aee3eaa3cb84457edfab211686cfa619e661ed1d46f6fb26d4d0dafa484bd6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e1e90e66eb9f96a20974f7fb105bf584867529b24531846c23e251c6a535e50ee0b7a00d1238dde15812425aea23eada600f6c90eafc958a0ad070a3934f90599bf1db33db204f30c976851658fade0cf89a6b268caf1a844369aced3b45cc3ea96245ad533d8f8a8261580ebdd7bd9ae8e9c7b0c4054a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d16d0fb1871c95b2bd9725b76809be95c53938d5470d82c9eb2b065a9dd7aacf04c68bfd99f6a4acb2fcab071a97adcbe77c804364976c5e0011a6b1fa24b66ed924f201d50543cea8dd41bf46508186957e9274eed218dffe8ef09c9ed34495b06b13a5ef63f1d4960b7bdab4dd41367e678465ae5f8679;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb1b0573fe6bd5aca0fc7dcf95affc61fafcf5b8ea0f3d5c71b14a27a4fca04030f5c93918ec58a8ce5ef40ee492c928ba694013e69fd04b77826cb35e383b6a336d76a4d24e54299e5d65291d6f1b50c2e7d907cfeb8bfe8b1f496b96b6c5cfd6c8dbd6154d2b726d9ffaa1f474bc45fca6a4343a03c6d50;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4f5d51fcc4587b2812b7d0934ea4c75b3c7a3e312032d8787fc9b83b2559785815e56ba8589ebfa7cb80d23703d48e393530c84482bd135f4a9548755b40c672f25e48c45364f996d06f2c421194b828dc2010dac230a97fa9ba24c8130e54ba41f363cc15bee2b91bba8c8e6569389a279238f0450e0797;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70df7a71a6d85a2a213dfca92c672d2dac7ddc48356ff55f0cb6bdb59b798ef6c25ebfa8b78413bfc45a01a2c00aa6a28ed4a20ecb6a2a7b769f303fe667945ddc053857d391e15bae761a4e34dbd10905b0ed303831bd9c2dae200c4866d48fd7e50392d2d0f64827058db0956893e7c6e1efbc1fc6f6c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h740d8af507fd8ecd04aeee0f0b838ef772e3c76cd5526f267c7cae5465d93c33e02c4b0ab7ec468136047df356767eb1af82a8dd9c6593b2d7757f43394a482793d5a77c4c455c4c334b2e0be0d70748fb3ecad12dc5784e0b033baeec35f30b3b288225e5e2fa22bc8575e7f862c726a5b19ab6e208605a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha2ee47bfb2e1d5bc53d8ee41ffe9496497a724785de8961e44b3b5774d726300ca097cb48ca839426b924e4ba95d822c8e4f0631f285ad71f0458409d3cda6e121b2561bd5b5574f925a99aa597af298dfea94409f94e80d7d1fa1ebefbcfad8f264355a73b4692a6c99cc4dbe69551ae8224cc85b7af977;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de2983663150dbd8272be55d867c34f5d108ab8b20f4e9191df60999d0d1b5447aa9d546ab65015e0191fa45033bd1765f666dfe4442d4d9e3e6e7a33c697d889ea16a1720ebf7a721bfeacfc82d86e57d357a824556e3860d2f81e08823eb59d06e2f6bbf8beb275f592bc33537e7cddff0e2e0e4e39582;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c222233989d0d97783dc2ac896a5cb181424707a6e6ef261632a62fcd58440d4ae3550e20c7bc3ecda9cf4cb63fe11e38eef90566e1b6ed6d485f5b31ab50bfeb40671214d122bb405187eaa7be76a2a46394e518766af272cc1e99e4388e0529b30ffa6abeb360d97fe5c51fa80981c52e636d08042fc32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ecbe474c7b1834bc89cf450dcbddd494ae3023526de2ac81f8d0e92530e702b3d2512d3ed4644972ac8e0de3811c9d6ddcadaffb39daa6685c4b50d44243dbf87a01f47ad678277f76b60698e66ff7b173bb0c72b333014ec38d21667880865ae929d714070e1c328af0c23368e4e97d39abbd3c36f930b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c51171a7b68ac080ccd4bdd21e1ac09c4ed82a9b12e4c999858ce7b598f2038b368b091032b47660a1c879fc51e35809a81bfd280889d18b6a248af35b5351bb193aeb053de902eec78b3eee14b38d285d0ac73f4a3ad683500fb41049e01b4dd8e24d7e6011ecd1c89e154a28077a6db8bc8c4790286ddc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h729be3ffe732f1946588817adf116eff94b409ca95bc7fb0b2cc855fc6a4290dc82143e9c1cef691340057484e63582012f04702343a1478e643f1149477f8a3e6edcb8447b7bfd2c69e709cc4c66ab6a587d8a92c074b9509e1ba674145454b234762dd71a68803c2915f85d501d9f1143525de80e87935;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1217aa018c06ae82be0d1def3fab9bf5eb025449ee6e0024adc6ae63fa8c5e224c042b4e01ae63fe25bbdc642515007ed21e7bb5d757597c530cfdbaa214971f7c26261a0d91630c379060071be11c605617a1fdaf690d1de1678ba5e348251d560c6e6d5d0b2816149cc456235af0fc2a6df5db6203e5999;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h127e920f1a430e5bcbc61f156de7aaa3e47ac12f3b0217e6f0874561d69a7235608d4b3b279998986aa1cd60ab27e1742feadb41c3680ec7b0a4bec92a85ae330e391c50861eff6bfca8054ccb06ea5a5af85ca127c8da4b6fc0e8ea35ce9fa8920fdd202f174ce2619eff758edeaf415996368c1932a5896;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1093c932671ca23553210654f4d14ac9526181c7496922afd02e188601e4a062679bd5b9ee6c928ab90d7f6343465c13a476867f1f80b6a574407b8185d023c36da305a31152e85913cd61a5affb615434a8ba22235c39f8c41881946e3d0d87630e9882960eb44a09e8790bf8a519e4182d2e3bafd492ecb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h135a5fdfbabb0e00f9ad1532fd1e014d36830aeb3bdf766c090d5dbc03b12f495a50f7e9c6e657e07186d9cfc7145c9ad098f008f002d8ecb7cbfd106c030b3c2342b68d8b56672ea5bcea5def8137189612252acc26392381ed3195345443109446a18e33eccf724a3fac485ddfddb415d61b30513b1ef19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1546731b06ab22f8dbbcef1f1cb39ce824f55fd5e63c0224aec8bbeb6987435b9ec34b1fb70e684a4752a382f333c27483368cf100a41cf3900517fdd9f1cb5646009497a46304aa38d88427623632ac6a1afc5af49394ee2d757a1f3c5a98243263fd3e330ffcedacf7d89d32d906879654a88232c5a5268;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2a08511d08f9a5647e7e93b4ba7ac35f512389520841a48b4fa1dddaaf98a7f24149d85825461b846880abd6c77e10b7feb1192f5c7569f37bb147d232f5bb944e1b34be7fb2a87edf507a1ffb3d62cc5cd5356facd3d7331481145ea602613c37dfc8152300f66f06e3b1bb21997d9d382cafedf799a84;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec2a244c8c1f55795bd2acfa7cced68d4eb61e4f1bdb43595b31821da9b9e0130e201972f8854e08d760d3f7fecfd1a06e2eb4510f9cba999747f84b13e2a6e62484cfb5ca88824261cc82b5c8ff5e1d7a8b736e5e3a3536a7f811ab70f8661aec7f8bf0693e0afc1dc224ee9ecf26e3371758dbf5e7cd34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc589965f6dfa4a7dfc6eddf053a7b9a8d3dea5600f3e26240e2428ca937df733412204d176b9bc7284d4fad20034d5dc6d273d9cd3fe5d81e2df165947f1afdac47db8a3faef2e7e344ae4060d914c2d37deb57dd8df7b2649ed5223c3c08c7db0d5c531642eaa512a22465d610380061ae6f5d4bf6ea8e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115acebff7a5b04fed88a271dd205f6e0a34f2596e8d9998971e69ebdb9508352dcfb9576132bdebca1a59422d9f5b8b29ccc0ea13ce775ed39bc107aa93b887139b85bf7396f15418529467a7cbd8fd356d9b13f58fdb9a12e31b692bae2bcf2fb958c959d194fa76bc5bae335685523779f93eb25ed2367;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h189ac019a09e3f9adb1cf01687880e8c45fbca15a8067ed2e2f69324a47563ac4adcd1c44e0c915f7213f5606e404174a4269e27465cd3e02c07a5a8c518bde1f58e17ba00e0d8f095437654f80b16e001927424a26a3dc5ed28d53eb2db774516cc9e8a0e6f386e00aab1cfbe4dd697cc20928f2383471d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a390e4278305cc118f2259fee1030dbc97a3a3f07d3f6fa5ea075d1dd22f04bddd65599478e3049add349070a36d607a8883766e792005b4c4ef40979de266a0d905f86617a191a29f1b7f3a1865990d66396e7cfd8cd05d134ee5e4c50227f9c3f88366e335de5017231a310091af3882b4353189ec9b7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3b74f3546541885b1c747966573adfffce966d8a077694fde24d3350ee7145562f702375501ed081227db6846cf499b287b0dd951d785003025a94a4ab45d98caac386afbf1d5d45e01b95f21efb5bfd00ad072905e3a9e974a9a09507a73f0f099c3b14322bd5fbf0de86351f7a2c78d8ac8628c376fef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d0a10400866133694dee91a1e9a2dfcf59251dcbb85dea783d407ea21924976ea13908f17793cc6cc8889b68d5528ade2f71fcc4104ce358d3407a81a57aa4d743c487368b4be6a98637791b92619703fd6126aa7e62e41b048d5eb67b959f8bf68434fef94090190d445e89e6835467be0ec72687ff16a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f17a038bb4ddb881c7e0b307040b7e9200214a59ea59505e841114899bf9e2b715ee55c45cd885dcd1500c9c0eba770d2bec2cc6d5ac374f544d2377750f0270a89a611b6dc674272b6ff40cb268d1a3e004df8bd5db29642dc2e5feebe09af45eb95024cf48ef0fa133c0a70965a059767eb75d464a134;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h781fc07048d123e79ca7fd9b1b9e8a2392f71f743f4e9a29fe408d2e3a4dfa9ce73848d6e6ae2776da7dbe979f1d246a4ac3d472796d2a46f47c439289f28094aa111e3aba92a483ba1145560ba48eb14cb22004db90ee63b458f3475b6ac9e66685769a51a09b204410d6935420651403652d167208bd3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5ae5389ccb4b0de236ba46b64daef51d19b64f5220e093a446b9917e27f6a6b98faef4d16234a095bb66d359e7246cf9f9e66bdfb89b9292d6dc992474b3a0d89f703a7e67df17c05ed663eaabd617a5686a23b7f7697aa933e58aa40efed155a080a4e7340eaf4fbadfd94d6efb4fdd0e36c8901a9bd79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67032f522ceb3d82d01ea9b85091ca872682ebdf3a7a389b88f8d0df2f58d45f22eac5f9b2721f9695ee6dc489e5c73c28e1d4eda78579d605e7484b8764e5fc0f1ba13600e05e835df431ae5d333337edf7cff782b60abe779522614b5a7863d06590cf10e096029749d0e9681777c357e7ca4478976fa6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14be1b8e9187fdb277ba90ab411eaf3b82853ee0a07160d3256094da4bd1290c7bdf1174f857f7ad3875f8216a73d054448e65cc0453119fdc50fee9406c4d9a765eab5e4ae5b171e717c40e7cddc3f2ad56d762f3987931fdcdab514f0521711c70774a20d0ce44c3d25d3212e0c71024c591f2009399671;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef857d3cb7effe7d6a32ad906c08f83282018c43fab1f2dca1138bd07003c3bd8a8c9852d465ca21cfead3f2f0ab90db9cf86dbc04f98ace14dca8233f0a3905bdf2835906166aadf56afdeecd74a9d6c359fc74c6f12af3f9f876d4c8b6e95fb3bb651f10042c87b0bf29db857e01a2b3b4b23f6eca7ecc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f689124d6a24d5b82e0cd130486bb2deb85d8b73c70c475bb2bff3b532571b2022e6479e9114a21417a1333e6e68ca9ac4e2f6d9321f7cab8cea202a79a4f8a44f920ace4da870394f82c031f187710a062424f1c83c5da6e632a2ad502e2f235204a1fb943142b888e6b25da2a293999b321b5a4c49390;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ccb50bb969d02cab3cdcb904ab43a5d7a606bfb8b1fdbe2b56ea236b2bd807bd4b5ee6a99b1e33dcb2a4b99e9009b221e75b7d13f9e9cd037168fa7c2e2ac879af0688a2780bba54874bd4c9d5a1ae33b1bca67cb15764c5b77c1a2ae652f627b12052ec16432938fa4f6b6e85baae7c5c68c40efe4fc92f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da197ece0dddc6c3d47064f21bde41133c73424cdb5630b0a2ea4ef3117eec858ccb587abc485c9660baa8a4caca163d6ca9e92529c5c5f16feaa38d86682d9e5eeaf70e99629f588a9616865192b1c09f96587c8f77c24d2b72add555dc9614d83ee6ff36d5bc4d6eda70260e42fee5a28a2791daaf54fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17958c1a6f868b90516b319e68810e377cce3302d131abbf3a826b4ffc40aad8496f5f8d893224986097c3328f3c13eeb567b3c06c97428b3a019e469794d5f7e54d6905aa076cfe7bdceccb40df65e6c49f545f20487d145504b1c05411a7eeb7f8833785f00f4adb3788c51b130534a62cdc0821b9215cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e083b89e8df964d26d81cd76b303d6b9d2c2310c18e24160a23adfe0d760133f6d5b625ee04a44c53c7591541a1555accaf88d9fcd505230b6b5ab6ad38b27de79f8c40ef9846a1038651b30454869aa36ab4aa2fe5027bacc0f5bd5c131d47b397ff3f130322cc103c729a6507ad61f16f4a342cdd738c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f7a1fa0fa066ed0bc01f089bfe5b882efba43c52c63f0eba2274496186b69432e14e8b4df0b2dd14a2c7bb980b224f71e5c30a1a53e3197ff61a6723eb7bc1dd66534db717326dfd9500c8c7a229bea27b78c6dbb981954a5e248d32f293373842df051af0a2f5a0fda206aceda03ec63fed13feba4545e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15a0734dde0b5bb441b906e651ded7cb9d254fad2b07ef583ba10b2462efb7d4b21390bb8194889f49c69a97e38d54d05b7b73f2c988f5470057e54b547c7f39493e87dee7a8fae8e036b310a90d7a3840407204734cc0eb7a188e2168e2d6a3ac0de548469f40932abc1e54a3a05d9c87275e9f271ad38e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a28409f9910e9fba10037a5fd01517175560afdf1cd01d282b16aa41a62256686610ac9b057a2e56f5ef316238ae680972244ab71f01047a13a6807e1661a5d4713362e7ee93128b6c94d49740f800d7d7299ce9415b61073b81bb7902553ece8d340ded8a2bc5fa3d9c7062182753673b993adcff5323f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc82d1db73379c0001c8625be29f7447f35134ef360c63a52314aa1c80c0e0bc87adf0c536a7d3f61cdf65e3e046fa0622ee7e744948269fc64effce91a3072d8b064a5f1766f8d3d6f0ffc7c9393d693c5d438b5e61da57227469fa19851ad9e5cfe8c77c0dd0c7b1f45c3c281cbda6a60ea5647286ece1e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e34b37c5ef90d25fab0cddad32c406a8e3f9f4e8b43c790cb3abab84e7e50d526a7b0fa53747fe73a1e6272cddd41a9a6b820442ba14c0ab5cfb385572fcf85193c277864c074d25a8bcf0f277c1623920e30890f686a6de57ba9f06f0ba1a8172b0da60110a897b6578038dd7726e828b943a9a4e86a0d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e0552769c9951f97603754e1bcf3703707d259d4e27b7b2717c5819c9c9cae5a2fd9df476792b77ae9e2cfebd279151606517e4427a5e4f9f65617a1c2fb8b1f5646a8986ffdf428b800f01f4a16c3d0d549482ae720bc2f681f2a084d4e44e2d627d50313d58ba0555804af8086981a4229e78977d5a22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1763e67842c9dc1672d1b325f330402d3ee685b85a5f51038e901dc1a059526d04a2221f4dcab540f45be6d5e6dac5c130ad62f99498f44589d33393cbad6f8922b7017a1ebe530a3a02c7b58fe7bee33ddfb9954c23dbe9d7693fc09a88c4a9b0a7de235395c938988f06d0f408b0cbc298a88338998cb4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1c660aaaab2983db01eef8b00012d5f44ee833e31e7ec5c3568372ee4b50cc6fa4bc65c701a3ef9122161f9d054bb6a282a96d9e78418709ef8142ba8e55b2f7abd97390fbae26ec7565686ba6f33027f8d5704d6dc5e530d61f924b87d1b49438ca6a570d270751fe2802f280790591e330073abe0a335;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1169983bcfb6bf79ea107fe5ecb156853bbba1ab10e983cf88dd42438512b329898fc372305bcb450db039f6946c835dc11eea4a5bcb2f5ca23f5692253f62553960ee7f27e139178b28e3c68174b42f8ad18f708566fb9054791a98e9485b7f40f93dbb6466685823aa679daa1b05324f5f18399d4e1af9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2f6d9f8fbf6e63d362d1d6cbb18ae728f02a2313f8b9bec67d117140328873547dbf9f21726b23c2518ff67e4a2b00d567650f397551f99c205f7ab3a4981db7b034a17fab4943c61b7cd9b0d221afe26fa0d97c6b6fff5ee0563d941e393cae3cdfecf8ead2594334116fcb23b7f4ec2e42d67bb766ec1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3e7e4f45db7ac04bbf3083012ccb37c946b27acfdd7da136adfc632facd1e83872c0a44c79b24a572123e98d8287f7961038fef8d5f2c50fd0f93f484ebbaa4ea17ed7dc639cbe373191549e70022a73e358c609bf79553aa7a5c99e69cb9a8293ba1e7fa2337b5ca0060da8f2e8358448b8e8d71e0f56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9dd81814a80146db7bef601b79ed60983c1df16ccf0e36540c234171a66dc2a013d28dbe68e6a6d999a8f6061dfad9ac7a83c485b47b8b5bc103c96548c502598716715ca01ce067532c223cef93dc2fa11d8cf9d8fb9dba06c95f1035fa9ce588138cf5849029d21547f2580b7d7fec142a5c742c09a765;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfe8d21772fdf3b4cf4093ce5b26665b0f1d94b0c4747e8eefe55542d1bcc255fa9332c2a1fb7c3956431fd2e331ad144ddc9ef89b860b9a5b8c86be1d4675d27e9575717fd6c339a6ad606408377172603e47edcfdacd39dd61c74131e4eb0d1ca37c636b1047fed76dd1240a1928949abe331d69dc21503;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h395f8d94447639d7ca939e490d38f5e895a53a79b807aef1e6c8ce0fcaab508c60b51c76ca0999ac9cd765ec329b934c4b3e943e53f99a700812420ea85dd397d8252dc476f6edaa37cefe2c8d2f6ef357dae5909395492f71c8ad513e36878652a0009366e9ae92ed269696e16e889bca5915fb06e4d984;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37f3f54334d276326d536324146ae703f3caf321f5e8e570219b0887da6a5ab17ec533231bf578fac1139e09ce0d232eaea72ad5cb19430a82b3aad141e0eead8ffd559eda4994978f2898c742df025a3568e06e281eb0380bdc94717729c0ede28812c14f9fc701398383a780fc985d7a3c02bc6c51cd2c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h398266fcca6ef7da593b80d834dc9ed02dafbe910c7ef6e00a07c6049edfd64e1bf2eacd673be1d6614e2920b55ba5d9fdc89161f50e3a28f36702cc86bbc6bb4219865ae998d22333f8a3687a6b14c38dd46bccc9eb571e30b6e8bd4371f4798b7710ad8d2b6c56584b1b069f2ad0c04c2a1a0aee3a0a60;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17d536ad907346052f8f4ca7eadc51beeb1484372907916d7d5ac7b3ab256e340a585e29fda14b67a9b9e10035dbe8dc91399aff5e46e6d0b243a3bcab7f1920e51bb5eb7861cd004d1d38e53614c8da7ee01dbbc9ae14b3651dd8b873e440633d544a8f6e11820ee428e72edc02a191357770ef416cf53ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3ef6028cd633d46f180948176dce9f9e0fb90b0993eda3afb45ff6a17601d395dfd61b4a571328106b041b8565b1cfb4835053edf01589cc3e8e03f428b7d1ec64719e394b3ba3bd5852d8c274515b0419e754bb1502d6e4a980747f6f8c9776ef33a48d5b59fec4767f953ad536f32e583b803f1dfbe94;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc1eb8acdc5c5c09b06aa62956aa57a546e2beb2e5a2043e88a1d893352891f0cc2c84f4136cb0270e0e4d1045174055b804a264aff6a07a34dc1d75eada443aa1a86e3283ed79364dab9419829d9e63a34ba511d92a73367da1b4e4493b16e8a88901285654665de34d09bfa0652d24985f3e0a122fb5b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d0d2c351ed42632653506658e019701fc2691668ddea4f3a46470b09484b13b6109312d4b056a38139283d980c53ad5d7edc77a39020c0ea14df5828f8525400493df20a565f8bfccb9cc18551356db2925a61c0373b3ff0a48b8369462107223d0611c9ae0e1c69f4ee40af7145716bacf86fdc8a3fe4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec4c4b4c3628f8d679774b85eeffaf360a806b1257241dadc9b0c10f869bae98b531fc055e85e8090d75beb38b3ac246bd5f34c350e53028d9061fcc6583f1937c0df3057a2751b41fddbbf2cdba65c615584d9593d7bbf7f210186eb3e58aad0cab34c612a2db591323899529ee0709efed2325ad98b18a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edf1334bad89ecceb1377e989894b13c05c0e64c42df3312ff5f0acad6787332e23971dffc721b2092a1a0c4b76c0058cbebd8b5e52a662aa4ca99b62fbd3bd2a2ad95f08d91b4219882bd979e9f4c82cdb40f0ad38391a03f5451d313cb971bbc0a33f2a042e43f041fecf43c1c7b660f5fdf8c94f47fe1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78e503f9e507e45f2f5c6585f831f6d59fb5c3f38ec4f4f15e20c9cd3192a95980dc8e3f2ac14de3818ce6c950b294d9cf68d6ac9116761421472749b7954e7a595f76ed4f01cc00bfec8fc4d2d32c8532b819192acc9ee31994a03acc2273d0781c6fdc65a5937d5fcfe97b74ced064c94c9b9366e3d81e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf145c4c51ac251b69a2778a01a4e2d40fb4bfe0b252180f22ecf58f276cd006ad7d9b87ffd7e054d5cf250a1a3f0430490f1525b25bf419273604d4d23a3c606fad2c364ae018ee1cf13591dd78d1bdcfe6c69a141be2f5ad523343207fbc21dd7dfe109de3552e8521548b7dd5c1dc0ba8a243f3516f4ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1138d56e375f137db565ab932d4fcc03bfaa54f2a03e7fb29b8bd03329ab7b49edad21ca6549afc9338e2c2b5e6d4aa50ab33680533d0456cb17de778fedd3121546addd4d9f5c9c56afb92f504b240dd9b755be58524bbaa0b1dbca26ea1e08fce3ef0033c847991ca73d181e31b3c72511015b31998e4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196c87da48230c4f171bcce6bb2fa98de2e1cf507806fa2cb7db95078dc06fc068eefb0bae79a28efc7e196c7cbb3621b93e8d0de967546e70e1336e0b26f74a3e602264fc3672ca000fe3289985bf0b33f3a5087565b951c6374d48fef1558ee40737fd7c83f2a25fc44787e5cf534c864ab15bd1d469838;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h432b3fa55c09e474345ad8686e746d4217a76cd09694db2368d0ab6887810b0ea2f49af1eba5231427ea05fa0d117749f5088408ee72c950d91c1fdc79e149b74b2af012d549bb3f4ebe9187ad720655f7d8915db5c95573e94ee681c60f5a4b3feaf0d8218d937f264420f4cf4687ea6dc6d051e612626;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d1a64ac1044328cc13a4a41fa337eb7fea254805ddf7d420d9fe120c7b9384c485d2529ccb27f0ea21f5a95d1c820ee88a5755d02f6672b81d907fce62f66fd74ad1b41f625c0cd12e34f4731d28d65e1037515337955431faa84be5f3c16460deacb7efda3115b8c3c3d3ddb3ae0e977d8e9e22303a648f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7dc250378893312e46e0f2a7f3f70d4d3dc21d326c60a39c2adfed8bc62752426cc72c4cf1e63063031414c5aedda3c0022cb74acb0e8450159b3fc7af5ca4176438ee64e20c3b91842d0f6cccef54d99dbe1c06c6f40d67ff102127718b9b240fa8aa40d9042061af8e70a62e23f638ee5ccf9f9484b4ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f766d1d5d3146fb7a2e93dde9e751c1c7b7bdf91749cdd96899dd7effbf549ec62d849276ae0f320e358de035e414516e767140330dc5345c0d058263a4860afb18a45f1e519fbddb9dc304eac9ba17dfa62bc88f9de24cd8aa3921fc100de5f1917ce4a49812010153a97c0f8d117296c9e5a0499ef169;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b0fed8f1b2105618fd3e17f3dcda9b2c3bb2884414be28e91bd479155d36e6cbeccece0ee4975af02f97a64fa791bf004accfd654a89934e4143e3d668b1b448f48081f97e73f7161eb06048241f1e910138df60b49879b0d906ea2206306a1acd61661a36c3aeec5be0af120d92e2935bbf3fb72bbebc0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2edd5e9e347ba40c20e217a4f5e9520905dbe17be2ba31ea8441cff3c1578080db64840b80dec5263e41588e75ee9962a40ae91603fb5819c40fe71002a462ec4f1ff25debd63591621c9e5553d15917a90cbc03e68c90f462c72fd69667f2bf05f6d2449950819f26feee165502f4571344b558bc3922a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1199dcb2f95b1cbd7ed15a787c97daa5bf664ee17817d3ad850a1d4b6b042d63ae6a9dd4ba2981f7879f1d35c977bcddf8fb04adea6132be5944c62e7e8efe3655faaa7402ba8ff7c73371069696755d9b10e97457aeafdd2877a08a845b91a3252cc9e4ad9dedffa6d1d6679988e9c169c1548cdb9e8a64d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1284b0318eac8e69aeb1ab70dab1dbbf26f590d1550196e052e8839d336f112622a4c8fb405ff87191db9ddaecc08b2f5085d8a8f94fe605d1c76a9af3aad02bf727515e3e37c9f7eb897c47a622eb8dab066657be98831ebc6e6f30dca72bed94dadae8ca3f423f0f25c7c02664424da80c63d222341d745;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4cbb49778c77945c46138dde170f30e08aac611cda204616f36031ffb5256680d81b8f19503dfdd4e0ffbb4d596a3680dfd3be9eb2ccac811676e851945cf841093648283b99eb37b0e0a335862cdb155a2a91d83e1ebd8b6931e282708159cb8029568a58fea0f06f3cf036323ed3ed98a01b07777a4723;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138431e26874b9bac4e5c91b2d03a42efd733aba9f42bc18c1ad560c483dbef375ffd32007c0658d38096a7d1a85cc49287acace1070d2899925ee88361e624acb11e12f3be3f386846703d4f181af835c7965c176bbeeade87342aa7f2df6ff773da1cdaf666e0cee330df14b9610b61b871fdbdc8034cd6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197a64b729e98ddee5b43fa4f106ba63a7f412c438e8aa2fc9d55a567516d2e2f537c47a3c867ae4ee8c3fcb649a1a2b0e07d56a26165a46abfb9b07b9dac345cfd9db3a3e3c4b0e7d1943b02d0c04f338559321275440b28c903635e82c1a793841b0f67bddd0ccbf77694b5bf27d4b09ca289440b4c7ae6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h21e0c15d30a11e27d986b1c8f0b9d94d59fbd7e73bdf313ecdc8783c3bd9434b0ecbf28e2ab8d397ee0d3712d46b2229c921770bce32c3a11d6a8b79a2349adfc50ed3e4c74191b72e122a77bc4ac032a52bdbe4ab91ff95fdb224b6c0a985b409705c5378bbeaf3d66b3b853730ab42480f513e5168ed80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfb2e3039c21d62cd35596067549b8577dce796a2bae0cb5f229ef598a49f620e37e29c6671ecdb355f590ffe34a6137d8200aace346fb5472cd4adf55e7a47a19723bc84af851bee236240568e7256f7e226cd09aaf7d37c7e0afdc177cffb5d90bf66cfcee8e1dfe876110385b9b46225d177f9318e422;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18367231aae60902210d57e3c5f6608ada453ecdac7081766d09a3492bb14b4623c89d4a848874ce8f16a162478810e9d99bbb607915147a20ae34e12c67f524f8b673f5aca3790b907d35285976c18a422a07b63591047f23da547886c9b553b7f6d249140aa48c99295ab49572eb84cdc53a5c6e9cca09b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12429750851384d95fc6fe799e3fd38e350f2b73942638999a487c47c84975c22f25b005e03eddade7c1342d257e36e19de747a04c0dc5c96ab51ba02771f29f51c5fb829c5d9ebc9b476feeda3969d652ad7ccfa792db364988fdae2b9f2e39402948ee1dcd7de20ca63cb7d7d196944d393b32c22eba939;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h92aaa930708bc14a032284682bae14ddfc31ae719c5ae5c5f0450d89fad2af39e62c3ad121c2e7b8d5c5a47e741a8e34510efdcb86be7cb991dd9441709169639f9504f3eb14727cf4bce90eb299ee4d61e6f096c4a2b9ddd0ef581e5dbaa88998df77f981e8c4852ef09b614c2644a8512262ac2172c346;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71db3e8dfddd3106bd861695061300759a9a6ec91f701033afe2da700e6c8e2efbf441ed390e6b213f1b729520c2a5fd64c3fd924c3c7f694a67cee179d0a64f710985d4e0b8b9271e1548d70631dec37f5717a52b460c6a68249a5ced3cfcae9ebee2bf9935a2d50ecd2e7479fc10c3d6324140c189e853;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ca186409d69876c9993c5ad3c6647052ebb7a84c674e830568eb96b335f7e642713d24449dca9d7958b1f4fbb647eee2e366c23ff5860892f7e5a6f4e2003eece9dd0321a8ead2c7d6f4120b9cf685560e489c91f1915cbb21ae22f76f91d28b13594f1ea6134c9cc2c74908f943009820911b89ca895ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156be6b4931c981e12daa9930ccb2d0f5112e233d44133f40f72f00d5c29801aabe4b8a607db579a17280cf8b30b5c20868d3eddf7dc2e0c2666245effc81d49c9f888ddefe3403f6417f168674ac34d4247a8c61b4fc2f0e4a72e0097360d41a8ce4b85f8d15c5b4b618ea3b24779645ccb5f99c457c04be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h510439ffc4725cc63e2c9a90554ca44ba8f5e3db2f7ad04fea0ae89fe171914781abad921a7bda4891213ebd02175ad6585e5bcc157b51c83c52690f01e1275d8a9bb7266098d07c8335c12702b2db7895fe5da908938c397731abf44107f948e26f9c107f0ccb62f8a1bc15d4e4198bdb0e83167d9120cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3205ddd9c9206d6d2739c9637e7268184a59b075e6767286fe7f8b08339dc006786a0c3db8877ec20cb1dddfac9972766649a995daf6f6e80e4717689846009fbbb46e568570c67137a76555e8fdc4aca2de52fc9b7cb18421df1d878f3504e7e4db9ec72874d59bb1de40cc5813e935554120a30df8400;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17eedd2a60a911129934aa8017fddefd157cdc76dfe3ea1762c39b1b3bf91a0f3f79ef6911dea4a0f12d5407a6e56af9870e0017cabef504ef23b09a78436373371e18b4133fcb465de14d29e93c29e95bd36f88f6fca8c83cac87b7b2ac8eeb954acbd13d5ad30a0ff099dbd788f8fe5bf9bf653235760c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfed3a67611dc5a3cd0efad75d39fa440d5d9f69eefc159464d80f8658128eb07acd49add7080496957e8e1f68c123464caba99f510f1aa05c821c293c124d99fd0314f24b9f4dd208a2b620c99e0a210fc991711f00eee637a30f83904beb482c11eb11a151df3d73f9a573c7d85bc3d034354220be9838e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10cdd7442220348cf3263e5866e71d3aaf6936370bc3916016f4e7659ae567016a3d94625070dd53dab4f3d3575f77d978f173a2cf40f8c2ff5b9fc764e7fc21e8d2ff35f2374e8890514b68a09c1701b35aac8e7f5f1856cf77e0da52de47b5dd83f8f321d004f8c6b7e4499585a549e6d1a0c38d641368;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h21c905d9826959b5e08b49a9a3e23ce2cce6fdfe52a69762902ec93adf5b291430c2b03db1de3c3c6ece9bb0665b0f65478c517461fd07afde46a55829c30ccb5e0ca92d12e30fabe50d2b237a6cf4a2391b0f4d420afb38f1a89f72ef5df0da96c693d77da88d98c689c287e5d3371ef6e0aabedbfb22b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h512430ee9c47b3f66e32231f6a7045fe77887fe6a6ca88e9bb6a55691f1559111718346d07ba5e4a7401d48ddd3cbf8a97f8d1ed9745aec8fa205e3868708e51356c5ed2002fc27f9f7718cd992852259d36020672b2f6ec6fde2c51a1a18d430409a19f6eb6529da9364a6183882682317f0804435a2e4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc671cc7e3a84f3da6dc220c04e753ccac5607411e7ebb640ac5ab346167424314c240af5ee58715378e9b96db1ae4748aaeda34643178aacb3d4ec706f46034ab868b8e1aadc840c60ae9031182cf0fd444e881d82e19587eddf0db38edbcfa0051f069b07d81efada20e8cf1123172f66c4a1b7c297b5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e111218286d15e4d64bff3cfa339fb181e6aac11750b83d285858e511a7cbef320bb60f4883dc7f87b806442d1d2c1c95376624ed90dcc0a34703702ee1311687fcc5470b6a835bac90171e38cd4b327a1a6c0a00430be4635cd603d71ea421756c17a0043fe0d38da23946656aa887638abe72a14b4d738;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193a830c2b2c5e1f68ecf0d2dd010dfc49ce1edfbaf8054636c59a4481dcf0cc79506d089e18ecf64394bbd5e6e6537aa584d5b29dd8910a9ca70cd173d0dadab5165f6800c948ac8b0194fe186f4a3ab6c6b71c6934006f9b6997783754478cda38b89de0729c83a2319365df8ff6ab69b733f907452fdc8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5eb4156cad22dec9a5fc709f8ccd258311e34252429e955b17db02b7c36871bcb7775cd7930601f2569504e2a7f58a8b08afd696e26674849304d0075975ad1215faf8d22ddceb44c023908bffe9795db6a25938144c2678a0d9dec12dc80af636e3bd4a2d8a66cc24385f817f0becd52d3f5df5aa4ebece;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13217a11f4b1a30ac5134efeed56c20af609dcbf775220bf828498ceae46dafde76a0846a52d912515086e409a71dcf530c0000e213febfd2b158da74ecc54a2ea8a6404caf59c15187bab6ca16e20e013acb83471b9fdd78fe9d1a7495c0cfef3c0d531dc299d2e839cc57982117501219e2e8bf8aed8985;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb73e07163afe643a20b40948cddb281da86fce9ab1aa976cfa55950fc6eaed10caa2f3f336a153218d4c9d3ef4d892b988dd6aa4fb47c36785c72afdd475d817632c1469eedd5f5c058476e45d384390d97be21e3ec647cefc7f49116fca1062a81d4fb29ed5940442d22bd953c5efd7875433db788700e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb15c5e13cd2c45128c3b70531e129b8018c630e87f9dc1599badc5befdab91c5253fdf0b22649e1bb5ac9d8c2afca065d91285c7b5eac73108e1b8e6fc03935d7f43981204629e015d83111695a393e38e070583f11a6cc169edebec5a562c3f0b921d473d5de6b62a7b5adcc3359486ccd9204952c69b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c82b0c05e8a26802d7da5758e80dde10c0639ffba4f54f3d2629ed37a7ecb279c53d5feea6a3725ba1582797c8e30f458c55027c501d91f24001815eaa63259b95ef4e6db81efd23b7af6d04eb730d09a78b116e93c4ece436e175551b90b35802feeafa7630bc01f38b66a0978c5aa6d4c331dc84c89b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0cc6e98706e2153c9163cb6fc3d36de590d7743f6846a8979a1e5fc7edf503662d3a7cd7064e680709dd85d3391e0ad722540c5f3cbe196a3298bafde7ce336c4231f255ce090965d73964517fd1aed40271eee86e84698649f03c54e7f17a881b4b24108bad44fbd47125421d69fab76dcca8061b96b0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1f00cb67c0f930d4c023d1d09efaa070c4e761657859d2b17cb316b44d15004108e72b40fe1051b5cbf47eee02d1d6eb90caf8e31f02901708135da4a5b41386e283a9bc9f16d34270e99a9c4d468413a477c9cb72bc08083dcadaa31a76599a6f910243c21e02e1718289c45754a092e6f9b95fe0d7485;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11edf77fc8ca545278bb164e373583d220df53130d92f2e8878c88c67d3c92de6b9862d6cfd2d2f8e3e802a42d15cc8afc45b5ed1e72e0d7ac94c63cf6f2345e2cb31663140e225e9db26176f8f49c5e3b0386d23e29a3a2105ded218b9712901ef931dfc88f0451c10ad449d1fa4decfef2284148a28fd09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b2a253cf9ace2a7ecfd8e1eee3c8f547b510b4553ea9f986614212126fde0401d56b04f6f5c5d5620087928e52ec3866b163eee24f8f1b9da64bb948dd135f04f0cb9bab438f109bc8f5eaa0ea7a27c42be6be40e79ee2b6776b041429dae5817dfe7b197c9d7307df7a32197adf74bf6344b381e4d9ddd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b53eb0a59712c8e31d6a12b917282d23a1d5aa47e1d979ade15420f6b2bd62916911f7d046fc8a6e7d463192f4367dea6d4824d98255c53e2e22b5da19be36fb6a105cc26a67f3073a9eec8b5f971ffce7b48b54042ce55fd0d5ae223757d056847792074c39cd94eef1103488fd4436d48b14139039358;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee7bf9a169aa4285e85843960dce868f45d055cd54ed4564d4fc848610e9719b7e4f0196bad76209ca520ccb2def17c6984c0a232682396e186b3592a057a48242956e7b66851d7cd3de0f1d5a6bc1413c695b3ba6e213c6f610945ed808d6ec5cd8963aff34d895d7e30af68af404a5f58d15b8a9053b17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1000b85ad2490e6177ff85f8708838a7b8be6105144d73f78a802ae3cae1d07c48377cbbfb7e7b986720f853529e731a3eb7b094d6da0f58c50f132bc88b1aac88b79050f228fcace59a1f4324e4cd1535519be613e0164b02c29c6d39e0948b71a58a03c7568c5f1180d8973ae874eb93876ad54d3a04b93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fbdab44c60ea9a1e25168c35525bd3c73e36f26ba4df5a5195f1da91ba6637620326781d0f8b02cd3c1b982c92ceb89e6080b261b390e926b61157453029bbab01b73f0136c61f96d554e3fc308ee052727948ba6438d088e7b20c7cb735e91be2f0b7fb1d6beb9912ba25777bab0d6eedaf0c7d31726c16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h144efee8ce12df4287b5a4dbf8c5e3518740536812e51f3d77f319615ea1887258013375af1a798ec3448c05d59dd0727bf971e6596a60e94d9df68a80f6430c597b79cb3167099178ccda6a3e45a1bbeb1af89e97204fc9ac91e2bd68d01b77388ccc7b1e379cbdfe205e4157910356480207bba391bb0e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0c270b8ecb5a6a6c02214a90e270728b2f94976b7c7e110584b032ab9cc61a889b0f5a1a4c62b220a7d0b1b281ab09ee7ff9af267e79eed15b89422cd6435da727f9225c9acdcf5dc00080792594eaffbf69a34bd10cdc9d63098ac1e30fb536357be77d8fcfc8125401c28890b584b4b94f359e8ccf7be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7739e6027ca37b15dc56c900201981cd89deb7c1a7075e70cf7e4fd62b4cb4f6e09bf8fc131e233185c791b9169a426756c5f5b3f1dfbd91cbd7a9d499cc6cbc626328ebf24e5d8f95ba6ff1cccaea0b84fc5e1f49172b1a98c9ac1b1afedde08694182da4ac01d4a36e4e802b98e8c0f997fbb89a8b3e5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e07d23533ce6761a2e4f95a831122e5969b35bf29543bf045faafa12d5aa932d28ca832c5c71ed4771c5e95e5938f6a937d9a0e601c4b255f35da820191290dda6f8ff0dd653e6198151431c6c96a78e9e450687f4e5b3bd248f6f3ae0c4a686ceac291dfd3cfb59035b671e78c4a4d5e3506550254c580;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b2d220d17f8455f9e8adfab2f6302252986550d5b4245d3f1353f3622b9e1ac495e2dc1bcac732e7eda02813762a82bc51890e1ff6b27f252e7e876a45f17f0e58f0c84d896c13a8de27786d4471696002c80216c0148fa4414f5a0965fd609d34602578ae06065a6c9d02d430b80e70c810c613724ae11d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb67c1c0a5542f4c6ed4464ce9fe17bd65dedf1cc68607f14abc73a040d3bcb49c76fb468ca2295f74e3705785801d71370275bac08c83ba2b30dca64787f17cf5ff32b8014e4768b4b20883bd5e20afd1ac02189aa9e0cb313dd2d37fd956c2c5de665821c9b361065b73119efbc454de72ee795d146abed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12317eb537f61b1ba18e66f6b631e15503f2225dc62b0dbef5df63ef340b4808591b557ada5b75951371b4110645c15f69e0c90abfefa54bd4319359991aaec1cd4b37dbff74f83de9091fce276d787df763100fb02864b9f10f12e9d4e2e0337ace849d3572b9a567e7f05169ec299e4f2d20f866fccacf3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h100c208588c5419206856f35a76dd60ae1a5920e7905b13de024ce51656870bc33064a8b72fce7de1f04df2634b46ad695211d58d79143e91a55f257a8708accd2fabd68dd5cee9555e4310fa9ec9546f57787cd8bfb954fad7e5ed50894d206bb3d55a78c19f3047d873577e524a6e5925bf39d42f8a63be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5c4a1a6e19d7e4df95e920e9ddda7554ceb42f109619eaf1db7bb2aeabfb8cfaa220839cc7bb486ea9baa25bd1defed47466ede3282bf2d74b449010cdf959bbe73e1d3b5cd78f70e0f28376ca1f354b65487a4705339a62b6281bc31e14f82a109981a264382839ac7ef5d1d07b717a950b6c2cf076316;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b224e3af1e381f329454b9d6f153302ff8c5d2fe2c51c924d301f80bb39f4e8ada0003199069471aa8f37a6da282e572325923ff7a80c9a4f69817142f72b03e92e9ad06290c0b1d4af6026bb7805365b1b84aa0c07c94550ec683bfe77e3f747e6d093aabd048f6f15594fb62d1601979b5ffa6b9b41a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d36f40d67a692bbdbdc46f4d99bd7de6f6f44d5b7f6e549430b4a525c7339eb1ffbba8f5c0df8f9c80335b220e3fd2227258ac4ed50e36ecd9d2dd357034a1e6d3962152d27453d8b254c13f0779844b8b8f18e79c1a8aec1c81ef52da3b9bed1dc1b3d072c3d5272694d038119225525b1fd93151eae32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h188b013d7af84ea5ee5f92035c88d7fef6dca65a30e40794eb95b227231c2391fb0a147e48a8862875e14860a80091cb7d6d642a9bc97a09081398dd7c765832fe798eff0b3814a791d767773b2cacd1ca6d9813e03a355925bd26fdcfd4914759aeaeb934064b46cf509fb2d70b3a09dc50c49c07b44522a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82afb2c735ee0069ddf89f9792d007e885e650db8c052a70696e2ee413bc01ca5b41d480473d1a48509a094fa3e83942c33e7b30591e7537389efbb79818873a92bd82e06ec3f273806105a5df3f1fa9a3958dde81a6b93a7cd019e5d3dab4264636706ce04493632958bcb23093a8ebed1b8151d2c93870;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc79ab30bee1d23969bcf35c4aca359656091c9dfcff448ced7756893b6a93aedcd1d7c4bfe9e868490fb910e344394bd6886c7a575504250dff2b63cbbb3fb62708d6d93e6639a2e0959ecd57c738dc3437d4b04bcba5b82f7fadb3dbd25c1eb3f680a50c80fa3dcfb664de797efdcaad27e508593439c9d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heabd8466df65448debf5b545e2bedfb4708e12a7469f1e57cb5b0b6cc3b68960d4ee3da17ab7d3b81073530e99b6609c9d8942249f1deed6786a5e0e48a871b44f65d5d312f19953728a81b66a034969ac72b81d47a3a6485455c9eb5656144ea29065dce01c898e7fea6f6bc23170b8f894a937afa4ae4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1000acfb17891343ce655af7264eb4a5acb3b02965d2a64f9df700d6fa6d3dc730211e758b54549637894fe6d14d84c935330a788fd7bb9f96da19fe926e2cd3d2ddc702a240a72903585296eba7e7402ff3a8174ebff5b946cb6d93ef26af2d32d1b5e36de655936ae6b47386a245cd41f96674c1972df98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13aa9621d69968362aa06ebdef5624fedabcb97f59ba862b3012d3abde5d2db19aeacfc49f1a9df5fd7f84c989f9d560083637e60c8d0986738ee62be68d2b431e31412cd72f4e2a9480cc22928f96ff0f6ad7996c10242598895ef2f57045a85d51750d9f6664384ba5fa23392abafbeb6c4fc849a5c12d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89f3bcda5407fccd278a02dd4203c4cc833583b841c737b3c678d974ee1b1843da5559ded52319e3e02aea36a468684541b1bce259a94891314ac9c5ca81c5fae311fcece0e5ece88f4e16e894edfcf28f6d6d6385427cbf695dfcbb211e99dd33f0c5f4196b61f35cf2556eed5188f18152197718184be8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2b71f7fba91fc81fec8de37bacd024a3c6374c3b72fafef887a419983e8aecc62752c5ffdc0f92999d764f6b6366ea7bd6fed384429343e7ae311c65b20ea4408306bf79955c82deabdd2ad89cbf4197a11399913a20777e2d966aeea22e4d06f8d8528605396ceb754e3cd78981b354f849c9fc5d16bb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d38c1bb6c489dab3446ff99cff6ceafe9772a1de5007e244021e2289b81e7369eb927d1a38fa9a3325e123125094b0ca7c38647b5e91187059771794cc7843275dbea7b584f081ba5e3dece1fbc14d1c05f5d83207e8b1af6970d71db993078ff8ebcba80b8b9a72f5cb1f833a6909a483588e13370dd93d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b182aea1c710dbad84f9ff6b5559a584e9ff77748132fbcdc70d785d9cad361d1b8d487a31e5512eaddb75468254e34d6a3d6af2e8f733d0b7fc90bf9b24eb885d34c7cb5138e231dbc8e6a072fdbb3920d9b6d8d35a2868e55f0cbe37bad0d13068b31840ef1432920667965f6d80e50f064c891d87d3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5fa0350bdd1c3579c15b4539f5e8022918ded0d46f914917b84a8d1820c2c00c923803a583c12d1a3a6340960973fdee08b424db9facfa3c28b26e9125bc8aaa8ec431f76215ab527c049832cc91fc857226c69626799e962c62935eed11af4ebe52382441a89ce24e683c2fab8b20eb1c8ea4a68027acf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef4f3e09853b4b39ec614a30d087e5c8987a80fe32fa3f0248cb0a01bdaef2bd28fa79562d84796fdb3627a6c3472afb09ba007980a7df3825047745a59eaa10fc5664108eb8b1067b5fd1c95d632e22cc6ee1be8d45dde60a3939c95d9f0b48c369cdde861d2d485ebcc169d44ea687d1a444b3a8aa48bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3da8fdaf851bbca8dfb634ac7ca54b575cdc8347d769aa4e16465dad840962c1d208ea8f65b3d5a99ca4eb9ca95a1244db3320d41697ef1ee3633a9cf80016b3ac10ced1edfc255a94c4e239b691f52d68787d758958d4401443e5e5753f74028f8b3409fe47642fdd46733bc3c157019d2f40b3a9c26824;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187c89b8ee611b8eb641b678ea87e754f489daa65d5bf8a10888a792d804d4637e856b3f9cfd179a3fc629ae9ee6244f23ae123c61e5572ee4da0abbb6fd4cd4f9377472ac93071ac763e7e29e1f6631c4138d2a482401a42d84c42b5d9e5198d0c7b71653a00efa83f462fb7fc839e456f1fad266c11228c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d76a9601accef9729b5b6c4aa29990bcbfc1b998e3cc856f59b1bb3deaf52c1c6b61bef0dbac6201baaa741d2ed38549fdfadbebac09e5ba027291bceaa84f81af2dfd8996d7d315d786a22544f6477c86a7a2048869c55d27b0489266508cfcab0801797ab565dfd713a4c30023dc1439ec5916da57a0be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172d9be9c3cd3d912419d0b926430f99bf9b57ca47befc5de7e844160e887b9df75d1f9c1f919a72c037baa456a808ce419435f9b362e01190b0877658827fece15b312c34282c914857724446a5cc2df5313be16d8c94a8ae0ef9d752632257dcf145208abe8259876f5c08196b94f598168fca1cf1b9213;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156c7a30771959701fe4edd1e123f6524b03c738bba262ab239d5cb36cad9452c5b820ada7789354fdc18910532b021eac60cfb7df4f8617ee18eca7fd41c7d2cf8863ea77fa0e1825e562aa923a318f1807e1d92cc1dc9f645a9d005c5d0c4c6b6e7b72185fb8f4c24176c69505ee8acaae7be39b918d95f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5537bc4da747c916a585f2e34633e3d8d892fd17b47bcd040540548800d4f2236069632398cf27a90b3740a53687eb92e11c414334e515d4a1cae793223ff67ff0d33b4585755d314dc2aeda40c67f17203e2b2be4cf0c34f9fc95f3ad6f8a5c1616f95b772cc455175592e332541f5b94f17e530465246d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbadec6fb8b4396ee195a6557b249d7b0384c723da49252308171ae5985865f606b9bb07cb928fe616c9363956f882ff4ad3c7df13a41fa7a72685238564328a053ce789760820c0ccc189c8bb6e2ff6c2c1a8cac815ed335317ad8bedc210db88107328fdd01a9b4bb57d5c25ad1f0c5676dde609cca6db9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h97a740e06d684f00191d70caef552dee329262ed2d3257bd1e518ff7fbe9cc3ad59c714b7a0e21620a5ba87904a57751f31a4bd17e8f8eb34ab0483c6ca44fc2612fa89518f394413afda5d0057518e9e885a3fcfa85b38581a9c43a4f361bbc6467c9b1cb4acb07e97711d17216d8d5d4daac05ad98cfe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115cb129d928c709ce09c10acd81e511dcf4fbd54f5752e7f9baf7dac2dc51a6f347672c9bcfce6a42a18d8a1ddd53481d09a2a425e827498ff2a9a66b8951680b47b7f35b351d64e5f60265a74fc2eebf752c1ae6f2409945e6a937f5630adc34011b0bf1f788948eb42bc39bc060774824158e33d59863d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13187b52fa8bfb5afe40fa3663d048e10246e065894c0c9ec7a3f5222a0d53047b2bbc46b784586f07e0b5a52f228fbcfedc03fd1cfdf78e445efc6c4c85f9dd46431329e9c536acf2aa326f064c2f63242c76fdfeb05a8f3fe0f9a3ae07c3a72760939f2b3d8d26ada496dded4121511ed9f96e8cc0bfd2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4f8b89d8381eb0449cc1171024ba49435fe22a372da144e0b7820b6593ba62e217da6452717c97c7a73396d4a9754a8b5e3a2936bbfa232892aff9df8b39a687d1e628e49dc48d30510a14bc7efee5c5c0d4eb12c30cc1e826e59cc5254fe1f41a9c908419fafb6092b064db939f4b3cfd6c6b718c7e32f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ee5372b7a8d84e9c1075b22d7bb6db5e6307abef488e28dd3d690943203556f7e64a83ad708bda8d29196a38e1e916aff81eae37a02eb730fd2a5c2490f98167592a0293bab4528a371d14069a32b2c327769c76acdf8134f2b815005ce017e94ce6d110c7eb047e3ce0acc73fd845e83ba8b1f7f71cf49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197b111332b6b4d5775c0e02eef897e400706f20eaa70ba4d3dca365413550f6b447dc5c05aebb327cd0b725bc7fd8ce905025b74c5accc5c743a665e9228e86c054955b970051cf936feff4411605ee858eebe990fc3ebe91085692c434f9fcabe1b4db3258651a7ff8f2c9a099a860a618ea16f1aa7fff0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d99af2d637ce74cd911ab8818f7c624e650fab6c2e16677347d648ca3de67ec9c6e95671d3c905b7e9b227360e0d6f48074bd3736396c930aeb3313675936d60f05efcd940d4f35283a58863fb393cf61df48d46ca9b065b31c50267e40e36956ca43edd78cfc4d21cef813a33ed0093a0e856144be04d9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h714628c3f71f31f560c1139f4e4b04cc823b32e84a4af427ad383ed93976df28cd979bbca7338f59d707bfaaa43eb20564da5ed1b87f631138dd6dd855a9ab6043937fb973cd79766f53e5cd62a6b79e746ae95e795647615633d0f71d4acfaf650f3cea3eda3e39278053e5fa4fbec682e5a932e5abd7a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14a158f2554b60c11fbd999a48dc1ffda98fe24f3a20d5403d684df6218b82ea4fe1745b9c0d088c65855f799fb56c2c718a1962a4d06da2332c2cc76ddcbb8c058ca550810f9d4f48f2ee6c32bde54ffcd36d0c377cb15283678918ad15222bc9a7811a191e53df6b3477685f0eb8ada09c605136072fb19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7bd1c153373cbc4138bb86c84401bc3dfe6af74d8081beaa0cddafc10b13453072a6696c23ae1dd16ca175fe5f6ba7394e4b4b9c17975f4e238fb055145ad32fb7d77c200111f1f6264613f6a5dc1b39ecd437511a359e47cf126d8b56db28cbedb7ca960a8ab42259ba28d548b783b592f80967f006c6b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha01d2465e4a2e3913b54d01afd888c3d71c50e7da44dbfb603c1da417640db69e941d2a9ae0a510bc7b174569ef30a9c8dee9303b631ef95ecb0e18b31d7144f12a7bbec6801b8af425a6e5168563115f2dabd6a44e4c3096a9f053677b00f2ea9be58767c75098194ac39068721f9d9bb93dacb6cc69ec3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc7dccc91c15a6ddfd5b766d20963933560ed639241aa31c368b3557cca3fc290a88428c23bff62b366b79075c1c587da6ccd9e13c0b779051e762eb0bf1a6608facb085d0718e32e47fd71537c807f989df697f7ca6041c60235039f9f59922fef7845bfbdee8aa40541ed6405cc80e4f89d24c5cefcaaef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3712f8d2def598fe5f726ad8fdefcbeab9dd10b27afdf91a7a1d8621810c28e520c9fd9b208730b920a0e94268fa4a669bb5b856c1137ee796bd6d98cecfd60d436a6db9db8de7a9382d59e22e1dbf75aed5c05233151f5d29c29c4bfae6654d13c23859eb6d7a5954a3a7febb3e10739b2f8135172094ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb5eebf5f8d9a66b5225b6510392255315f4f26a0ded4cf360399809e91ed893e98266897caa4748bbdf04a5c5758f3925191cb9c87e8c2ec5dc069bbd2be9cb28f4b3eea05342a435829a34fe68cb55e8acce09b284a635fc1132942598585af35ce62b4ef1284bf1ba191e5f3866daa2387432b90369d38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b6aaf0fd5db757542f6e48fd4862ba71a7d5d32cd932e82e4bd6244cf7a7bacc97d41b049b6152d06d0fbca6e57f60bd46affe50ebca07d6df89909aeb5560cec2f4e5328251cbe153fd3980a21895f0116889aaf564ce6f393067279189985bbbfd47d272a6088f51bbb2a7982ee74e96a776896e5301b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b959a0a4cd1242d88c6de5095ccff7689a764983e4ce79e67cfa1f3f6c7758a26c66a2b7ba7e1b2df2d30e41d815abec7476720f0befd9839bbb78e68c78b0c30bfe41432da0bf7302e53e7774d5f2804865e4340680c60383632000e084edbce9ac50433ad1e6cf5f216e6d584f376ef070bd6bf943d93;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ec4e62589ebab690ebcddd32cd6d7d609453405a66118ad5dbc9331db25eae8d2860132c01d30637405ebf79827f894f397cc5189e486a0302191374cc928cb3cc524c8943f00296ebea341578d0c496114d9611a7b680ae3eb9a9872cd8c08b8080ddc77d36254d0fb230e2f197796154539c7252618b51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d3f7da436155bfea6ffa2520944f571bd365f800529e152f6e93ad050c24be0e62eae9ecead7495bcb0a5f102c9625cc1e35983d54f5f5f11bea3e1304b261a28576d2dd347d83920299fc1308f6ee85cce8094087ec576b3495512710a438c46beb6eabba131ec3d7b6120261479236b66ae63e4ff00c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a5c111053abcf4d2ccd79aac5349328a8af3f216df673273ac6b85594a9eacc4d6288710c6c8f0512897f2cafb9c91646e7f4212cf2f95bd87f3b00f24316d926392ceed5377100f823f1c74fd49a98ee92f33e08162a922f6fbb387b94902339decb3a456816be927eab2d486cb58c8745ae8762fbae8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4dc5d7013392e263dd9faa71fff8651299a38001e0d1c4d0f6755f07ab08bf33807bd084bdf3e88f1b6737354c697067673d70c8e9a5721f974abc7631d07abc9651e073efe85ccbf02eb023e6201b456a18deaa024ed9f12bd6f041afe46a2986d4c8076afd5c3f54d324c7ceb9736fa3d7c61ed58dc22e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf815dc4dd6c81b6d00b84a2c2a10ca8107a2d31bb2b8bfdbadeb5f1d338ccf6207a5fd1a67688adba2f5b7c052c651fc2e0afdc17d24e4519f588e2e89eb79784f373a1a42abd00368e0f1b8af232a8c0b4eeb4dd38ed981157fc276c53562d67149760d4640778f3a48da937e44fc16b9927e9ad494acd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a55ac7f753d63480942475fc96011ed035ac75415e879dd0ec59e781c7f04a6cf80d4e11eccecf0e881142840cac4ffcdaee2a85f3864df14ed06672106b083d6360ebe404e54cebacf72bcce3739d7fd86822a2227aa75dfc3d94dfc3df92fa3acd884cbbb559e43a1d5702243895dd9f431736ff523e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h145e2c89b00cc5076903e711715119d143cd623d1ae4d08e5449752f8e06d68b2ee12bf29f8a71f45a43c852683a0ae57b4b277c5b28e5ad046fbca9352281680ea2333628f851e826b156f101bf8edac9caa28cdf26eb47490fcc83fcb7191d016bc592561f45c1e291bf8a7ec14664b5607a1b7e8bf7cf9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d02d55a9c77e41be6fbe896905ace31a746a7f5b3c722563a2e89dc55f920f2f6a5624aa619bcee6a09fa13934b17d8191f226b1c4353729194653ff4352fe73a2d2e230f4d3c2148af7d6296ab3e8de8d90dbe441e376c3e1fe8d01ef5648510f88fb496eb9d3111d892647753e16f8c2de54f264de1553;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84b32adee00a0be0067ddbbe0f5743a23cf06387f9672c0b1cd9af560232a124178a7416b7407777dae5a6d1a07c4dc42bb7b3a52fa7d26b2b7be04075e771f691be87f46389d68ddec38d4668f01f24d3c5702d6602e0d429b07f92f11c663f9bd8b48e71ce2180da594569ca84dfb4dae575948105a4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13175624dbbdd3e930a501b8b80fbe4a414d1999e51bda6a8176cab29fdccd9e79abd11eb043666cc4f0b30afd6d3abd50bf9381a4529dff27c7bf5e9d4ffff01166003c7ade6cd865660f84d6e7de717a7f9726452ffba03f89ab9b33c83c89b58943426c32e722aeb98c1e7aa189b043687012cae6357dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0f2cbeeb6482c2c73e7eec2d4c6684bda3eb0cf09b9865c6a50396b56793e22dc8b0f38bb0f9c83780f60f9ed002d5de51a16b63bf2a3418b0e89e37490b7ba4d4100bc99f300449a2f877627626b768c847e79ff00d62392067f5be2c5505d1473212568ec316bbe1ef062a533a970333a31364a89355b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb003fd2f33f7875459f6b23ae7c3f9e65e45c277ebced38bd726539eaa2db8c45527cb4860f5c1d8a326d98d1118aad43d88cdbfc6556a55a310c294fa934e7cf55298bd99b2be5f27c4c6b065752bb3650c72d4fb618fcc7029d91f74a176e9836c258d7728efdb7bbc7907c269fc22734c8bc42c6fa41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h116413edb012231fbae7ca687aacf5f4715ddf04a42db317a15bcda8d7f2573f2a2bea7f644a23ca73c549a0079ff96202d906179462ea4b61d28c085349ba9deb753f22245638996cadfbd3da46e31d059821e0830c3f03ae19bb458d13015b3f0f826dfe7eddf079a648adfb25728cb6f57a4fbd89402e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e8b3e1b323123c81bc3c7a0f0d7a509e1d509bfd2b25c25c5740ae1d9ad03f9b34747e1cb4000c467f78974236ca80a9ecf00838f538e6d12f6b3037a2b231d495243c639a6932c0a67cf62dc8e750d8c7c9cb9e9bf7368fb2b7f6a0d97e56184836365aaa4d1faf4e09355be2343f880cb41a9cf74b9b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8df1b857027f8acaf0e44309aedacdeb45d4dc417bdb0662e90216011b6a1e869b223e32c897aeef8fb51ade34e247d38f5c0311e65c001f25d24575bf093fdef0f6f9c5f899344bd07b06e03f59e409bfe1d20cb665cbedaa5a11b4e729f8a419ab87ccb7a3fa70c3355dad7228a3f3be7ef2a6f4fbc2c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f2b81feec3e50108e3ba10041dd128a5fca43a346137c758b7b4e4debac19944be5520d996a3d633a9aa8d20e9f815b447ef855f27ffa9ade99adbcfaf059cecbf11a47a746681411350c93b17de2d387319b08b179dde110a3723d67ffea2f9c315804d091f00c1460cb1043745fdc97bec2ce789777d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5136afdaaeff7f5ce1c4c93f7e3feb39c0ff68fe4c817615ea9614e7197750bf94a0d8bb3a317fd54ad6d5abfb6088d3d553f13b497ec5ea3ecd6aebc36b682bae4fbb1f428445cb061b9ab04fcd5e2f7ab06c6aac2a28859c69b82bbb31dadf8332c0782b24f7c5059af9879478e2256a639f4b835636f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2b236a713a3abfeebde90e93010078f5f972f20c16a7a879ac5a600d9fc55b8b19792cb94925adfe67ab68729c933e20792380c2b392e9dba088ecdc08bee5ad80cbe5375c79441b0fc9cbc4b057436a02af771f527c6b3c6a50a9f13c026df0bd192413f5aba2112f71bc6a044d6b94ec35638770dad19a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ce8c4ffd0464ed09fa5cc5fbae20f1288c826ce9983259e1c06d042dc6b9fe82ef1569cff2dd8fe4f6316736378156755f28d7e21aa21222ec2ff1d21929038d456e214a0bd71eada3d22293adf6f901005475059a66f5418c6ad022d2dac930de6e351e3f3ec5963a09187cc2c89939a4e0eef5aa32f2f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18797df75f980d9b2be25e16fc9d4bdd38ffe4d206af405769dbe8bb26620b8f92b5975a31ceca99320c7a6d8f354f1101f7db36728fe62129aa2000cee6e28ba92a6f4adfc209aac8a28e67e1230b11f76da30a5d8e81b1291bbf710009895e87727d0f42c78a94fb4ec612bfc35db6abe112acb772101b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160d557ff229e3828e2081d635368b8d3a6aed2895a8e42c1a3cabc6598528f8f541be11859c1c3f8d2a5a621e21b52a1ffd12dceb3339403e4a91130e928d961ccfa2d4b31c0947d4d7b56bf1663ef51a945634d2fea7f1b4bfa53fab3c8b126efc30024dd0c9a7127a9d2b80881e77d55be7a1f78217219;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h110e2bc16a20f9091c577dcd90f064baa5c3d1055ffd06206f893b768cb388f3fafdb502e08e11216e135a7764b7d4022b0152b419bd9d9009142ab6fda11a354dd25495f0d098d64d3204d40f275e295325e356dd9bd831a9dcdd735fdd78ae45cf104f4a38a17a81bdddc6f033eeefd024dcb22ec483221;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14369a6b8ba50a04ebfff5093170ed78d865c7fb4b45ff979a0ee6f70776e6114d05ed88738987117b79ab8c573b15168d916be15a6fb0c7c2bec2900cd81de17b4a4863a5899b5dcfaa698a63867dd639f04a52c764563184b1c01f753452c660e928209d247730a9fe302085c0b095c5e818684715bc808;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1074a2c4a014cdc6cd66fe90bfbcff6a52852aee5cd6d501d4e786975e79143a2d676b5c41fa84b3d86ac4e44636a0c4b411443b4fb6635c4770b3a7d5330f6c50a16c93de5bc478842584428f9f5ba60aaef653acd9710485a07fbae44399e53e6f5d7d6d2d07ceb9687d51087852c1f9828625ce30c463d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fdf5e459611babb6805c01722db8ba738512c09d681ce658c25cc9c5c43b301bc9f7a97ba38af04faf7bc452fdc0daf7300ff179029fb1686c062666c7db419244972f4c543a5f9fe6f43b334998d78b5ae4952974809f95c740bdd1feab19afdf38e8f077d4d9c21c57cf4b33388e84c3a3178c4db97260;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c6e50d43ee7414b85a11fbbc4a062d86fcc95211d624bfd246e22ec9ffc5c24be488c7bbeaf6dce5d4bfe077c3932e53e7fef49d6832c77e6cfa0d92c3192c79963b91f22ef0985b890197396ead1fa2a8eedc2a24e1b43665c739d0b1f1cdf4a4a9d67e2a0141f5025e3564c7faffa5451c31e47ead0ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf169ea16ee1c771288351ab8479a5c993856381ca6ce2119df99fd6512e1c4a4b0657ca633b0f6c108c0f988ce089a333e7645ab1049291e4c7ca43c306782bceef7f22a57b517bd193bada9c20372b0dd4ed28f41d6564009d832ca8432c3dafb476e47b2c79513d749cc9a1a42c217e14d5bc27bdc2498;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdaf590c936265a8f2cae2d208d50156c4f09bfe9a63ddd85f5dbe56edd3be780e62c08b5031cad9c0a486b231bb220b45e75935b9b5eef6cdfe95882268ac665e79f9258a706d9b99fc692525ce929cf4e392027c8d035944af1840ca1c28449823f88f0afc0a58edfdf4a07816f292647892a57944659a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a659509916a5c200bc4d5072dd7031e3a32b75c007b337f28922b2648152270300c876aaed32e1679846b652181d327137375357417afc5aa0198eed78f6a0b28fc44b94bb3a76c5caf83ce774de7a7aacd394080e80a3508bf3ad62fbd48b3891f9128563483362b6d81f645b230f90acc7eb3cbd062fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc388735d2211aa964c56098dec13d02c799634a687270ed4bc2bf7e77093c290408cabf654f240403bbc2cb61723efd0577c7f43c1bb6f3bee3502c6696cc12b143b5046d9f25c0f196b7ecf875e71e0b4178acbd1a3ea29bf3c450e80edc9de951acb52384743d6e431b2615d48f93217df5de6c300001;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1138263c759ae55278740d73a2f6e35ccefb917a79b7e96cc96ae6304cb371b28fbaf8589e17279aad6c5821533b80ed0ebff04272add8656d935b139a6f2b627514e8300808c720d2999438a323c5b4afc66b1e648253b4324cded262feeff3abc538c4e85a5c96c4102f9db9f1d9c02c9334416c7f51573;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h171b2b9a269018eea1d2ab91574e5d9ff5d8e77851a35c0090d40c7111a5bd707bb363cb3f6c5b49136583d0abe85973e921319ed3ad964f75f804bc1857451c89a32d3f4a49302bc8b83821275d95667c37a15c4bfc4c51d928006f448d6487bcc09bbdf1cbc0ba74b5453789dd591c90ef35c7ec2a5c57b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16892d0ae2264401bd1c687462e9c97ca5880ee54b6533737a09c1ad78fb78209e2f2549b88c1b3954b6f57bd9b51cf30ac90b31062206fad20a2663d6744490f0308657e18816c1beb56c0a35d5428f127eebf46d9fb9f76445f2578d46004f0182c97dcac2bed2e4e1137902108b6b3f8fe5864217a0f9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17228a0f77f0f0c048a59608a2fc853aa63b4acaabeed556a90d9341dfc5c075fb48b453c8d6b11985f9dfba94bc81653ad4df9b792be2a32f8ac09fd0b8db0c61c9182dc183a937ea67f9fb860b798917f6a466b9120b8284d5de42b7198715417149a9a2eee2730d47e0d1c8b2623cb6eb08e5e8a6ebf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11253cd36a9be57d3f01e586958907b49e2c8129df6b1c938db4d1cf49a8521b757f591bf47a1c8c1cb645e7d15e07b91d2b71a7b6ef8e3f092b3e8f99fd60022567f679ede3a3afafbd98fe5640a506252eda7134a8a36f2a404e7b6e73f9dbe871a8db5325ba63cf2f262868be8aff9db0ee4ccb1e9a170;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1efff42ae999cf1b7688623c31f1f6eed0e8e8f28c27985d4ed15c5877e840e154af1d4cf41b00d27c107b598dede847109a62461b13a18bf1da7293ecd1340c57515d4e6151903b169a52630c990f8b12df8a565cd308b20460f449fc094e672bd9b089738d55f22d0c79df90ad8478d7f2e295edd75047f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h235c7cae88cd07243b977e5df6cd3eed53e8e7ae39555b2fad92872ce74a38d49853f7e0b23a20d089524cf6c492134f358e248c7928a0c43663896d540601864b729bced16537e32b4834430531245c325c4716086d52fba2bd13613efef7751446e36520a10e4eda6f9efb6b461c2075e6adc4e8a9f6ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d75fba68ee848569be8e2b791115a6d0511602de16b5b83949a9c808e810e7a45e3c945d058859605daadc963b0f8cef7e1b837e337e3a0b524fc141f8b976c5d32c729320ee5ea10138ab77ba3df0e4cc80e62e72501a15f8270ba6bf33e03f8603194552fdcbbbf63680869060eca1c0c87358bb5187d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2fa85f849c8d630341e635a2fc3c86565f5faf9b5ca9f5a0ca40cfee5e6ba8dd203f64a6f0b6db888813b22d6a2ebe6ddbf26a067822b3cc8200018866c90ce880fb28a4eb77416374a98e1305c1af2736535e447bc0841ef89da3e7e1066e32ef8efe6529cd5daa19d8af12d8ace55aa28b816aa4c7ebcd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h153dfe44e4edc86ed7bacd11cf42fed7fafd2041b413930692c7e3c199fe38cddbed3b0d0b4ee177a137d19b9b787fce87a85caf63d0493b2aec2cc4124cad0c6ff26fdee5dbcf8289eaf948a9acbfb8cb0166673e7e0c0897fdd355a915c1d6caeab9f804a90a68d80f9e9237783fd65d463e17a0dfaef70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9ada53030fb23f56b34d2d968a332ed25ea6ecdb062294fff06da546899275aa18886ec42112fa9ff1f83f5a9fc5f85e4d3aef8b623e4b97a074987898f918a56a13c0e6513e8bb88ab53e54b309e286085ba447e6daf78a75a9715b9955afa639a1ec95695fef8f991b4a3bb4d857075db037da5fa44c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha69484655e3003f55043d38c371704b14216d1c0c16bc337250651a835020547d2f1a05e4eba6ff1dbe22d2a6296551a9bc07412d842f39d10aca77dd9951281ef6df1fe726b6d5f69dc18eb2d515efb1ad05338d6a7d6fcb9464cf2abc0f538e1886443575a334503a60a11efcd905db584387d20ea7d70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d92c3c0655e9ba0b6bbf7bf478273871cfbd2e8f4e0ebb31eb031c37568ed21ae16e085483bd17c1b634d3e65312d3d7bfbb66743390c13399f1bad2b926f4f3cb722469f2f0e7eaf063e0c898c600fea5854fb137418d47456e423d5cee2ae35d8b7c2d875a0ab38b43e3c01de5d16f471b00f51a435a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h153c2877d8fd6447f581467856f849658ebad99e55a510e8612e699fd1f4a6d2b3086bc677afb9a15451f00eb32d08adc905caccd6346595b31baf31f856717d93bdb9a9e005c2c85d81cb63ea2e4177798eed38d8a4d48ec4f9e812cdf349211596b8a98fb234324d09771b414419c1c02ef5f846f73c59d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3446c394223e053c0809c15eb78ce3706be484c9b39ce1ac766e532c0dadd1626635a66a7350271ed4ef2f649d22d8691ec5c55f2bf91579465c5471a112a5dd6584c4fd156d669a661554d846b7f98941d50b152b345ac401e1621ce8e2a33cfccb7035595ba432a62890205faa209f1f7a131adb3678e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf08c8692f29a3f82331b00804514ca4d88b875589db3b884415ed8f79e0571387ec40ad4b6aa440f27fb4596948f8f4a7ee2e140f0f79fe8e5f83e090847eff613d2c07c74e7b2922c226a964477d6497a5dd04a425c5d9b1a9ede22ddc22c98ccdc8f1f3e59edb347ab461847590bcec7c6614a194809d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4212afedf0334e18be23698a9f322d7ee2fd17897aedadc32a61754e55309e190bbb56d281272966121e16b5a83836ff14a0f683c336dc5f951a4d8b83cd2cc988185c8372a60024ca3503b3a74a34cb031593a6b8a6cea974ca04e02202b819b7c56df90dd01d28b48c671ba9ef5976352bbe4df426aa11;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e1422f2a68ca65e419daa66883b6fa17d2c5267fd6f94cfdac29768be52fef9d592b725f1f539a92726296aa31cb459cc978825f28510a222206d2156adc97c25a20f28f1fcadd9af15f587c5c5d1d651ee223c51c7a49a989cd84cbd467fc708029d053ea5c901ff6ebf5657ee20e67b2e9a8260160d0f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf28c7667a7ef827ef77d102eeac7e65e7f73e9515a17a9bdadbc990e045b8b078d2145e8934508f4d7be76bad2ba6f6490d0a2036e730dd464196e3ef3a491b901e7d8b27827fa3b29debec26832236e61714b24edaced73b7b0b7783b1d1d59340a4db1caadd28befeff681ce26a7a99bb8ab3c29fe0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd62ae498579e5dd0cbe94836636d0d7053f9ce45b5ed0f8db2539ba4e063f93be698f732e217b71b61b75af25e86909c2f506edeff100cae5a615ad48854c9f47d07689c005ae4c724558066aa520637c983a467ad237c6b0937cc44ec21ef3566ee3ebc1b957287ed2d18d41474fe0de243f7387f686a9c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h726532be5a3159894d06595182ce5051a2e3fa02d74b36c0fd4a35c1eb31ab69e91feae59fad9c462d5d90e231928435f6c0f4b3b4d368a2ee1d18586f948724a4ef4d193592a817fb0df5ccbfcb579fa287008480f88e578a5322f3e2d4bf8ba936a14d809a9ee11026985102bb65dd646ef63976c3b20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edff90d044d648c8ff1bf2cc803170e5743d4a529dc1e7006acbe9b8895e1c2ea17846908be8e7f7a7e364c9cce5c66b8500867e422f661c6df7026b103df53a60efe294a243f3ac62b72bdef87571fbfe517297308ddf5eb2c189a8f85a89a523d685eb5ef3fe74f3894b08ccd7944bf23a67fcf1cad157;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fed22d4048113e6b89bc300eeb0e3e23f4b56796c6c3ac96b41cac0c0dace06ac0cfff3d33aa9aafa33c3610a7f994deff707061b80a076c33ba8ed67e3982cb13ae58065d98d14de0a2e278ed0f01a4e75ed9e396aee936eb5dd6d4af12b7ac6add57c0201c87fe9a8bfad4b41650c2ae5946eb5ba4b468;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1447bd4897394ad0c059a283db852be107549c967cd213cf523f3e2bd0e1a14a6f6a21c99d1972274802b5eeb02ee415d407d6af92141cf00c97833a320238f96d3a1be6ef1d11bb6fdb1b41a43a85d1bda79662faf840e5f43e28eecae6a009896815f92444049717f961ab949ab7421ddfc90772d8e31ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb09408d35a51837d6630ee35f7644870e42c130b97ba7366c5fcc24ce2fc9bda688b940392eaa6bb1a23805dfec7fabbca30aac08880ec11196ed8ca5e624aff17f3017965ae7c0acc04778ec59731abc13e276b59c5d786417575342deb49cfb7b290690d6e2c7cfc29e1731509e6c771269fb1c6b3d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c533c59aa3573f617de767c4763953033b4785d0bcbc509452a15f1575dc756cd283fa8d4f3cc4ce16cb443f1908052e2dd88dc533fe311b1aab0f1d0a2c92ebde2b6ba9af857ac9fb848851a0addfe617c1e43a8ece9b1680456c97565decc831e6ef23333160f3a391e643f325b023fda9dcdc1e7b3a15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f62460c4b0fa444ed761237aea24a7e96946edb97e77f4caa3b396f2207796025c1ae2b9e57ce22eea12f5bca35ac88faeafb9e501b41aad5a7620c5290c6cdec555a56d0ea4ca02f5f25d1db2e4b01c91076fbc8f4d1b7e2e1c28b1fd90bdf0b81a40a3c0357d3f512ec7c7947b44e26c3ed9ecd29a6d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14722a1f68ee0f267b2439b1376f92de61ebf0deea7ac4694356764ea50711f9894cf073bd5c5230726a20d4c03cd68c1af133e0f23c7ef8a7fb1680e0ec5f45a79cbc845d84de848b7fb4d128001d8abd47d54cd2ef054e364a536b7932dc090c6aed04b4ad7632f95e488237a6bbc2e481ac608032c22f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba64ac6346ca59154beed1742bc7f08febbab2926cee38912183b587d9da56dd8ab85bd823bffa4fdc039227a15cbe043917d9cef5c6aed56414c17e6754bd398bdff6a822ba7245b41c208d5705f30a7b8f9c58b154442b6e79d96b733c03d3920c3378af41ed2e7070da402c0f881ce57842d3cbcb0841;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b386e836468e7eb9106751803d78252540094e7930f0f526a959474db9806555e720efdb70a1bd239cb5b84d3e4ff702dea019d0fe74d345106fdd8510b69bf433d80e439ae0e981e5af5c254e822e004597b2b2694b7a9db7729f7586e876a709e9615150311b6577e2ba00652aba04ca5c3e98e36fac9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19fc6380163521b5c69db7559302e06f629e7534c60dfd10403dce2db5c0ee81874a9e319204e6ad175a63b5cb0ea7a2e796089eb9cc262e1b5c0c856c48984c5fe0b6356cfec8b6655f5384dfa1e33e5c92a6c8ccb556be04b2c64143978da17e44f7eaaee9229349c48019e2c02ef49d86386614a408231;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17defd5a88f7a0ee0778c78b439c32e5b32870e3c41d867813356a042e9874c80b3416e6e7a04f2fc5491c81b72b5a81d2b2e138df378ff94d888b78315dd036a5658012d349d65faba45c9aac9f004494274ab8102adc591cd0515cbd543a4c17c20c2afbcc67c3fd1dd85cdac980ad4941db82c0627be2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a47020bb9841b8635292a8fe6981794c4ca87e3b7b9b119c45b91a980ca5dd48b109d4f322401134d6c3bdcb7a9f159bad9dbf7fcf113dee24d0fca52c73571c08c03cc1ae4666b4cc1fa15468aeca40004f8f6eeac7366adbff618a441e558b84b55e9e7681c690cdc5b9d7e53f35101b4cea09ea151ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda7101aee7c1d731441d2d1725ac6830a5603cae6c7d09db485024e011b226651147270c42c4727a681914d34f395f7dcc3f3d278d6395d89ba9dacab1babac6cfec2dcee9d8cecfb5a0adcb375a7f4fbb5e8d28c9acb48b0fb5c5e002ed1f1847252821f97c999a511ea0866b6fd555db448fe1a8395730;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f048c282ddeb6511b21dacfa80f0ae15bb8109c7382f4a5e3892a4dcd535151d94b77adb3a4e4b3f3cb091002893faf467a9c62cca4290b051bb4634f87c9139a7eba73c19e949b935e2dbc6d58077e954d9a1dc6d8029baebff28b0c95f3aaf973194b7dc0d7f0bde78d9d62d69d4c107ea40e4fe5c6e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d7b689dd62cada82900d86878f7eea1885398a89ed3c09afff957bca07e29508085fe25fd78ad3dcf4a445ebccf30319f5894d9cded35d8c417b7f77bac2a96e65df825f3f38848dd24805fff20ce779e9a7bc122e3e5230a8995740e620a6d06557cde05d5384bf17f4217cf37c45db597177fdb6fa535;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11bae5a960ab8d84dffabdcca91a18972f6e0d9b906310e4eec29234e5cca3c35ced024c43164fcb92695767f7f9cdbc32c8951f424bf860b98f721581901da90b473be52904df64d91e6a8df96094189b64e316110f61ac64eefbcf54f355c5ec952c4d518078d7d716229b5097dabb9c8e07fbfc071a3c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194ffd96515bb2be68d014a04751753cc5df74efce40b7325f2a520ed97f188021ea5e55145516d859419a50c95520c37cf3e26cdfd81d4e56dca2cd29c74dbdb7bae463fffd149154bfd4d318295a2fac162a9f5db5cbfd2a671b86a39916622a6a22f61ee6bb588e93bd2c59714e61b6a2ffcb9752a3afd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ae4b29ae239d2545bb8ba4d54f5dc46f77f52c502cf5575410e52a2bec015934c62dad306a1e77b84d34fd62b3b6e74e8ca0ce0bbc5d500821a00932ce1d8522d37cee0e468b3e9e264850aec1322f3b20cd9edacade05ffb15c8fbdfba2e986cebbb834595378a61a2e179052253bfa332bab3fc9ff95;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9eadbb3cf7d8585abb0c1bac01b6373bfbe567b94d125879bb6dd41e28db927b6c6019ad4d5731f6a8cdd97437e14d1187ff7f214c4bedccb68a3b0f477427083d173a69b42c3e587b8953193fd9ae26bff2dfd7930338991063fc97b156b7db1a1414dd0085ec12ba9125a7bb2a3b851ddc2db212949ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbba8443f37fec68409f17e1d3f716868d1e3f6ffe3b308737bc9f40d9940f28f5914a81f26a8ac13804b1129af8d61f1eea2bc77f9fcb1ee1a397e7cef362585a30a819a0039f0531d25560279ab496dad30215a3776dcb4f4673f36c1dfb69c1c957c377d64335c164422ec4115ebb0eb2c8469e672887;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h237e1d4928bfb5d907c145b9181746a9b8714859412d510ed19909dacb60c3cbc0021f1c8b66a57e06a10d5abd2d2911b8453673b02ac173b26f2b1bd47305fef730e55bb2995b37eb3da2735cd666b19596f88535922ec231dc34161a6b4856863afeba46a1642deb11b735e0b45ff147009c769ec95106;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha0c0c2d234566f207ee622309e3784db24ae5874a6cb9fa4902aea295a8d9a7d5056f9f6c70a880489fc6bc6611a1e8c9d8fdcd3ef1f9769cf0e365862c793c9f97cfc56a6dc2f56dd0f5bca40941772988a1a6a0bc2892589028635b154883a8553eb70f3d447e93f4ff4fa10cc4415eaad0e83cc916df5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc0d6e61c14185cef6b0b91c190d8786089f71f84690a5dffeff50ec7e0b52eca1849567ada81ebaea7c95e9013737e8dd9ce58e6ce1e7161c81935aca976d98a958297c6abb7f5650ef3487e8f45544bd72aac6ea013a3a80a9c7d96ffad1e710e9760ab8d80b45fd77a74a554a52558c8c767a8c14512a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192828a32956ed3aee20667cacda095fcfa2b227b35a6ab11af91bfd223c97dde65185e7e90d143c7857011ae7d4ac78023556bceb142bd120de341868fd7af8533f193fa18234766dd41a453e780d083a40f4699066a4977568dc36193c58da33602a03a5ac72a05f299b0218b74d44bce9c87a8f679dd71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde50cde359a13e182f20de3aa16b8ee14cfb4afc1ae72547e7c513b3a4baf0a91b908adc08fd0f8e859a84365519d4f3d698358df7d1cfb532a9d120ad099395ff7d6c97d5637984876057a0e320ea5032e8d32ac84671077238a33b2bed07deccaf5a631392b75010fad7fb9718b93026fa03d5ab415530;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc3640b1e671108998a0fc77b922e9a8e3fc0ecfd69e48fcb9659e2fc870a9e2e2eadb073ff505c2886047ad62d75af1d45ab2c5c9624e5193ab1d569121d7dbd438ec43fce4cc58fa8d1114e373ae1d2c7fbcedaf0d8a0a83d42450c60d5decc0066c94f15705672481f1073d08c7fe15d793c95c2c66a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd90d94c48c771be397043341abc47c8fd84beb2cdfbc2892642d4028247e3b7f4ed67ff4ff3b1a8d01d4daf85009cd320dd89c1402f9746d0f8fc21302c2d17c8cac2819f71bfa3fb0f4df376176f49a07c4ce9e7e68007bbb06b0a615e76f00c589168065770776ba2d651d46d007d8eacbc431a8ed5147;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h128517d31c0c566f010a9c388bd4f59809b673a783bcaf80bb6fc19a9195d18f04407b985356b1f10b4b69d3456a03e93d16a8a018cb01af0d6817e38513b9fde73745b987aa3698eda0544d74b26c9b442d6e149ec03f8d6952766d0d4b0f4e59a9bc079b586679df32fbc6133499633751846b7171a5e13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c9eaae8d166d91196eb2d16828031afc01fb0b83525567e578cac8892d2a3c2bf85f727770fc5d90c1599afa7a9056e6d544cc2180a5160d3ed3e3ccb0357fa8634f590bd6f08bb4e6fc3a4ba7c5ad183cdb0750cf08509a609af3b62ddf9331a2df8b7bde1625d09d572c2194bfa4a8bc83cfd8fb63e0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3dae2b02773bc7c2baada033387457341b374c26fb171716a83c012e45f654c5c08aafd70eae269948a2a41f54491b053b1c7ac2a7feddc498f8e6d0a51a3984c7b211d8f771e8add407d568e369c6255c2e4e86d354316b22f4d9cb2277e5db32f019b17dd6bb17ab5e89dbd3c400f0d7d94a57e924e56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d62d51a03872e552409d4d7961adcf92c1bb69fc342c487890edb87f8737ea1757e1bd2e774b24a7ff109f9460018428423329211372169a3d1a2d32229fb026fd1ce40bb8622448e24c00750a715b951b4cc4ae4e12bc94317749183602681fecb9b9ba6415eeb6a6a719b58cc52d41cde981a608634eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ad1f3478ed2896942e271dc516bf52f9cf979607f573f74080be09e687f7abc29899c3dad213de9bc238ccf763d46cff9f743cf19ef9c722eda10232edc90808a0a2e204ada9d6f4cc8dbaf75fe474626ab9268cbf1d682be8de89f56db051473799233ad0cb06cdad0bc97d270aa725676c851aab8b3d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1093fe407c040153191964e6e4779c3a2c520987d585a4f8a827b72bfc35c634a7fbd6f5411d32f33948f2120344a642aa849f9721e5d28ad3cc2e766cd9a09abb764591c031f9144655eac13ab218d791bcd2a51acc4453084ff630c8fb73607903c4a74f2b20b22662c314c03e171d50bb492d38e2551b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a09f0be7a9fcc36ef45baf3a2515fb97aa6101661111280dcbd30ca3f430ba9cc575642dd8e42a780a368587112bc6434f720cbe4aacb7430c31f30987754572eb8b84761c1b454e816c1612a12826e62c3fd4659f260b485c4d20b543c814afa6123f7447064b6856cf0671e833618f4a6313f35c9cdc5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1234b7631b953c17cdaaf57be60f9fdc632076244b30ae34d8a861a882b67325fe658f58f6ffd02eae9a27f2461aab7a719fce5841b0441c9d1b4a8058eedb89efc18073fd00f40d0e9e7eb6526029e37461154be164116cc9dbe95cc953a79b683c514b475d4e7da65f2943ecb19783205632f52c30a7522;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heaabfd1a579a86ec94ade3739c92ecc770de55b18343d63e15f26428ad060c3112976da2e2159cc49c0ce9d081b9f4450c70c1fda0aad303768e1b29e0c69313bb2f057cac20038cf54f3639f4e66581877dfa14da1b4975cdcc12470a6c05be4b993fb8e003d1642aa78d672ce8cbd2fb7dbf907e70014e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eda640b16989b1071f407a7e82950b842d65ab96bf8f3fd3a620fc62cad33a7c834a341d8ee5df0dc469f8fb2ef47390df296dc7afb6e9bf4324cfa10dac928fdc2dfabf4707fa6c66d9bd5298e16dfcf0a93e96f556090a2528395659a96e0b214fec5cefb70c125d80a36ffdbfbfaf504dcc4c2ef5398f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1135cb6d716963fbd11ef5771bf2410ff414ee1ed1d05d6e3d8aec243dd049975524f9aa3949e522c3db2e048a19034f1b5a53ba7b8a008d3189ccbaaa92eb1da216d27ce7749e09d8b24304011cb2cb08d8301d154077cc3d67bfc690557a7898ae4b857160f74b4f89acd6687de9ae196891b127666d758;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2786eb2c4c1ffbb8e25af4824866b59116425c4cb10a816208617d3498b6e4893ab034bc1b1d84f858109a8e7aaf9e07d0ece9c82044d177a4f30e714a4060d079c1b052fbc1b42d51e508ddec11f45032ed3d8c0c9afeaea9bebc8e05a061d7d5db1506f9b59f7acc8f85e16f137c5cafca6fd7a9fbf4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be2010bcc4a693a5cd04a47034217dcdcbb075b4311cf4bdbc83f13024d33814d3401b824d4847529514b71ef3b142c5ad5c1224b701cd9a4111e66af5f5ce95ae6a31047b5ca740615bc9650e944410d5ca68157df7269e5bd8488d44630833637faf2f1f81f2605202b2612edb9f5af12fa4040ffd518;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176b5e6f6dcd7a6a492bf583330a5d91c54593901696ceffa5687e57dd9c03bb76a8cbb7f69010ea5621252070f6c071f0c6d087fe1da49a4cd62ce661ab522e348f7cc3b1df7e420da1c9f73434f1c1a614a67526816d63affe47b7d05e4fc2bf4df7143e033e764c5e1f85ac3163e72dee80bd291869bb0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5700ab701c1f248a268b2ac12daa8e02ac059178db65548df735ff93f34389f481308660981275a2770df25c19057945f2fdf3957ce37c741c64fef209726a0bac570879f9c2ab45d76f145d6567b349cca3c786188c35785deb48a35616c1d11930cc882b1430fe020be461c561ad4d0aec830dcb5a6ca3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f231fdedfc47af3c0c8c269a6f9b173ad13652b0133330014700d60fedd393237b7f9a6cb548dd2a0cb421afc4b0714abce4be8d25b854b50485e4c84ab654a94bf72862a32a4041d2a10316022fa4620a53e179acfb03a29de170d64991c0762b7dfac3498f32d21bc5b38074bd0307c1b7c61c652e057a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f922089e73631d2d1acb3604ccedc355b9985403b36ef35ccf483d7044fd4c4d709625a59d5575bb4c2c80fbf830dd1a1a311366b2ae35cde9d8ebeb7a0b5ded864a84eaf3a818eb65fa67cd9310c807c488e9cd601c2c446d6538b1b626b6712c9b20ce0e459a82a5a1cb174c519f0c9d521e397d627531;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d47e6b27f7142b15824099091029d3186062f6b7f2dd9400fd0083ce9ef3d53b54b2dc76843e1b7a2e785f02c4a34a2be62b2533adabecdeeea7315941a1e7855b102ee13fb235c557481da0bb68af0febfa750992057aa617e776672d470257aacb9b288c1174f702c6eac7109a931ee602dd4dec0b02f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12c6a711812957a6a532b0690d10bec77b9c65e4bb2495d4d4bfc10abcb99b3ed0a4a4d9bd7a385c48c27815c2a568c454085af12fead0a2644a9c85f77f8bc8746f29111a1d84146af8a27850693a7012c723b1185818b891fb20010cb5ebb0564d347cf927037b6f9f94cf32edb44032442660286953c62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd67de1f5967316d083b9e3f5e0fc5db0e820d45f61ebcea6e37751856c86d6f98b3afbf125731bd6dbe29015ee99dfe28fc94024a785b565568aa3b7a67b2e4559fb2d8675d11748837dc191f8c40c5cbcecf10fd57f0ad7c67e7d2fad9f92f7a040d4cbe67c833e3100a1f499849591f177c63a63d8214e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h886ae2be9f9d8319778b3e68f56eec87fe209d9d5fe474bf7ecebcd89488513838f05e06da6956e6c986903f66c78a031616949df8595d08c1470e01ca8460f82e37717b2c476743ca733df3510d68c8754d1f9fcacc5249daae6976c8f9713ffdafbae63c634ad5039f947a74f26866356aa6a8b152e938;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd41aa7314a0243b72d519801942ab40c6c6cd4df3722a0efa20f7783f20c8c6f16504eac4401b5425acfea8270a867b141e0476e55b31f91a8152045ad26d893ba12b59dfeeab3b94c4c8abc853d7768c2f2058bb305c381c239f0395346f2db0ff045dec25275ab7cfb97ad12ed59ae098976e312a2c12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132721470b0b8da570794f0a598184f51c5a809cd2713e113822613c669d47c48a12458057a9ffbaec994e64b61b5895720165e2e007c892fde3fe5dd305354095b78d00acc5c30eb49663be284fbc8d66954a62c8a13c654fd93ca90e22a2f03ea508f6fa3ac35f0f5ce9cd61b07f21b45a5190f3f3a1906;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14968ed75af88040f914e89dea1dcd1d7dbc4657385d5c15acb2c0cf766b0a27183b346abc940770d9ced5c2dc689e93ac3f6492d47fc3c416e1f97dbf155082feeb9d9d3f45392b3880818e9ef4a7eaf72c5b3a857ee95f30ca701b84664383329e451f58a03e18cf7562c3aa8845b0b8ed40edfb8f4ad60;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha08ffbab8997e7c87e2fb1ba2d4cc932638f07f95495a99eb83b408e8f51c5e702921e3e2cdb1c803e4735bb9b0c014e2af1c3f664817ec20d59907a5e21e7c976ffad4a1b5e60c15d22690f7d565be48da7c5820c5f0f387277268255128464bd00993c3cab05ef049369c78d8e4f7d338af5e68d82dbc0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8fd237f09647c9abd714672740aedf6ffd9cc14f0d2cca7b66c876ef39938586249f4ca7366f4c1038ce8560c7a6741fc98f085cb12a3dfae0226c7ed2dee6324aa65120354f58d7f50035003da5ea4bb531de1529b8e58e2c44f1f9c6e654503bf2042457789ffedceacc8e0ecc608f507b3f9acbb6a3f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h884eefde0fdacab8545d0b74a3c5eac915a5aedc2d4710f73d4060ed2ac23ca0033f2e51ae9a3cbdcc12db30ed527ccb5fa02b013636651214348e5be89e0056c65f74cf0bb11730ee83b5dc71c91f810be5e2059e36484821eb3aeeffbbf96444add4d611177879d76e69198a2fde0fd9a22bf96d190d2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dff182af49361ec266211010581379ae126d42403a6c31c9b510ef1083cf36a9048d8e60772a0d3e243620a427b47a6f1897780b39b6c4ca02d8f75f559afd6f124e57638bad9870fd6786a7229a5e443c8992c7421220f55f297b9e8b731dd7a8128c46063726180cf49ca9054030660a6b68ed84d6c1fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e9c178530240747107d3514deb45ac5618c497ba9c34f820f375bb4011f38d52d3aab57a42790c55fb01606205098d0cd75dc8f7a4c413cd5b5303d18179869572bbcce62cb4c21294d837a8cce459fe0d2c76258b0f285c29f39be4f655835fa6416bf5b10b3b80aa7d863aa2bdd0f630fd04f7403037;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f7a349f1bf4a4d0db9612690cf1a61ebdab245de217ca19a45f5ce542888ede323d7d08c860499647ff68aa1986162d89f32f0b6cd9059c74828828f54d2310d3b3749a73bc35f99ea06f54936b2d38a2b7a332a9d5a8c4d644a6c3f4c86d5dbc87ab5b87012c44204434aadbfc983ae18ca798efc263a9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e8f7f15fac754764276085f61bd66f2b76503b2437e6ca673e0212b425ab37dacc22e47e9f3f4a230b9ca364b116e6ef18041e053b6ede2e969134eeb74aa6952489d94b850c3f07e27c8e86a37006cd621e60822329cf5a58a3523e4c4c112eca607e11045a33c75a3e9136c50f7d21786f25e45dcfa3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h69eec218ab1f9e15b002cabf0ff49917913c7e733867546425cd320fd5915ba0d866c160ce7ed1034e9f20c29088dd59ec78a6ac642e877a434e4a6a5bdf1d63c0d9c8333743e68882b43823357fa4f2d49b844332822044d09158aefb8f8e2bd4b6597c866a2b94f8ad17636630d9d3c9dc40471b4b61d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd74d00c2a52de98cc460f427d4c220cb4e587b68175d80106c9110fe26ac9fab15a055f33ed586112cb37372390273a83fc89e28009fca5bd76d5637bbe644a170d78cf6b9cb2e420e47a23d5b2e8f70724532beb79315dc833d3b2344b96aa78d24083fef3695608ec82ece1ed9696314f032a1a0170cf2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd2fd1f1f89ba17b39cfde27a89aca2ce260e0c468f29d4b3d7e87a461fee83b96f9adb823908cf9887a5ce6b557915f32fa4646ccc1983df69d454fc5911e22d85495b484975fb5be1dd7431d1fa1e4fe71f229c1a870871e53e49d529e547c078e84ab3d4fee926e8b8a84a9beea27b1deb1cb7c37a1bdf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9e5d7602efadf04750be34dd7a2436c11f4466acb68f5b360e347cefaed12da5fc7ac4295dea89a6f425db4fa95a790b7ae76a44569293881da97427b0d987355c1b68f8c49f062a0144deba36c8b13b7c34e5bdae95d89b94b3f75effead2a628f0e7dc868499649c75a6df76f21dbc81e65a1c35961e2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd234d79635af07e14eafa970f9d7b815d5c06f1641c2bc5115f1451622b69e64109efc67f294e841d5dae32ffcd309a92a4b43ba1e4455c2cad0faddb473d9268f3718f6a13995bb7a51851fe59acbc3e226a8d8079deef6ca1224ec18e6ed8c3710fb2e8a3ecdcaca74a59054b455875113b7a737f4e26f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c099852661d62df5f751766d6346833476d380349e70f6e7879c6ee3cddce3fee61427763e34eb60f387821d5f08d4c55497f2415a0a5b6622f93c2223674c6f62acb58bfa148ee12e002659a0a2a2f96a0af2e3a9cc6af52940e3155e9d6010fc17d393ec8cfe9b6a3d76ded5cfbca9e37e3e721dc6ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab59d27b292f87f3774bc93f0e2688110886e847dd4ba6290d9de7e926c4b7d3c3200033c825aae5e1e00f914836fcd9a065b7c3bcb54b2fd4a6f2a112e03a78d183e663444a4572f8ef5c22eddd1dae3914d6a55c0269fb65ba266e453185c47ec557a33a29da4289e44644ce16470a895b6a1d937d8ed9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4d0acc9672b0e5d079d901bbf69b2c4be42a7a8870a991fa3c604e9c5942cb5161152aef9167dbb23e474e279e048fe79239770ee3d556bcf61ddb8d769a656955636f01a1b4bb69f7a9ae45da857eb77281b0d39417a48fe1efb141eae180838fe2d3f92f05ffa19d548c192eb910b460e9f94d4523728;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hace4fcee193b4b30e3636647ea8ef0e45ea69361417156fa8f47e3cfcc547640da16c985109ffd6b896cddc60065cbab15ef54995cc9796e3a92708a118fd70d00af9a3fce197a7888d48a13d932a107d84b5fb5ab8fd67894005c130d1b3bbe29de53c80ef6ff4a08e7bb6a50c3e13e9944d5c147731cbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a77c56c87ba4e113e1f5bc06f121ba5e5f920aee9827ef92e12075a41bfa5a377ef5e39fd182a3df3899e130e63ba84fa38ca2196f744fcd01efe402c1c1c4208ca33ec0b25323926467acec696e3bb51fd3eb429c21ba8081a9f020fb81c68228acc0952f950b503e4f9903e1765a9e05a8bf2c68cc4e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1215f2b43770fd33cfcda506497eaa971151ff55bbf75ef3fb6e38bb5aa7091bf6878d14db862f7b2a003347aa59730fa5237d87cab5440c7f34eddafe298f79df7de234b13cb085f7d67c27c7b7bcf60f8a1ec849f0bb1eb9648e43550ec3042ef0ebd196a38ed1ad0c0e0f3a7672749593dcf8676e91a78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193312dc0170e51ba013b024fdaf110c5eb6cb856184f45489680fea8f61709ad3c74189eca9da3dc42b13927cb762b317a755cb12c65b5545317eeeb29cd9100ab4e7b668f6c218ac81160d677e8840b4b4319218eb43199971b38e08844fd60385ea60d23293405daabf5d353deceaf334de59e3fce86c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d7fa25b666d2a248f9eaf7d977219a5393dc38f73bb8a5738c08deee7dabe214b6a3d80a9cd5dcfe00dd61ccd540e4fcde3c9b7b9edcaed089ff1d34e717f3ea9e8d714d876371f0eca69a149fe4395b176d4392bb5d813f442184201dd3c0485e569cf06db6c4754b5c35d885e33435e8fb529e44a89df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187b623a06d7d5714571ba45e3516acbafbfd72da228b181bb778484e716c19105a6c65b9af630ed62b5453665dd327b07bd5b6721c6010955b9573e240d079f874d079cb8c743d8aeea0a73e26ae6a2da02bb6459431f0b388cd6bca06a04eda7c6455f8c9c356e9dc9256c86763a2fb0a690d5d778e4640;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9fd6fd84b217b59c2a6ea8108f858ad58540ffe17f10f3e3756c259fdc81f3ea105e4b0d3c1a8792d51d0ad4a6bd13907d334ac3754efb862c202a9353045611f14a2c028f037ac38b8042039863edd3169c36c0e0da32665e501c7c05676415d796bb223dc6a2236d9b266b6bf75d4053d353b4f2b6ba8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f96f7d1b40f6556ae05916f9b3822acc432702183e8c86e18343e2f6a0580accc527062d1538499c39caf797c0f22ae87126dc4dc81157e7b8661e11c6bfa2b4b8d351efce30e702fd4675de4c16e0ee8c824ab80d6e8b4fc479da38d4f2f8fa96c9629b43e0010aa4d056cf751a15218acc6506d7e95977;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h196ba5842676c67904b39312dcef5732602aa6b108cc43792eccc1814f8b487fc4b31a7c1c1a5daa079e1078520a17e6e59b148cfbf0e2f2232667734f86bd03dd4e307b87a15a208d2403b9f6a963f15639baafc6bd80225485aabf011dd0c28901bfae0f7edf238f6b8f271e6e3a86cd801994eb8124ef0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb485f8a1edd8cc66c61fafc68c6bac8bad116a79575ae49255c8364c4db1719035e34c310c39df26f70fef1c1bd02f6c8eb718c7ac1b9c0fc67d1b80b8bec1ff0e85cc633487fc7b3edda80ba7a242be5c20447667e18d091ec14d19c418aa58e7bb458d25bccc7bb9a0f8d1068ea98db3e0117048b9edda;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha063f4b31e8fb76f0f10802f8e726202cae5e0b3a480093f1966888f6701df10b0d8472f961fd7911d12b76678162870d53ab60c03b916f42257f445bbd9705b7b8cee164646b52296b9c5df7d3e63ddc1179aafebba27bfe67bf004933f4f78562746177ceb683b071a3bd858f77ee29029c4422c28623e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10ea06842bb8fca824d8778e8dac0d89a809c86bd9be943c71803089a9e7a6087ef4ae2760bff3011c18e5cf0b189e4b56519dfa85f2be19d9f354d50c5494ab105ff17c8c5df9b6730c53025047b6df786df809e409f1a51ae21e1ff28fa11260da977cd7591ede635b46e10317493b4d41a4b2b541da3bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12fda6b5dc331621bc1a488d532e6b981040bab5d554025cbda227406afaef95c07914c1613b1add4737adeb66eeedbf88df3ebdd755fa48cf2680bb8ffb08af1ad7b1eb034245efca906f41489fad345fa099b84dc7f1540515232b8ae4b785dce8d5bc1368902bb1838a4f5f0b54086adaac147c457c87a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa67ca5dc7fc6a186acc621cb2f01fb21cb7022fb87c1159b9acbfdfd1d545c029d69cf49cdb71110d6071a259345a7d89d23439364568a1f82a91dd400b93ae010ea313897f362e6554caf7a72393f77a3d9492a147e5c9cfcedf8e1f8b7e25e4ae2b7574ab49c44dbcd9d7b3314cfe225e75b6531d0cfd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18b635f7b96f899696e5cf590aff6643971fea474ff7b4e467d20b1be172af5dc0c4a0411621e0e8ea7be41be2d06be6e8cce0daade951c283919474df747b0652b5accd70a817336f3bf057dde68da34fac424beac1af3550914259183417ee8f3eee0229af3b45c859485a66d20986074a2e0df5b4ff95d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15290ce30d261bb126e4d10184c4fdaf03eeb1c0f59606dfef5f9d1c490031282f9899a99b0beade3f32353a9308aa9396446d52be515daa778a77eda06c69ad293e823919beef34a068db755ac5f331a047a3918994864e6939824efdbd328e62bee70b551710ea38835bf9444802c2d57e926c05543c081;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h180c04d22c669613999d51d9e0b8a99604e111a1627526a391a41177bc7b5e068d40e999e333f4390d0c5d30a4a70e508bad044ff6bddfd2df56440388718da8483a52e9ba90399e3c7a39d0049fdcdf036cff0f2156c9d6b8633d0de5abd6d78879f6a9c0b13a347e911282c4d47601540079e89721b5d9c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1272e760e5e5e01bccd33a11d51dd278f3accd3017cf238c8d1e191662eab7fc24d0c6983d68a5a1eedb32ebecb53f946e11a44948e09a0b3e6fb216b96a41a8c4b955d572bd794204b1bc8f86c45fb97ed5fcd890bd25f6f06f3302e32db28b5c632e4acaa5c56ebb2eaac7970ffefc38ce0582bb37d782a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1567d3ed57532faed26f34b2c7c530d3a8b0d8886788310a3aca29543dc03ab3783f271659986eb0bc9cbd583181e254ace798b001fba6d6ea6beb0b49d31f4d561291f9fcd13b418c71ee8bcdf9e490a6cd55c353c67a9e23db0a5e8a8212c06b4698ee91b2484f132ac4215817a2851a000bc9a6eb5ce80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19205a3406e48eae338a386cebc158cd6bad4d525299f8440e3efc9343a7d988352ecf0c88119d36d11f3a63601bd0510717a480fef6ac7b41abc265c8100b5e5ed158529b47663e3d0d0da395530655b4732152b4291c821d259e8a516712770a47951af12b7aa67c7be3884517ee997cfa261748edca1e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a6e4e6098bcbbd153d9cb7f064249eddc77056caf389dc3322ddc933c3ea504ee67368f0222a23f725529bcd2bce504bd91581439c8e2face508d01c5d1c3137203a936097189c16baf065d2ec5299e0d02407e59b20e962cfa51732e4d9d7905fe7326743f32327ec3b966ae20990fbdbb3d057237ef1d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae784fe7410c2b99fbfa7a8b708cfff5ffd4ffd92e4008ed4b98266e784965e19a575a6b43987e77edf712f0fc99fc5b0569a836c721a0a71ade0969aa571673683de1d3103f783f23639f33f3ef44c200a9f2eec339c9fa39bd3fce52ffe1f221e6b35fb3995ad939a9ab644f9ea06fac067bcf3f600705;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e52fde4e1c203ebb16f0b16bd3916f2899a704bb0bfd13df39ef4c9c721f02e891d939489145456701a28b0239abc9ce1d8e7d466aa25d7ef009cf633150bbafb7c73e53e62f29b611e92c0e37b8dab56fb0078827143b8927c73590152e8a1d07dfb27694296f6b2b17a895fcf478209fdee449e5bd8237;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1afde4ebefd8badebe0952ce6fbc8a9fb5f70eb5005c45b66c8c90148cfeb00078681fc4b444221225415a61a3727c544d52bcbe9b1ca4c96df0c9859609b6e867ed587605eb2840f14a8fc97c3515b48a1407a665ca6d6f0d45e5b67c57421ca1c1a71006c98ed2a86405887ebd63085ccf00ad4705dd362;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac46432eda77183ae1078caae928084eb6494c75850bad8657dd2edd26baa29afc9e5657140a8e445b28954ea8843b6f35d7360fee325dbe70957bc5826cc93e5a9d7e894d6a1d9ea76c849374143bda7a3988fa46f44de99797fea536099b578386d405994d97bbf96fdd82e9b63aeb8cb464fac78a805f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13830a42aa30b4233057074fcaceed0af8fbe51ba9ea2780f633d1d1e536e6883278e7816f82e553ea85fd91ce9ff070ed81e7935c1fa8673b25c9fb3f0b8b25810496b029b306cca65e5115ef24887ecf0027aa6f68cdde7caa3d8ad370dd05f27a512a07441d5e42da70b7ee5537a7beef90769076a31aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d341c7d2b98520645247b5f84fa567f1406e68121bad6fbfddb39a1cc0ae5c8add4322239226ca2cb91b85561c8a702d73074515cead759e748cd9c10b68ea76a6657a50220c4726719339401e807e2756533373fe0d8edc9d0b8a27efb2d2356f082801f559bdeaa2492298bc77e7c58002ade2126433cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dfb70db9ac0a9dc7c0f7431f9d5656b497cc3287054b319e19c4c662b923b188da9e75b1684d995b16f395a2270f912821591497184f6c370f59446066dec7c31c38d231cc457d1ca41f55d447ee3caa85fe40e87103d7e2faff97b35973fd4e9bca02f8f1881ee4e75f43164bfb5f4900c42c6883e38df0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aeeeb21d98d702bcf9a7d02b6f9d03985421fe573827de97b809cd466bd4ab0bf5163cc9d58cf9b27ed9d541ca2166d0602f1a4aa89330f317c610c46b6851a3933b19b0e1d1784b782d605f5ed5cbec0d09bf8468ec513af10d23773f554087711a55e3fae912b1457ee391b49b0a6ad0db1456dfe48889;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113f262843b3bc890ab1b7f46433834bab058e9c2a4c0cdf55f77252db9d80b924f94eaad07772deb6196f680fa26fbf770deb1a537a550659eea097492a8a0941604379b0dd4cd1c39ab23b0ac0f66f73e5a6ebeb8bcfa43447f036589e019246355a52d89f37472d56b7f37e046f4d62cdd5ede58e32fb7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h783a7f4157319eb7c3e29f1ed6375efcf5462a476c9440758ef3c180bb1d4fe3b04f306b0978720d0289f549d3be359026556b727550750c3b6ab5d782cdfd7300d15f7b989d4400b1069fca1fe401c3658403262aa13ae753c1774b7f36a1f941d9d2fccd82e903b8e7f462fe1e26b5eb012a1f01694aff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109de00b8687ab92d36db3c284930dcae234f2676720b0d0875efc57b6bebe863f2e689c0200971de4c50cbac6c8a51c66ebd482b1565571ea0cf2485b9903f97f4fd241a9dfda5cda411718e1d42dbc117d2b7fc87c1b7e5dc07c6c45a63067c2689ea0dc9e3cedd140f5efa6ecfb4372764e621f08e492e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a24fd8b0fb6a9405f8d738abc21fa24f7e2f7c6d607935f095edf66c13aefd179ab79058ab712ba70316ac41300584b7d72e025eb0473ccbd43edfa23fb4a296e3b252e7f01b4b2a1bdf3a37e84d1aa6150f0f5daebffe93b8bc06f22173dea73a3f95dca7ee7f8e8b9aa504a59431db3a6959be534369a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h211d2c8e10fab91e48680c03b33bab9b723046b8269e82d192bc9da1c3c58750caf0c880ed73b0d091fa5a07f4a6aa40b88e3f22ac2f1dd1ebcf9f28cf64afc6760182cec4dc352e4935664126979390096e2ada7be26c93412d95839ca6e1aee2f8f04756251cf3b157d9beb672d4788880d2f049314eb7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h473662c5b8eb98ca470b502a3ff4ab9f5944f33b4b346dc99a8093bc45e5e9b957490e1a732b3547e97fdf6418b3d1c7f25fdb63bc0f55f0e901fdf7ed5f937be44f96095c7002424878f34fb133bb7d734576ff78215e901e752447c992dc54cce4e454d02fa46c44dcfddf67a9c269cf172aa47a10b9c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78ed43371c2cd18f414032ab40b34955818cf33ef6761c366c41e46047e9d38ec122dbcbe154d4862914eb968c33d912bff1a768557af91b2c32efa8d2a2051849a187916633b9d5776190068985068e468233b59b021e8c470fc8f6e22385142455decf9f9ab8fe9a95789c46a4960fa2a1c8cee157387a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8c3d58531b886b36f3919441e003e85ebc350f18de42a7b075eaa7d3ed3233273148c47838ddf478ec341e95c7d76f6fa3b6788c1b5e5073c6fcc867b849afcffd28d8460c88b19a79e57d594ff949e44d73ae23b13dbcb41938579a72a1c103f80c3c52ab043c1ab0d4b1d9741f181f8ffb82225612d72e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1079db21d9a6b68d06cbbb975e495d95705ee8e8c7d16e6e07499dab2381b935ab3cb6f4f82d904d3f02a6ecde3728f6c8c8929187d9c2a6844ac28180c1372e4b814dbd1f6051bffe4f7a8cff5cbb5cb080607279e71a8b3ffd21d33fde9a7a6c7b2e69f984aaf6b3fd89f6b1a9a5db51e98173d0e0f82a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha8f37afe50c74029f54b73c0f38902d88a0a5ad571c5d05610d6efc2387b0386fea2df0568bd133e33f9dac2cde0bdbb61ad498b08743e3b115a80347a41f11729225101a23c534e10549025bcc41df6769c935aae1511be15247c9e915e753957a05dea01d195592b6d14bbf57bdd80b5c0d1d82827f74c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138d54cf144c7f6219b8967cbb4762363f85ce3a260f8cbc51ee26e3020058624f6d2029cc9573e3b5bb4299a37c774966224c0875eeb69195f07f794f04f3ba424e418f517b7c1b0a42727f0341172c3ed4ca3da097e3f62152dd2831750552863047481b36bede12e87806fffe25185426b0aad1c5659b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ba5384be7fe708f5f58f1dc3751fe08be29bda0d6264db9a25c5400004709d23803521fe1df856db18a5edb422473dcd3012a8bf5e7fd5fcb5bbabac327c47f0c7c4509bc3587c8c99ce08d527696c30197d439dad47681d3aa36a8435d17a04126db1220290d2c2f8c4adfd63ba504dd5e9ae4ca676260;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a39dc0e27dda44168858cd672a2c3e4b5200ffa2e8ac02d49289488a6bd495c7c788757c2da681a8af1a76349b70f0f763a02cfd40c894d87da9e02295fd7df3efa61c65fdc53f726470341e80ee2f998ef9568fb99847fa0ab100fd8939225055d4459d0d0898e0bc53ec34b545546dfc0c5ee712822cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e7e4de0cf7b3dd66209733fe11d8c87731932002affce1718deb1a1efbf6959cfac1c6ebb9a421d265a26483748200bb97d20ec3b007716a904747cc9fac9009820882c91fbd3090ccaa73fdfb2979bed9d9922ab0b09a3aa5f7272dc6d07b347e8dccc93d79bf3ae20d51bb5d3121a1fe5f5bc5951b103;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h853ba1141c5e01b06591c1145fbb80ffd8d678ccef1344df76ff5c5aada10c0838f796977a4be20425ca5f13582f518d9b339511ceca6eb853867605f0f25c6865f83e645f355322bb5b09a0fdc66c56e9a97852daa97f109e443a6dfafa2803a8c31f9030cc05b0c857d6151a223d8f9a19121f98654feb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a22eb55cbabbc2a8aaf185305991a2ed0fd475752480c90dbc2fa050d06158021c7d641b6164b94c960d395d2955afa34c0d774d7e540a36aa1c2318d9d563df83f525461c78d3b705687e927c14686497a0a76c50255c80560a3f306ff2eb7cc904fec97c08c534cd5001553b1f8ee212ac206f449045cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8828c35e1aac91c9884ef3130483edc90011998915f80021debefcc5d0e7b099decb096d4d2cc73006d37b072c6306f2e9f2568cbf19572d2042a66bbd7344412339647ffe959000fd1a0743e22f0590947360fb96081194abf5c19c8f831a681ecf4cc7744801022dd44170d5a6fe79bef6e5d754b1e5db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7b2d2e2db72e141a65cd50628644b5a72e6044978331ee20a79e4afa8db22889b0e97b19b967062f644e2453fb213dcefa4be8315f9cab276afb6d1b1713892104aad191f8707a54f16acfa7730960d92f645490ab662d615b01c66ae7f1150413841d33abee5b83d4decd45b82f0b5c1e519d0a6d66ed9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5aa18968ed52ea4df717aea93d32570fa21d5391a879aaeb8ed0dde2dcbe5561ab49caf8961bf49bdd91c73f95201f63c42694fae1cfb1258fefb393d065d0ba3a9ff4f130320f0ef95c2764faa6b236b029bfd4c6fe5a052cad1ad448ea1b1f50bce315d7a34f7b14bb7eb077988d2b471d501b3a4a12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h141fc909fe59fb92db68b83ceaa15296661d3ccf2f792f7ecec275ee8013e9593d136db1dd9952953e28158bf5d5d33e2e6d242e976048502872024da3872ad70d9048f4fdbaa412fbec183022a45041203a5fa36db807c1cfbd6aa3a813d49d4a88d8a195a0f7a1230021c58fa14b73d1af0f247ce152bc4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47294466cf9803834e823006765d129c1a22197619fc6e3194111e88de450c316d687c3ada0c2e138428d071a11abd45ea4b7f23f7e112519fb2aeb578c69d51c6b0d5fe7dbd5ab08cc563c88af6d057f4ddba6eccb2a4d121fa48e0b6159b765016f49a2dbce3906d27406480358d95f2c825435b0256bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8e96500e3cee55624be69149ea8d3edda6649c279bf816e5b4b25d48afe17e7a39e067b50ea201e51634976b3b891a381713bc4138bcdef31be4d99aea74402740c7f6283fc3984170dd43985c377bda6501c5d1755f5ec6ef947cfed9587fbc0d9e15340709388d0e85010167423eaf8f17c2f613cd4c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe4149b4030942842f48b54e99e4ff9909ed86dbe3f13361b982ecacb0a4d148c35bad92b55f78af80f87fa8b47d6947476062b1d4153f1b37b42017ee3e116a425793af59dc365efb00245eb59fcf86b63323e8ad9abb21bedd029ad2e8158471fcfe84379c6078b75d976587ce69348ca5190228d3711;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b7fb3d36e30fd26979b1802ff905ba57e50554a2b2689505c0d43188fa9a5e5a903bf2ee02871d9b7bf211b8c8e5e4072ef22dc95dc241415cf7247a6523800ec68b10917551d7ef38000e61bcec50d8759269009667f8d4858b4b967ceee14f9c7c322165cd6962fedcb08bc8f0d738320f3460a93cc2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195773fc32c8014a96995ba754a55a6ed77f8d35c5b4484210179b7d2c3c754448fa09850d651b7b98412b5decf75a41a3bad6a47b012c7db4d6e08d68bf0551f2f285bc199d402d1d1c208d690979ad372ff387d25c9a1a88193c8785f1f4e5ae42a78d13a28ae9cafd61a793fc51ddd8d2296e30b8b99ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h481b8d3efbad300e43146ca62f764dd8189103ce92616de3641a4b7fada5baef1d6d79ed576a769daa9ac75dbc6adeec48510d3e383f02f399422adba239ca0a38537166994051c2b7e044cacc9650dcea7aa23bec8012fe01c6b9f04c0e9cac6ff9eaed64c44dbfe9d1a94d3122c8fd8e4f62e2a0671893;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h380d8fd2d91de7b1b260a24a6848a41f2e156db7ec85de80a36fb65f22201aa1ee8bfd3e910aee75707ad348877a456db530e6fa14e247cab3bc10ec1a37509044193f01d9a9b923df1367cfb6bf89fb6b6c56b2c8d7caa4d76236596f56771b6abb53fcb37ea4b69ad724075c88a2f61227506ab3dcd9fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f858b1c4f57badb62c9dc25686f3c15c103cd2d83632db530beb7100df576f6618c7f502a5fedc130eddc1223913085f14ba285724951e74e6ed8d8d4d3f07e010afa3a2544dee157f92c5e3aec6473aa6acfeaf8020549cbfe5f5697bd6e7fd12e593d4a29712b4c1f9490048184758016278888a34aea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf23b740d12748c5abd1c4d027c5e9b489b6974cd0e8ff2c786c2c0a6f3bd87549c44263a61e3521097d5869499565947d20d1d331925d70127d2df09844cee2d0b3c94003479733e8f25b82db06875e5ff93c31cec49cb080435acc58dce9897c0c79bd2a379861c2d87e50d844f4e2bdb17c1970a4a862b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3e0896235381989d12647dd732fcf6f71476c4cca52d4297669486be0fa800fd1288a29d5244c85201ad30c4aa66703160707e7044e6fb0a9bb4a5f6cb07dfdd1d467a5cdf4ba32214f9096366aa45c982090e852d663a58d382c8c72fdd9e5cfa614b23c281d3cdc210a07fee6016c33e64de6a99e82ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19975b44eecd2895350ce81654445fe35cb8a751036dd4e334bfe7a5013f4c965f5a7861fe9d96d19bd34fbe02103e2f00204bfdb13af6c18df79496d823c436afaaed796f7136b9029319693357c9a3c05dee08582535abe173501fc02d262ca7ad9a6fb540d0e20d75b6fc32b530b22101076ccbfd6aa84;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6f3f15cdf60897daa9982f555e33d0320c4e312681dc607356b17642e7e8d9887672b5b77aba7f6f2f9a209e1b74d3b32e3aaf38ca89bf9ff901fd5d1fb1f548a16c8d045b052ab37b1d6574d72c66604ed1a3ccb875b15f87e5387d0ea0b1a06622857bc3cf859af93acc764cd83b4b6db755bffce0838;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3754fefe86f5e0a8497e9194b11d8cee27b120761053bec8e27c000bc75c27f828175883fc2f7963d64ab3bbbe84ba0ba460eca8ac9a8f48fc9445d8a187c98d2981371662345bc4fffdf6d5b81ab25d229081414f3bf04db450984ef4df563ef9481855b5621a3113606c8379174ba19b70ddfdf69adc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f65d54c23a72aa04f18ba03e36071b2507a3e322cdeb589c175b64609a38e01eb95a9c71fe087ac27bee2387de6341ccc355f91276377d330a0c0704fe5b29ee427cab190c5f79fcabfd1cb90718d4198e3de26ad197f826ce5833bec261b4af47a8b7c5b0f18605be5a624d346fd4b70483f6ca4377c07;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e40a8ccd2a3654abc915bcb976f2149be128a61aac0d948e250d7c9e0ba6713c54ec62fff8e1433d85ec70ea57ddebeb5bf67046c88d56e1d5b3a53027ae4ccd55b1ac063c3d9804a141e34b48551ef8c33173d8f48f0100d8aa4d90e7f222f760499e1b39468fd69e55db1bf2443d342d230d05bdd31af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b60931a319ee3a99055f726a1052a543d5945346c3d01f9f60f3f80e4f2d15f45dd85a6661282a1c0acde4a889b07547769c63ae8a9d88601b912f3a3b91d22750f789b9e4a1ff45efe7af65f270445c1b7234afa95181c7b13fc76cd55ed3699ce736c5d9ab922d70ca49e5119f7e71094fdd36a6dd434;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f56bdf5b24f66f5a1a70506dbd77c8694dd3e92265610195be4714d6f2fb88b610fd1aacfe34928518193801cb8bb933acf34edd4ba18a75f50f2fda9f06513d3c15bc981271c059d884dbf31088adb1b70a6f77f6b4b73fb6b8bb8ad4d26dc89e76518086735c2b6de4972fed9dc22dfadcc6ad99aa629;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f5c6a558d52575f216549a9b4cd7315da70e5fb1ed2a7b4fe08c2298e5b3aa7fd5b64bfe96a4c24a305995c4e59f39f3e2cd88767ee0556400a19a949a670f01cf554e746fc4180b43946b4f3d52783cb0af32585561570a16fdc893880047e5add71bdc2698918e148b3cca5dccc1cc4249ab25dde3292b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c56cad637217bb2b7ccbd21c746083514eaf9ba7739fd5d51a44481d6c17615beecaa3df47494057ee417b2a1bfaf14d09b4b07075f16798655418272486b370ffa6fe0b2a010166b78f27591737f6237aa1e260c67c0b93acae6e474cf69615c12e6ad68248fe5afa8f7023062844ff21fac32a81de83c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eeb1aefc7e4da7ea952482436364709a73318cd0e13cbf1f8f45eb4b57b14e54e16b001ce82f81314c7303dc25d5458db1b08f8947912f5acb77efa9d7fccec2f3027fff69d0f69bae26ff37924666b27d1909f926def3e93995c415188bfca851aeac6de4cafcca909ea764ce6d6d92cddbced7eee4fd38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c26a9f7a8cecc041e5df18a6175bde33fdad55a68181cd52e56ae4e10e01961abc7bdc8b745245c5b887bc5329d30e55addfea9ec7375d568c33589f884c95fff8eb755b50d098ef58bdaec8de2f4654ab643781974ca306e9fe45405f02f58c71380f8cb23f6c81089bfc7d2e4bcb2eb0c304b01ec4e1e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfed098c49fc8af2e40e7e47f33c59f0b94a99069e21db74f39c25fc240544f6cb877d1e34affe677510cf84b056922e30db02f3da7d3977ebe5ba46b820d53d759a07e6765a5bab3c2a9db4ee222a8f603fdb04c4bd452455dc836be7e014d188208a23f3b9e929a64f3a76a3b5290a6baa8d8584360288a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17508cf396c963ad6b8e4bf3069251431480c523b461e39195e7035439b47e2d1eeacd66af5ca235805ad9ed10fa51e510f0f9189fc836f47ecf19c735043fee9f0a7a8c6984673bce5c568312474ee33e7d0348400f83fd8efc7d0a4d0161871dad13e8bc66f3eb65def8cc03b1b1f7ed31ec2b7421323d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1172fefa2b88a5d98dc1805f60e5c51439da2c373e8feee69f8f45baa7afe899ac50c8419ff0c8bee7c6e9618c0b11f5438931fd90f94e916e106b0c540bfc014080f56d394ff1eae0794cf708ab577f4ceaa860d53948ecdcf829acfaf154b787567faf2cf1f4f4694eaf365849dfffeb87d50c5f72623a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4a23dc8199d75bee7885acef102d70f2fb228e989fa00d34e4e3157e886282bd4fc52870ff8b6dfeca7db11a1833668752dcc2df165fbd785c461d3b24291dcaa242f9c71fc7b9c220bca69f2a307e5939552799b719071a4d63f656210c7ae8fe6dbd5b4ce4cd04a86819ae5a7ee17a6f91e41e0b57c68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b44b5b1cd3d674eed6815d2cc494eb47253f586548f41edc9a6608178eb7f35a038ee6b2c599744ef0ab906275d20f2c66b6ceb07aeed6b6015641bfe3230d848d43f67e7c0d646e2e8457bb8c28c0772f4c12182a756f418d8114b60f6dff515bed70a26d4d074163f47bec11e526e5862d54a2c1c459c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20710e164f0402ba9f9f3dd32e9945bcb191305262fb99e98872bfe7df6d44ad1d936361bfff020a5f8d1b885f1fb4b940f05cabe81ea7a6c77e5b497e57672946278aaae083d05f7ecd1af7823f9dcf524453252d4557e5f2e9ac7ce5f4bffcf0f3b9ce810a4841e53a016888c04cc3c7246a50b712010b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha784dcd7b4071e6f59bca004b952236aaf6d5d2b9015752fe34dec60d968f8a9b5635a76e388fef5e946c57a6b6d27969b01269c8d1d036fcd4c54af5ff9c3cd947287e4c01317525c4f27e2973ef72eb2edf492ae029a3897dbf58a19ea6e1a661ebbc8f534e902180790ee439010020b18d4f40b516ac4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190c72b05daa163f8d758dbfd86c684c24770a8e79917a98c8f70a08ba530773d7adef376904ca4f78f0a8cfdf896305e5b57e49e0f81fd31548a051702bb9a7acc261d1d126ced2a1053cc938573cdd1ac6592648e9b3cc1d62aed3efad8b185db90b453a0956fc853e67b68fd03545b9549b2649ccce162;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129e1fbc38df9f10bd7a027390aeed415f095c67ce65b06ad21fb21a3928d926557263a8a9fe306946b126e54da9a6adf415ca8aa3e36c53a4da7b21a848d97a4e3111c773c669d69b74ce53de4343e077ff23cec5a80590f0e64e32b58ac9da0f5966fbac1b712136d97d75fbcf9637865db764d1387db0c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182400830e39393987e03790533f74694482e674511b2e66ccc678b85e07e731bc6b39015aaeaa5e4188949488f9d06aaac31d03a479c3ea1bfd4921975ec6b884f1c85fcbf384a5a8affc9412b0af83dd5a54a56d34c00e57304ca9c053d0d848e245b47f1a64df0ea395144df33c3e0069eaccf26b75806;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfad7ce80f3890903bc352c1be551258d29e433933f91d468e541c74fb1e03a35f36910c306d8fea0b084f0cdbc32aa8e559b073550f51e27c07b2b3aa5e5603ea25afd7a016c913e1c5612dc2f89cdc285a582447abd8736170326287bec0ec84c7cafc74a70a74b7be5e19931f7ae030074b2669562c16b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5137eb8aa200a5603824b57f8dfb676a3c8e1848e13864b7e96a78bb0c2212423094fd3cede483853aba4fcee7f04922040121368724719631aff6e202ea8f70ec805cbd9484171afbce394ae034cd0409d77f9aeabb49cccb82fad27156542f54c265b0717b0c0c762e0ea248c77d8e9f71463669605094;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f7d368f2310e21412ea776a5ef8bc8c510071e1b48b866223d78916d665fb21c53f9c65fe14643b7e7a1b0fa5b732e14412ea95fb76e88834c6d4d27f90543d349c2d1a17ccad1b0712dd67fe1972bc3b31ab0fcf9cec53ea8b5b17b247294686917deecccd31fa84981afed13f9f2cfbfb6274c01e5e569;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1692d44fd9e3946f136b0ca35aaad14c7cf69ca5211f7e364fc4cf574815329449f8b2b79a11c75648daa3ee26c0918e14b1282e56219608492bcfe083f9ca5110160cf3a771f8b3ec7cb2e7294bbc82891939d677d2762b5fdee12e94494436625f95e4df61afde60ce8e459fe78bc526ef89751482e0a3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191beb3e646420b87440cd0eca149d56aae71b9ce22e7794e633a8ded29986a024853aff83f39fea172047838fa16609d12365d82646088279e5f92e532f063b3b153645c19608a9ff9c4e2cdc1986e0e92c95e601aa9b58ec4ae99931a0eaebc0efdca9b66218eadf12072a456aea05e7d01d4f00514ecc5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62b945a44c5ae04c41149a913abcfcb23f69d781c608b065e3a8f968a6d6ea86810f390f87d0014374d4dc2acaab248ac1aee9cdc0623343f01b950e0a39a59fb1ef34f7555369f8cd0ec2f4e05a4f8d626feeaa402b8e63e22b662279ad4392929e161b1c2b6044321f15723f20f21ec553b1f04a62d2d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e395c150509e0fc8e4597699f55d2471db533070309a20ed056a6503226a25e5986ee3ccdb537aa2aac209b531441517151f78dfc0ce49d7fb836ba9731e43089fb2fef207920011d3bad43cc5d9ea67a1d9ee27a5a6353f1a6b2fe94ce683a3c9378411031a9acc132051105ab474a5f1fadac7f3de20d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd15a83830027a4421eb292b5ff82b0c04a73a837c37d15cbf3141cc15b5b894c2f4e68ab005f38e2bb853f1140ad05a33da2eba055ee4c5554d369ef02d5eae92fefb90fc23ffbb80498bcb6260a8de269d1dadf15e7ad66ec9b26a95be7fbe12f43e1dbb9d0ebcb7fc405cbae874ab7de5246fe8247b61;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb89209f1f060f0bdfb6db890a9781a72e2b8f8a5e2f3e8fcc0bb0b03ffc3dcd70a64caaf69f40442adba3bd1f6e717d9abdca0059e71b176a531a4f18d997f8ea0a2f878ea1d8878313bd673431196fc9c503a20f2fbcad22c81522d5003f634048c50bb1631a382bc25d04895045e221dba171913429a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha58f974a864ace3075a22205d6e6603974ed66f4a27ba33e2c93f05a4df0cd3a7d9f570a5bd2d21457e13b24356c9a245a770095f36cccd776e1d92d41f9a6ac9faf91dc9da5afe47f32fad7f1610a0eb30084ce351ecec5123e73e5820545ccb39d1a001b0d0ccfdb0daa5f50d0031c4a69e6b2fbcde788;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9136e77edf1d53a30a19ac0c850ecb5712a41d026b181f663aedeb9fe962ad9d501748d47ceec7dd19a993eda2e8aaa92ee7a24bbf1a66e1e97b310c2181a7d6b408abb1e8940dab4922749b2e827675ac0cc11b5186e4df3eeb3466978d36ab6dd4f7114bf3436b4554ed403f889c1c46a356667277b937;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15f523ceb27f285aff4f69e4a875da7c24cb772bf484c10758ccfdacc71c2a5fb86c539adc20a1c7d9b24ea80bdfeaf4608ca4cc2f024cfb0b357afdfafbfe37713f4f0188f0b8c4fb5acc26c39b05fd6e3708f5abd9ad70f494f7c9e3feaa9510f47578bddcd6a2a0f7e491a6ccf7c824b2b5b925abc78dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f23726b104ddae17c289ecebbb6575b85ce256e604df9057d6bef3cafcacdbb3556317f6ac799fee5c1f8b6848453791fa718782dc7510d109ee5fc23c53874d43ccbd9b3e38791d75d020153536aaf547c4fbc2e0a46dbeb84d3891be0343a4e2a13e7bccea23559c8436cd2531e53552295b27bee56ab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13a5f21857261c00ad77894cc7351d091cceed0bfe897f261a737705490c86e12b0d35d7e7e7a5bb01fbbed20e5d414313555aff41cbf215adf04b648a052f971b762cfb513b05580c8612704db8d0854df8a9690eb7091681428d800245a80a8da9e967b26c838dcbd949120e5ea6729790942dfbb597e8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h100ba5d116fc9693e95e678081b3aa9b2199013dbfdb400b673999186e5d4eac9b32ba93c00b63fcf6d69e5ccc4d199c9dbbcbf37ef45d4f9be3a564f21d2c97a58492a4b0f72732cda302aaf78edea80f9d6da9c12600f09906561254fb53dcd7169ca371d714a422f29066c767393e03c54644ed6aaff6d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1afbdbaf9df93f48c4948e838517c9fdcdafdb07dba4ec75d561a8549b5db30c2e475beccc04ea106bc240a7b4541f644b107097ab474cfc255a86c6647f963d9e272577c615c0c8d1e68c1ba14b0dadd9a421b8ce6afe06c01d0febea363a50bd59d2b83d156d0d7dda34e447d3c36ffad8c7578059a4202;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd16944280bb098632cb5eda2e57e90facc4e0bc7472cb591ea7d6a34e447bcdfc583fa461980b30c299ef9ab15e4c789ff5b62f36120f58bcaf9b64cf325fa0ddb7593e7419a3020c9d4ada27ea78c7a262535f8fa531cb066d99ff5152eaf327fd9fe89369cfd5e07c954b7f5bf24859535b90c5c76b64e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10487a19e216fdb127e23e745bfdb67d3a95de7be5cfbd41d260221452c5cecdc059d302e9ff790d5ade1e4f27987821478443ed35b4db5daba6b8f1beca04abfaacf22c56b89a88be3632c2ac1012cad40728fa33e90c2171b228264c611a2206daba99e12ce535d71f2e5d47506f41ed731de6e0a77de4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f87673e0e4329d877b6a11a98d7b17f0b71ecff18b68e4d63fab7046eb5a70ce800bca0725b4981609ff481f224a3fb086f0f902aeee6130395b20e5d5fae0fe709aefcf8db9c7174ca19cb86217c8d803157316a002229816b4218a8eb318f25146e10a49b2f57f34b7af755e2e15c7ab6d9d9625a0892;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12831d8cefae82cfbd1b2c23f0c61838e12e32a41e5ee0d8767b40d4302cf5d262bd1f2786043128ea121031dd0b7f805f4ff7be7376053156f58e9abf17c5971406df5dd2a3aa9bb3c0ca751287f3cde562753303b6db3fd48c41159b2620ff87bdf6d8a9b25eb7df3be7b8085cf0e7a1821e3f0a47de4ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h109ea4c3cc06751d74e4cab8a61f0d72014027e172522e6496237359dca159cd77580d8eff524ca61ebc52adc255d872c0f59f3993c8035044cde77437c4e88450bbb2ef67ee7fb63e190d97b78e7cdf26109044c68b585f769358f5c620cb41369b9cfb60b74e41577287e7ae6ad26233c66a2532eeda648;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a7d65d65e9fe50662413452602771cdefa54c43c51a03478914ae2ca67642c065d9eb2a95cc46d825082c31f238b4681208e157b18a7670a4fa2ee4f138106f24aea17004d87e0a438b347000e9e775f8c5570532f8c3e4edbf1bb9471ce031af92e8fece29a2bed89fd142852379920bec6a5e0951ae27;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd5acaac31c99f070d724c3aa60e64d3f757b403565793c1e86b4e5bfe1195773db161624bbabba55f85c434d4829eb5c2156791b84c09b653311ae1f0baaee288d85054216845f172d6910610f135e4f7dfce21bc6f430bba2e528962c284ac6810ed818d519bc6d33fa22d4f58e53b327394ea8bf7da5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h946a8d3fe242e471118c12992ace10b2ceed96a79d3f57563e1d5cdd2a0e2bf0a050d158089f6ab4946e8d7b1204d013d23856eab388ede43054f0cae4ece04092c8ff88321305c457ad317c0801a0fcf3a5d54cf4926ff3894a87491ca221cf7d1d8c59c33945910ef6b125c018fbd70b3e02da925f7182;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h141869e77d61868f20fdcfab67db02f7a0bf73f6b6f56119ada4653ed52a73c9fbd0ce2d8a54562a0b86125f2f21e5088255bb0657a2a7273cb7beeadb940c44d3bd7f77930688756c4b05442a720d98fe64639ab2f56043825d81b7ce7ac0b1f40d9664abf56c6d8cf5501e0aff54e25e61d9560220f9dba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6cc21d5df3a2a397bed3fc89d5fd5d7f17e77d9186abda3e51f060688b72794057340ab24e51ce556094a81f355ea395ffe9074fe7d78b5175d4212d40ec4e138cbb9e8a8b9b4d118ac4140d4d09b438698ed322a668deff613c826d76fa35f8cedce5ca677f783f07b3e3751b535f0cb97f4ae1341512c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h57ee9982e3023b717d2f543b0baca65ae91ba6d8b2ade2e5a0aea0be1b3e159610048dec159914b124d1873c6e204ea392121d2f847481661f07f3145393dd1aaff06c7e9ceccd84825b12fc283de33b9df3e9c10c901c5c1dae3a226c264d9d29cc0806ff51350ee785d169dffcac0db71538321d240b19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c183afdc922af3a2c4d31fde87e287c58a8e55a773de943f3eaf527f27df3c96999ecb671180c172898e41c16867babdacbbb9b10be3c34eaa4b280349bd75c0d0417218a3cddf8948d288e7bd9acf09cd248e9a09736729321aae8fd5109716a6e78424f65bd08a3632073b4fc4a409e9445898295518f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb3f9808223456dee79aba99d441dc0b17054a02fa787aa379b02e3859138ec288b8c67eaa7c6e416e3343251f3156a42d40f7180f0bf4ca668b30b36f99f3c8dc44d105d50f9d2ebadd6f0d4d02bcda7d85224f1e802b9fbc4719e82bd84ccc3239c144d65317224b37f55f32705af6134a91f68ea5849af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34b687fe6c52ad2288d54df54bc12b71fcef89372dbbc281e5e0e96b5ec6a9c34bec3e0e8a1f5107963c9604a1826c20956429dfb2859d6998255c52099cc1f1989e30ab3525905818ded8fc529f4bb634b9aa1d0f042a0d423a18e0311aaffc95fb468b5fe121f6991380670ed81795752f6f77ccdc98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4991c4407eb3d620fd5d111ce00243cf5b475e71a6f2095115f6d481f985270319bc63f0bf3915e68698a3ea6b604906d62e57aeb080f633f53ffd45dea874ed7f8ee63429016cc95095b00cea149a62b11d33c000f007316952535f4f10af4d26c1dac8d8a5ef9e15aca3284a1ad854cf107ece89ee1a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h132f00ba45ae97ee2916b2a80c648a6d349b4a3c40c47cf5e3107fd46b09ce0d4ead88ea7ad82a5f611067911a744eb6e683e92a658c7190e848ef87959327eab36474dc7d34317524b162bdef3ded71433c436ba2f44f9dbf296e7346b14f377cf56c997f203ba0e0036ab80ac6d397a7a628c5ed77ec873;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h435a1ba860516ea8b22fbdf29e4bdfd965b93c3e319c12a622a8a555fdcae086138bd2d871ffc235de083c7cfe54a005a9f782e091bb044dc1b9379016f3095d7788722fe71d05b44a09fe296d185901a62d1c786d4bf2753fc7d786b4a2037da5c1fea39f2a3d3af4c93729e6e0f788d231ecaab96cf648;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16729019784efc09d3aabd68631b3ab9ab9cfba4cb3fcc1684ba34cefac70806308cb85df6332b10b7b0499c81ad9ed2315af762dd34c0fa73c343262da72940641bee6b6c35905b511aa4ec05ef620e60ce42e068cf63ce7414c79d34403d02213730636edfd995bed96296087ecf0c52fcf3b8649985c03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82fee7ff59f97ae41d710a848320a7e8f40120ec799121133d58c032e050483f8d346f2f94af4acc2477f7a5952f6e0693a74e69ff3a5d99df901eb0e88dbf03ea1ffe4d615cc922c746c000a4a5f4e9348bfcd6288215339648499f1ca914afddaff214fb17c5f38e9ac5dd00747897519236d47e6aec98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6162ebafdb90ebb38373c14430e9d13409fdbcb1a4e0087f45ae1b6679806e23f8d0491f101d6e72cd982796243e8b87da482bd119b009246fd5cdcf2d91861fdf4b04fe4fbeb504a485cdacc435df53fb4819d2ee1bb09176af6fd59e8c543575cd6ed337214c6266ed1a3e7d89a94aee009ed831d32d57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hebc476814185644a69bedbbf5d0f18f23452ca8caad5e6c062ffb7c5d78ed5bc5f8df51b77a4852e066f8d358a6d9642a824b759046d3aaa7c0ca3d7b239e40d92fe40e5dd9e5bb75449e8c95f52a395d736c01cf8c7551b88700335021c6cf114656403a415a7c0b8d8b034b37242e20064ca73901cb4ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e026bb1758db148311bb00962533d85cad8c4e70be96222ba8a9e95cc2f5858ec11df59ad4ece57477dc45add4c6b0860d013a33d9735184424b8176765cf907568c41f55c0a25ba07479c0f498b6bd4204cff718bc0d9b71fe014a8b32eaba3e1b170bd2ee1ddebc119ac8a54c9ca20d647fe9a4a6a7b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h492fde04c3c56e39fbfe5f11e0610cfc549e70fc49eaa19579943508b5bbd99458b01ff7ae5218201da9fc0bd67aacbad4ff8f06719f231e019a6090e6801d848ae733148bb997ccf4270541964601c7808cf8952da5c3ef6c8fcfc76af5ef28e6f018e6b1567ccb8fe3719677c7384eaa86f5bf881123fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h177b01f0960df6e1ac283d3d2b5e3735c3f29557af710ba2de63dcab70a41580ef9a34be373386d62ef05419a0e934044be517f778a782e1d452892f3a8259bc7b275df58eb5167c57980ba82cd5ceff06a297fd8f4797ed6bbefc6ab252683433d92c0762ea645a87d53cb54b34646975c553c74e262053f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ac2723ee93fad4f132b71eec1aca7d4b459fd5e7e57d714f9934b184f1ef54f04dcbf4095c0d6c9c94a885d8c826cef62bd8f82b3d3654783acc8216852ce68a2f7635627ae79ec32c94c8606c2752f84bf561d3f5b1e46a3cab357b61c50076b758ebc793090fee14a9a15fa706a965e23b6eadfc5bca9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d138135bc82f77a337208ff4567d4acccea02422992ebb2a1e50b48edf8412d772bc31023c425282b5620ad34907044ce10edd6cb3c4e96a848b62bd33e12b23bd3b5e80e3a0c88b9d21231a48dfdfb1be16182e3bc9299627ec26fad029ca3e353652b09ca17bbbee7b22d0f3dcd31a49d00d2e4ea2eba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8044de9d33b9c302b21df00a8a351c309d128126b5533538617a6ae2437094dc821053dfd61c7331670336a176aa3a1bb53a8bc0d1893eeaa90f899c3d7c808c9293accf2bac3b7faef8154b0b567c898b0dd54d0b04b39faf50a1c8fdeb5f95704058bbe075eef99c6e17cbc2e2bf2c1f4e07b20ed9fa45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18d2fb8157a118fff83a1417c6c6066c9b3b726823c3a06bc20937ab7165bb2703555398c95eb2cdd7f39fb75f342860550069292fd08ed308f41db9709f5657dfff4537418c239045f81a7611826ee55f2e5c1a0d5cb9465eaf6472dfc58f9a512eb8f9f1602e5f51d72c9ba3190556efd8fbfae256e8a31;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8917fed713cf1cd9ccc718d054274f72b5a827a7487a06e9060d188d00b90a596a6e00e89bfedc8ff5759d042c09ac87deca7a947a5d927d49e6d6beb8735fc8def3a97d8bc0564ebc8c994c71df4c64a4fcca03370a1a47a5ee7d77fc495ce909c26100b6dd8ffdc7324090aaa5ca9b9907983b2dba37a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h870d82fe665c864023b57c23a0f164c442399352066b71ba52757bbb8b0e42a22a6d03ef40d9c1c10f32d868d93dab914557a4e123297ba0b0d848e5b0ef2b990620043c9cec13d1c06184c5ec0cb9e72a153c9fec2ac5349ff9471fa4fc53b348520410aee9ddd3a816a91c1c3b03f99823bc3d493abf1c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h126658312b550340ccc597b7a376121103f0b5a459c90cd20393be2612e606c758451fc06e843b63be05d61064d10ba931d2f6e315911c66f458d6b2b997fc5d63bb43bc1594f55834a4dbcd9cb9a33ea7b523b9bd0b7c53141e3ac87f1c92fa7c97075cf6be8b049688f9cdd182aa400a3ee9f4886e2408d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h530a98d178115f980c9970d64e5075ea0889b249d5d53fc26f0fe7721252b0f0366e36fc02005ac9925430e7f7bb540212199588a6a65d995bf4c047a77ba6577e1ffdb502ebcef589dfe7d50d80fca8bd299195d45115efc6f7844b499502cd69d5672260e71f60cdee25cbf389a8788855791ef73359df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h117889fb26f3cf34f6c13c6c4da7d1e2ab428c92214f665d0d34b1ff11cf21e9086534cf0c5303becc3a808dbb27115c4fc56112b9c4e6e6d423b86ebb0ecc694fa5ccfac1a11be206b556405a00a5b5206798e7c1a9dcdd3d9e95bb3e8830fcdee78cfe443137b66395f75e405339e6ebc047ce6064738e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d626eb3fd6225983c9e9daee77f24f33923b5f068330386025090be2f411f19ad5d1bfa6827dab49cd89f6777991f746636090eba82f06964cfde9b1902c8f5c9849ea835c0de181daef733e50eec88ee1803e178d39080e357b7376b5c406ffa882058d36c8856a313abbf4da4c5ecf5cb18d74fc9c30c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3fe72f9364f5be7da1abdc42b89bfd4f7429e91fa24cfcdbd0c386016fdcda68ecce8df1a7890b85bc3d52c6f67a542ed818655dce2ed4dd850417f93d8d77d3980111b87dd5516fbaf54b430c27604477eb4ac61842b1638ef6900cceee5d1e0006f6f91d1132c90a8bb9f7bc86c9bd6e04392d56663cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9b05ae903ede9cff3cf1a27befe16107176e91722399209106bd87abc9c1484b7ca15b96bc497b282046d15e3817bf9d12845c9646bed8b69d921f9b1cbe8476619c5df7b60a6e2d8ef158a4adc84acf9f291bfbbf9f63aa179e614f95003d9230b83720fb6f04c4c59a4ac39762bd987a4342d092c1a91;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec3894e850f76ceaaffb73ef81c9f13783d006da257779e7ea85b49c5820e9b68b2ad4b690075654931828ddb3bcb0baa4eeac241082b72076c3a157472d633853e7a866487f4037959722cf2fb2803b0c9ca6a25cde7e58bcee4856ed60981b56ace7e1eedec36c46331aa16f03757935b9cfa66a0c3626;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e63b10efcb906519bd1c6be838d274228efbeab80b00c252a8cc3b4a5090b196c1d2b4cb65cf8a30046cb426ea79ba08d894d4c0814d4f28fb11ec4ed707d64f04dd9bd2792774a76980015c8d30820a15199f9d2c1bf9b49710a831344d74164895e218b98305be6e7ecc58f08ae6bee07cfa65cf6985e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7f619b53230efde9afa303ebb5fae3551357e4f799034def6f74df3453c68fe03a5e3b504b19cf7c3d880f5505ceb62bca1f46958f5d09c87474e2f1078a3480d09481be6c982641f30f47c694e133a40edc00f0a50989908da075a0bb158fd72e34cb9b442ad53fc3cbc4f0ee9dd419d9a11470f10ac13a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0199a18a2d1e4be81f12ad917f75fb2a61d462a678b8d3ef3aed17989381de3a2313f7b50bc933c974a8835317e004376b8ef0ff59b28a5032fa2e05558e2166c213ad08b90ed0a7005d66cc86b707cf3bc62dbbb82ce7ab6e3e1532eb8b805719fa44c60be27abed69f640e7844bd0f74b7ec43f1b5a5c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc699a3eef8cfcbd98e53403543b7ad95d9e595e7f0bf5562a13c23628026f812a49efb75ca190586ac15ac8e4568764f56b2e15dea96291399608ee7c5fa1f52cf1021a8cfb80efe54ce444ac8a2686738d6663de40749ac40abab89a7d3816011314ab2cc7ef56bde93907ef53598bbc1503d4e59fef642;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha0591ea63b70d780e314c111c393ff43d0da7b84900f8a24416601249bb3802402f4ad649dd297d93c89fa5a2bbc9bbe21c1e01140883d749f663a791d160117addc87aa1b9fcf770432e41dbdabcd908f07bf6065461091268e0d9b4fe0e0d4558ef7dede3c18e5d846409acc2ed164444b93a079476b05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b45b19ebb25a5a9ed0e53ae75b7b2b05d772276875e2058a5d831be8275af6609933248d2f875318d644129a6eb1dc0d73ceac8fbbf2890a65845418bbad4f4e4bf8b24c337514d43aa5204ce5dd8a49bd1a4099b7be1a906d6d33204ff2cae6681e8674e024a8182cefa1af21c84e72fbb5c7351be423b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h819517f1601205aee3aff53e63bb6f7ee8aa20cf655716543a9c68587bc326722899c3f1243723c68f818d27f0aa3959874d1bce4ecd0a223dbefdb82bd053b49db4a62ad522c808417819bd44a7e21d3f23ed3fb46404d88b3c4be05e2fff3a3bce75927afc7d7725b6e3c20dd510bdb3459f1d1bad455c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d83719ffe6a5082dce9466a5e1a3ba060a756bae3394e7789170a2b644f7c89e2d08318e2214af39e337742ef729da4feb2e6e7798f806e8f4867b532361bb08607a8055d5f1a6bcc7eb2a8f6a2227d6a0bbbed96303756fd9bcd577c5f86733cfcc6863317d30211f2cfcda960723c223b1d804b36a3fdc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b7c61069fd93ff9df062ebddbdfa37084a25eb3f29eca3cc351b6d9521bb2aa51c46f2956982c1146c4f1c741f945a71a031a631591c1e58902ce8a7240983e4b07b32de6273897a17a82f6990aa47231a94ea79b37a01fd7049c9df7121aea37e014871c1aad881004fb3518c5e81146c51b22853847b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc128522920a5b8986be2db3b47c98abceba9324f334b36368c1e1800c9f36f02fa4f000fe454683550460d83a82e60be6ca5f35db97eae0efbc7ab35762cb20ecbb0747d1c65cb0f6d4328d04bfcb8f6dac62e7bdb1bcea018f001ddaf4a4322a804518505bb23ef0bd451ef3cf35f726e0883a2f7432992;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h62d86aaace6d0b56c90e9bf5fc756edbff3ff2ee0e059b88bcf76ca790507fd706f63fdde531f2732b244e572f31e0b4f32ddbea66d81ac0cfc8ff1c9960be981ffdc2a63cfb4e1f41dde1848522f3adc565a3d4077953c7d62e86ffebea712e7bd9607ad51ff27b4b11ae712c39cb90c503f9ad3a5c9d4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c495d3518926d8dffad4fd1c6c372d25235f5be30c4a90e892e7202869542143169a7bfe73db81167b2a23e7d8a2bbda9e5698e4a8b6c076d54155ff9a7e8174f3d0fcf8dea534d8c95252ad6beaf2169d6f23636c86f833a6a39d54b94f55b1cdef1e04126f83bf57d390c2ff08909388418d054157579;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13222276e5a1abd17d2411e3734b8c8e46045847ffe89c6a00b8b51ddb275e9a36c0684a4390ae7ac7efe2bc94e729693da3f6586b77591a428c20598a8af17f569ea7d445ffbbd0127407b5f6defe42edd14f413e6a40053f64c08096dc52c862cb2529f9e08482bdd8a36c76a7cfcfbc393ce742d57d409;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be5aea04a0c8b6b13dadd634befc302db097885e502b2830b5ff01c4ac01d55466e6a398ae747820bec7fac2013ea299f4e604030090b4e26c58d251220b48d5b6ebd3188543ea02a60d224c6b7a2ac1cdbe52bf761d8b31e841f463fd205c8611985f398a461b7671b53d8d7e469fab499458d7553019c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be0bf2119c5027dc72af04cdd923e29d2a3b284e27c00ba6de3b6bf1b0c48cca2b90a19644c2126031a85d4fffaf0949d127647cc6c9d4e8f16c2ec8f40e07e9c11a96e4ae5d1c5431deeb88c389c4aa039f1efb5a3a336cb03aab3f529c89854411fe3362a0aae27dd6560339327b363d580a0b5a7dae88;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f50ebf3bf2daf5be231be9dff062db2b8a968ed301ca7d04239d70e2ba0f9dac62c614e7f73e36a51f74d2cf63706238014095c611defcfaa9353b2c3cd8c7d8fe73b4dbe0999730236a76a351d2d63ac3278c523bba5348389413c6d10c7a00fe88a07ad0f89c619aa644aaf583c3e3b3ee16b18dbf61a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c5fb3cb831c9a1e69325959dc76ccd717a645b09636be0b6848a2b99709cc4ffd08bf95b2071ca1d0cd1375319904d9706e10a59a1adceaeec9970d51fa118cd305ea19d2bdad4f0f01a759ec3e27ccdb48d5bbea9626ae8f772cb9e67fec5309436128ea00fc39c017716888cb933f2cf9b1ab7fce3663;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h827b6fb2ef6e20c45ec3ba6ae953f3d30e1c3a028adb1dc4d015d764f4833163633583e380bac64262884d96f332b6afb3030ef33a247a5001fbd905182aaa22fe0c269247eae4c7e31d67fef894ef6530232b825741e74c15ceab2b71667d7026965fb593389477959193e28311feddc3e9a6a5caa0e9d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h470ebba8baf7f46f963e633a15d7ef7ec674d7e1e854d6a633062fd19e8f3da87b66f057e2da5b7f2cb850fc7c1259c36ff8f299fa4b8c55d219023b097379744eae1f044e6e4a58185f72e3003af9a02e2e20d9567c092b5c81cfff014e5d70556976dacc22fe961f737ec4d88a4d736a6d68fd1d81a16b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13194133ba83aac82fb7ee2557aeb0c38f8a5307cb632fcfb14019ed796399d99b34d8c8c78a7be41b49a628dfdd1f33edca600c852880bb561af3a39ffa85d7601a160de7ea328f48c09da86ca4f43aef958f3ba8c3fd2f8df5be9ba143fe1260628d8ef84d9c09f3610ab82bcf838fe9b483ff654b4043a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5f221bdfb1409b23b15d2a8f35ad85a428592e52600fb59b1b4ff59f0fcbb0bd12999e07b3425e073f737facaab33b1a90845b725fc47279120f7da5dd27ab1bd83c94a05d04d1ba1f02887c967409d9ef4b7103ba05bc32b96d5829a32560d9226c2ffcf243f547e80cf8197190c0dc91e9e640ccc575f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16acf9b55a1d41ecb0c56cf8be2fdb4c23832d30b417a80b6dc67c43afbffe3f6d7b32089fab8cc9d643b6f2c442c83683225c0bf3f407a984f0023dd8dfaa448b6ebd1fc67c8d8a1dedbf24c0831c7ac02f5c79c955c6445d5a9b61dc717306be5678b244c7c34e2742b8216d4e728c97c8e8d900856a995;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1390fc750295ad86e978276e850f81ca48bd508b1d025f72657a1b92035a045550f2aa1a0a066c52af5286ea8053b48302e4c6600528252816ad3af2f4f215ab1d5c223fb1f1f307287088767d66f601fd438f504c67ec1815b693d037613e6d573418bf45917c745cdc8e71ce103f08d118984435c20ef51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h75c98bba72e45e231c9edc82be17f5df52f54bce2c516eb8c356d83c53cbf1289530a03d706623bd4eee5725cd074808266e7ede73e56e3cfcd52e806bf48a247810c830e2dc32385ff883969e06322c41ae2a055c5ef67322c57cfd9626656f7811e48914f1cb3f1f6ed6844934e9d591bc9726c39122a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c82aa54bf3ea3536c8c62ce0c3e16487d5f118e8e4de718047a689c6acf97e9d9e7843951b19700c1340330ff8b890e2bd8eece9dfba2cc8f3a8dbc8639910732b98c37e18bea8d555ddb96d8ed5f250f70541834bad28728cddc43c82d180f0670abd7f861f502138959264424f96ea4df6456c04a7baf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5297235cb213a534b570dd7e7a49dca2a1bd7164bff9f66d25ee44e6bb6a4ec4539852ffd89ab14cbff0369fa6dc34c99161ba81f87b50f0314c62bd25ff999b9023661bb9d75052e04e8e82bba4b68566a83b0cb84a39d8c9ab42d62ff760e81a0b126ef711841d40825604589c25385bdbc1ce2d2d028;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdfa0cf740409b214141d0028b420262c2c7c3c80c3afa3eda0861f5893e986965afaa0fb8ce03293a3c91f024b3290a773ba5066cd90b81cdc4474fdadf012c0d8a92dbc009920c5f27a8d2bb382c41ff63e26810d832ebb331df7dd2a3e2faf281c19ea3b795778dd8051d14346391378b83034597628c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1871a44e089965822fcf0e33dea99ac8be3f7abc001857bbfb05868e0a289fe5c810225878a404803dd179c2d73736d5ec25527abcb22df0ce2351c5590f5e1aefd142da3ac0e2a462705ef47d371f18773067dddfcc33f04c04600de4a0c8e4d8dfb1d3df32ac5485af80c2dc230f66b738a1be9432168a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b8aa1ddbe61b341dc3acae4aabfcfac5c1af33dc18de35308efb17ca9cb1acaae7adc58970e5ad1d0803482ec09b7991c0ee13df4006e0db59b5c00725eb451a3d5f47c4c9624e5ff1498720d8ca516938fb5e8e0a8f1526074a8fc46e88eed55aaee72657b5bc36cd88a891798aee62eead06e42c160d71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a4357283336b96d565f4b6af4346c9decfc658e12c7066312ba82b285054bd44f544b40d9d9e72d2ea4e0fbd7c66b7bf1cb8f1cbeef2c410d6968fda064e99efc79be566949402b26d10a3cbd5ed8b608b8aa1a8dcf0ab7850bff9e5aa89cb1a0d59d7a426eb3dab91745a3377de3cba0a4194e782a3d64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1293eb3a9d2240facce001decc5ed12cddf77ecc49138a536a0dd1d7315b126172626ccea81df19b69e2ecaaa66872628cfdd2ac03705d9ccbfa90d393f3a7e83486eadc01e123496b830e2aff01d81414df4ec1d459ca0ee3bb22d5e01e5b18f4652dbb872075835cd0c25f00290a868308d03ac582c1e1e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168d17c18eaa3de9e56fdafd1722a1a3772168b60c77812dce3ddb575fddab22844e0e133e2f1eeda1ca6e117de2b21e33c66ea5103b21eb6ffc891039a569e696182a8e38d506057c71dcadc0a6af3ed5109e561d8fa271347a5998919b61f3a3c4dbaef56809da0b1516155a72b52afe1d1fa963f681e5c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha487a7120e1435b4646ba5cb9906ce93a8a3206c26a6e349a45111ea55d2680c920bbaeebfa8d15abad6ccda4382eadc172c7d1dde2566b02daba7929b34187eb1613817bc11559a0fc7284923e614a36ae249dd7e5145d8e9616b66b0b89b58da58a013bf501d1db46bbcdfeadf3ec30ee8550dea848f33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154cc3aa683d8fdd0068e67da84a571c40841da38fe57c42564943a42d60478f49ac0e434faaec10902a7fb93640bec0506d34e8021b0b930facfa7d96528427df1152acf04a8c72a8a35d5ebb0cd9d9faae033b9d787b289ea03cf341b07085b6bbcc81286a8690b4b6b6c8d5f9a8f9fbfeccf97e3cb3612;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h170b0ca296f301ebcc1ca764532558787b7d53ea8464c2856c2b48c538a4128c1d39d42f31ac1345b5090a54db6f95b7de375d0b4b9561062e71b58c1646720829dd79efcc91ada8178db6b0f25bb3b50b1b2ddf63b01bde82f4f29168715f51b0c53ef366518c5689a1434c31393ae65f8cb6381efb93b3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h178eb53cdf1014cb4d75dcf8d5701ed9c96c2f608890f3bc987c8e20632138b51c4a6b1ba205986b30f6f65000b05d733e7b5cfd42da3984e6dfc588ba0edc64ff9c83bbdec95a98d450f524a73ae57751dd0bf7ba4336ec7c098c44186f57b2c589f4d168642be6f83f128ddb94497191b1c4d49efd89248;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a33d06c2587d60850b02a1901917f0c03873202bb36501f55000133010099c27c979fc4b733fc4a13dd841f674de1db8f3462908f8bca14dc7514d6496c5aa23d891d69f52599d379c0d70f26e3db3743cc6a8b9211132bb8bea797b171875025bbcc5e71551605ad359ca7fa7f8d41abe9459eb9f62ec70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1060b68c08180b85e43b2e941d986310317a32b63da8957e6570027a63ea7010f029b38e8b3621545da0f9f7c2a1c05e4cc9609ea523095413a6cfa3daa6806238f96a745e094559c9367e9c37a26b39e801d726c05d6634a74b51ec6b27a991add5db136be1474ccda2d1e75fa71906bde5a9aecff14287b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h452b73aba6cf57f282ede78ca9f829971885823418ec376e289a89f035782ca65ac34d6a4fbaa4061e99d2520784de7fa85b7b35802cc6da7f9845aae987b21328e2c8997fd91ec17554ea5dbfac4d4f3c29681dde082289cec0e0bc0a29dc74fc00c06c9d46b106d2bf686b38b8ddfca17647170a621faa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c7a916871b7ce7002d820b0bf1f0e0bc58d53d2dc075db9478199e0beac9f913f82a2980c432278b5a8db12a6b0e9a12af65b389e7116f8cb5a7a5f054cdaf798c8a2199485fa2e28b00fcc73e4c0c481d66d31bd7c7a62d387f586e89455d56bec30a568cb7416b042a6d996e702bfb1db384d76a14327;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc79e01f929e0730f1d19c44b044f57df57324afe5509fccdf194b100dea7ebbda9bbbdbdfa6ca6c4d4549a4dadef05bd41e9acce89b0f0fd981a15de709bd0840f1186c921c553020574ef01368151c85e371041ef0e12ce38e69f7ad3d1d6684802b76995641d7d0d36589e218d5460c4a28657a1621c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ebe3cbb27a61b9d0be61921bcae47e3fbf478ee8a6fe0a21c01a8e0767a5536cf8059d8eb2bc8535a07cf579812833f4cbb72593e7ecce705739e5dad0e86ed38950aba247c2bddd115aea00e38abc82449b410697bdef3dfcbf1fceada101ef92f7aff18b88ef6e707b9759796796fa5ce33ced47925d78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17029c7e0430eddef8f38f6a5290f9f9af9927707c09fe0906f74fe86e97f45f72f4e9ae63fb09aa50ba1ab1ba6e2778bbeeb4881e428bf75dee0899545a61e7373674566d4cba3f8be9221385d0d0308e81519506cb2e8b6943cae4afbc10f93c8fbe0f3b62570c48ad740a9d2008202782c023978aa02dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7679537fe7a95bed1c4acc4d6782eeb65255e3e2b6317a1940b81b2c8c091786aaded6ef09fd53d279c772b4128ab1b3a0df89d123037bd899b592cbb92fc6c9238c2fcc7a598105437722858acf14775a65528df92fb9cf7f3bc54c7ac8b9f912508f940cb045051f66a3394477cc32b49663827767b998;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he7e6e416dbb3e6c96b795b8f87d0e78cdc55b89cbd59cf95f11fd932d21a10b948970eb67f16f6cb9c46646f9fdaf59e2deaba444f410b5c3520fcac9955cca6a72b6769c04b6bf3d2e047bc5bbaa65e5572128d8cebdef6601b8144173fb425bebec201503d7349e9cf87a11fa27b43cb8c5a701b56cac4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h198515c524fe88dac31ec9a1ed808224d9db02b841476a9246136fc0f27f1df999541f08ad568bba83b5b6b59d86dd2d349a6c47968c975d21158d32ca8177d93ca053d2cc5e1f60d5f9ecd791af8a159e05ff80dc0a4efd43b533322932eaceb61c8446a5eaa313679c073dc61fae7fe011a524f2ada6002;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39974447f217c1bb77d1a4c0799a1f03ee725df2ae157186feb67314062585f3a4408f6c4de97c6056be677030e79b2fb6de9d16386fe0cd1d2012b0d51a25f68bb9172eec736534cc94d6e4107b9aea3be42b813d237a38cb8d70f389ed631408e3613016dacc69853be7c96e4a45eaf893d8af63d0ad67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f453f9ef67ead3b32b75c316480011f38885115a24c9a8e163512a0a01c2f90efb43798d4855c7f056b172d4e94bdba3b018d9e39f3008fd955742eba78ebd5ba2ba013bb7316cbc5aa45261b6413fdbbc1c6c7f6de109b9f8d12f3e3e909b3374d08f4c37033f796ad96b0085026d5543e893dae593635;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7225cdfa60d074d0800f2d536fcbaedb7b1b9a76d4f356a7acdee71b38447d887f0da5ed146ccb45f3811ae7f30ff436a0dd8f780bbdc767a7022bc12022962816a4410ab33aed865d4834a962ee06a8fd7cfdd62cfd8286dcb6d79014180c01148fd94ce8d951fba289c6826dfe8aebf2a459fe45224894;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1871af02b9ec9979eb989c455c1cd74dc4b8a85c428f713f411f47d2d96d70801805e5a2aa67a5ec725107f56f102f726f25bdd660a7ed84b2ad09c08adb4f28642d534cec053b0d679fcc9dd20da6ab1d4025e7171810993598fc623e87d8bf0cf1fc646b7971fc8cb5bf6341d20267a6d6bf3df9de84e09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1529df6aca1419bc38e419ca4919bcc6f406a647e20c9cb0922587ca76fcc9b2b7b0b165f1ceb1fdfd92329e9001df55a02dfb160b644565724b9f857f1ace4bd6f927216042b76dd820b7c9067adbee9e37e5e552e1983f156fd3a0f330c3f425e12372b80d581e02e6672cd6434b2ab7464ba93e36064fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6eedb32b476990b9efad6bbf872eaa3ff0dfc0b2e9e5c31d9c1978ac41d8870f532d0175740d054c066e7fa3afde1c7ce46783c2d89e06a9974ef3d91150e9da6a44b44d56adc306dae1cfbac96f635a2ab570857d3519e69acf296f3679a2596c4919034e02ad6a4c1212738fb21889e6c7f735f92cdc61;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdcd733f13bd9fd535df0ac38a74ce67159b3745afc18507640503be8413f58e521080690d93a52e112df4dce91254867c707e048ea9687fd2ec199bd849de1f321e5ad8ffa2c379739ebe6379023e04d6010e716115d69326dc7bf59b33661bf636cb76f05f5a628a2b54ef066dbc5c15ecece96ba958509;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he60f1735383ac8ae7b3921f6fd657469cd728de4d6bad917a11d27b94943148dc216021ed778740d605e851b56cc36164d5813e78731c83c843ffa6269dfcdc6687c880f05cf08e4eac782b54c110167a3bdb648b26dc53217c4dde131cda3d609b1226dac4bfa546489e776b34449648c274cf2df3237ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb80c4ba0d07d909874cba5ffc7763f3db9a2c766f4dd31e43d70d3701cdc547d396b9aec6579090b4f0679d9393140fad85f939e439e109174a110ab13ab6f1e844310e5ee0e35280354209f81cfab032fd69be1dbabb2c330a36bcd588b01f44ab0f629661ce18a08ca9f4ee141ba1714a8e4a6e5eb083f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70965046b5ee11f386ed86e03236b5c8ea2f336e6a3b6e5ab65f8305177822a129ceffc20f49c847a1d4bc17919b97c39a43542922c6c4357e01b3cd6ddfdb2af0e126783b8731642800873fe4bf94fcc01079d745ebd7bc12fb86024e0d4e342a28d1bf71f39b9dc3f23887acaa32c7e1949f540dbf2323;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb671727bc2d54565af7ced4a89022551f625ad88ea9dec530dce99c98cc5436776d49678bf8aeacc7baaff7b59d38d22a89b379f4175a9df52b07a3ffd4eaa9f0a36952165a22e9fa023b91adde60bdb204a88d697437df7f1a888ff3501bc5ea8de41ee6badb826fe30a5359eb337d4316d644acfc51afc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172fca32db623ecb9e3530b57883e63c0176f2b22d140a775d4295d7803787bb84f28bea8d43e3163a72a589e6376e57950d8eb635a43e1a56d4e9bcb3f5a25389f55145217d949a872188d8b6ce9869cedc0fb517517b7c7cb8934485a3d1c3a9a41c0cfd8fccef70f4b4bbfe86e4146681b5838b96ed324;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12da4ec8d10737b66a45b3e2326ea0fcb8a89d4b3d7a9722a7541f6d495693bb40573dc0296f8b1e6d0ccec85d8171658b4bd279567b8e0da3262ed6e09bf7ce73ffc081f830321ccbba00da59ea8d302c7867344d7cdb8405c59122cbcd78945505ac7178c2ba0d596ee1462791d2370f4c85fced7b1a505;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h51bf690e8d9fa2d2d9d9ca7f96d66c13610513ad2ca18e279d424e5b4bcd1df880bfd6dc9b0f240989a714ecde44f3ddb8738747d4be17976e9cab4560f5f12b68714cb69d07bb90ecba00923a2c4203cb25df4fe268ba0be6dae5f3fcfed16b96af61cb7841fca842ab2085b4d1550a20b021eef0c0569f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bccaeac9b12609493f17422edebc86f2451e49aa633c77d80944f79ad4e3da2062f7aad404a028576a53f87decefb62d02ab6d15b70ddc8f1afb8c0b5e07dbb0ecb00a507470c79a5fe5e3536d33fc91dd62024b684486213df5702310863b940f681ea591a768a7192865d9bbb904233727a9e472ae8e69;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2478482e66bc7ba1ceba98233058fdcbec1c12e90340cae5955c1d7ef4f9e6ccf68ff72370a37ea613cfbd01778168df95700317916c9480cfe4ac4aa21afafbe5e121b0e83f88c2eec64925184b9eb361c7bdbdc1355b394fcae034403e84bbd6ba66d433822c12d763473ab0f533c227b09c7c5bfb15dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4596b95bcfed15336bb69a8ce1746c6196ee8023c6aebdcfaace886aa49d0e17b4e93ac379722bfd44321d26f5fbbe55782ec61663042337bc591fa7fa6dcc011ebef84e456d2aaa4d09db3ae6113db35966dbc61ac2373362938613702898d8843cfbd776aae9b8c283448ea2656cac407959537bcfad6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19896ef5611ed1077c6b43a693495a2561dbb6766fe17909ebd1fc2c3d96aef3c5eb87abc0ca9922db8383318f1fff9fca766d38dd47b98ae7f51e6d6cc18077c5d21f5c0b41138e1ccb0f977602a8144e5cf412a86148780afdbba2454ff4f1640776d81810d3dff5f2d5776d9bcda25290f3c01111443bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1002b3d098d94e021de40eacc8c144a5cb1777e53392fe6d4d0c0c9e0fa673ab3c14ff1ff78d706e55a11ba0da0cf6767f5b198265da351e44b46ccce9e9f76c3b896586dc098f259e9c6d0a8edb44d8d88e4100e4b945049a3a830651418ba01c4a853a957fef0e5f34f0286411712986e9e01f3d74e2324;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h110d4e8a8aa485245cff62457ea36a5828fe91fcde907e0bec9155f780579903a45e4401b7b3ffac3e55f0b34e63953599306f8a78d5962797429cdadd888c4b528843c258330b6b2f2820fd9261c6c75d024bf136a36ebebd6f5c95edc98129f439500df4dd71c2ab8f040accba6af948e822116271a7372;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb9d645659fc5b36d055228586602f9f9fd0380facd3a5a7874136f8ecb37545c9576c7541e73c5a6e138dacd26b337e0054c319a3322cfa3b555702a865717e76b6a2d65ef0841ba0486a768de4b5af246077bc10aedb8510faf5d81285380b23cb62249ac796b3f962db48f492da78ac17976c59d5855d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187dddf0cb5e26d04a58a424a38b33285a7640abee3ce1c01b94278c422d4074fb927101556516a1adb9c4b8514092d52dc5bca07e911aefa9431127d581f70aa3269826096f7d1bdd2f5af34c9542fde7a4f526cc939007c48912d6c3270b4af9889271cf3d6d1944524329ecb2372409d09466b548d41ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b41d4f0ff95008a78fc7e1db51aaa18ec3e02d23eec0615bb3386af832893002eaec4bbaccbaeb2772fc4f3b0c70b9edc982bdcf2d7dcb47399825ce34fe9661004203966e001f63cd0fb4d9132cc7654a81a2e8e260d53f6500f28b610c91026eb8e20d578bf27842a2770774102ab85b3796afa6aea21e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c8fba2583e9cf57696b2f1bfcbc54d060fb01e1c26e9b2cd8e2310de7dee7914fdced91d2dd6ddf4fc50cebb4faaf72730869378fdf70ca0dc9fb16e97b135b59c27f5e1e4ae8f0d15fd31af22251a64b87b1a1b8a5e780fd0b65b7450cf733a2f407317ad2942dba4100ad3158f084075f9ada531684e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h82933eaca67a5bc3b7658ba06005ea1974e6b3c48cf666ff92a279f791d9d281fcc84dc077c07cc5789b4519932d80a771963f0cdf0d7f5b049c259fe70b50d12bd9d73b1fab74551e6b4d54b59764987daeeb788fb4bde6dfb8285bc9367fbf57891370eb8bd3780dc80e1899438dfd3aacd53a31cf7808;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e8d1a53cf06f2f495076cc1fc5bf0eff250f35dd7c525cc01283026e8f26ab11a4bd994087f5b1eab568a0505d614367b1cbe738ce1876d6d05809e9df39666983353b3bf736e1654c0d7cd83ca16a9f61d39ed9c6e9ed4e8ec58dcb281a8590c71b5f9e38e4a355d5d08bd4abfd32421c2cf51291092b06;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1edb7677e7498699828bfabea5a6e679ed25dc2d560233e80a532242068f77bb2703bf79121f3bcf477d90f55b8aeea9554a4a5fd3aaf71690307a8e07ece85a51d5ee3ca360bed92baf344b34a2c34c7ce1bcd2d41d880289e17f3e1e5e467d66f4f8873fc088c66eb1c62627c1375c8f74b0b3ebfb8a28c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb154239a9879a9176e194be5449948187c069e69ab806dfea85b2422cb69b5c1906f1fc5a0c7cf0baf57a264f9cf33b28757e9217caf7438ab01a89d1dd6642fc69dfa890623bb656971fde8559b1b7fc21c7054b58e5edce3ae7dd36ceff7e2862c5ea4a2d3d925516e183c073f6066531f81cd8817227;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f8cccc65c9c4fbdbc287a6dc7f1f868a8b73c99e680b70a863198edc0d1d98903e7ec58e5c705a833d210f2d1351ffe05bdafd1286ec43cff1b3635e169a11e13fc0fd1549a29c831034790f19ec237a9caaa504e4034a6a6cd1b4239705f832c83d14005d17cca24759e3dd742ed1985e6386c4ec7e093;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h364bcdbc62766c90d48ff8bf32e74eed19c935cb7efc6514ff3a8440198bd8383454363307b90f2b389fe12c1ecf8103f05b38fcf6dea8b6f6d0fecb40405488246b4a6f1e248d337c62fb7e7538bdb979fc8b02fa50d4a147cdfb112b27533af6aad005fc5cf8086177b2d8d622f3ba140866aed5a6d786;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d8d0ae84f2841519c50d4232f4fe30e6ddaa7e7860155a05fc4e50816da5f47282f69d4b4e0e2bd61eb5387b3dfcea529f3028561411bc960bbb3911abe3b01d1e11575e46477f9560cafaa93c46ba636904d74a669d114a79d8c5c39615f48731d404d3b99b7960cd3279613dfe939b20480528cdc3890;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dddf64a469c2de3d409161c6bfe0449b537b08ccef6c276089fb6051b72e69563cd05ece5f24622c8f3bdfe96feec10ddfa67e6af9504bc3be0868cd029c7c4e4cb84fd6384bfb7ab4a8d96aba05343630e8119fcebc613b4521862845141d9e1b5dc43e87125c27c49d6813381b88395a3401caadf7a6d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf50a090e0c9f643f3292e2d064e197535f9a95730b2f178c2af764b4aafb012b329cf5be1121fb98e0904e1ff56e4cf921b734c4323cb514e87be9ea11ce21106f7dcb8efb9cda35d11efa4b8b7fe71cdf6cdfcdc69fa8746629a4b6e36d5195ffe1158b7d4f5e2d14b8d7a3222dbef54eeac9d1519b9d5b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd611802ef77892890f6790ee98ed47788aa5d1aba8a623df92a0a7039c070c148133006ecaca175034e0864e37d04e3e53ef5c4821d61e3fac401b9ab21231d556954014d8f79bda20b9362a3f23453a0d7d03cf933979b3d41366b0a746dff46e670e24849fa4524665f21a633361a1c1d3161675e341cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1253a3b0ff5097063807eab5735e31881bd11624c1454392930d2f41cb5e5b066bdf7114f1a795a344a275bfcf60dfb2604dc4f4d263b4253e676b542e193f56fee8037b022a104250504396775ef08e808781b25262c6c012418b28e19e44d2e02b5ad6872a2160cae30b7b8334df3e816b0ca334b5fca9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2698d52729954db620cfaf983178d0abbc2447af2f6fd372806a538c0b31a72cffa4751af4282dae1dcc24a8e23a799b65a4fde94b20e2c564cb6f1fb9f143e5194991d353df81be24103f54b73ed3d439a9d287411186c3b480787250baa2880a0dedb9bb06de0100ddda40f85d9842d7acaf5805bcc465;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc726fa84abfc8272ae4f0f21eed0ecf59567801eb4536ec4ed091fa7a93005932e5540f616c6a7c8780e32cb47406d319798b851e55f2d0e553e100df341ff48e9ed42a866462e4fcb3d9179dc3edb41a9516b099f01d79c562d90ca3b3110398a95d6661ff0626102465d3c3c0be21bb738d85738838d2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h173e33b930454ad6c0574135e1fb5977c5ea33b1696b5acadf6ed06a30731ac60cc2b1720845fbd017ffd5651802c2a3bc909dc281196eb76e2aafea4a78971f3ff3818d14665fac70af4ac34100ae91ea57a7aed14ada1c8a867e24ea1a212c3476486a3324c4e7b4953a44078f74877a70f72c49b0774;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f79ac534ed6cef9acd3e84f9924a4618f35ad766a01e4281c7accc8fa497cfa333ba3dc532ce8e22cd9171ea62a652c6434ca70e52b05e32c42307e09b3d462ac13fe2560cad9f9794bbe959dee156a15ba7a48c115ea44ab51dbd102f936591326230cfe6ed06930fee66ab53949704005a0228426dcf6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b4b1ab285eb9ec814cfa9adb5ff398687d09ad81dd212c1be2323975765c587e870c5d73d1b0b358e10f17f82a210afc31c00f13804a837595584ff600ca787fa7caa6c825b7c9e2db794c60e1ca584b997ae58799f73c5957100c12494dce69ea4d797c98519adb293d8becf2bc025874c04605b7e3ebd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h151c6a4e1673d62a7d6c219a4e96c582014cd4dcb5b1a4346d8cd0b483189c289e73129635fa6568dc9d69ef948352144c342c9f54073a7f0b6fc1ef18842a906860a8d09745d0fd43c720df6cc6e191a94e83389b98e80d25803d1941d0168cd4753e6e356940975f22e908d8f244d1810147bdffa68d39d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1b88968881fbf8c0884b8ce94ee32cf7e623746cb5cf7c6c2eb17d8b57ef9038df5dd3d71545f008d863412445f437de6032a1c70af78e9b6028137e3372aa1fb5b6dfd6e631475fed7ffe6fac24727e3f463f18a2b8de1cb37f49934962a3021e38a7c3c05ccbeb605d2db94cbcd64cf274c44d5cc0072;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e27eea26a1be50f9841c9f75dc0494c7add6f66f550d4e218c1c43b9875f88319c2049cb5719040c5a43b564d468cb23238df0659b0072f3603b830a570319ab94615abe52c268c9c0aebd407501b7928ab23d7fa02c78c104f5017bda126d626b9010d22bee23afc8e6532615afb4a95288ed838c857b1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc9f63d4d3cc8a4005df39f2c765b4f40c46deb2f42430990e2278ba0fa46a1eb0d7b700984d77d18da30117c7ce0e81ee830fd90d678c85b8b9b62468eb1e92eca29c1933b3ac7285a426f46b4acb977fabe2ffe95e3dd09612e2fea0fcd49085281b8db8ee8b302078bf3bd2d696aa06f4edb69d3009f86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5d02dd92610d2c009de4f3836eb2f0a2347001e2594908244282190fc80e47ecd317533ad8efa3f51ffada35391516dc1bef92d3e95444dd1b99228b561de107fa0d459d5d76828ff5d0c1ef2c6ea331cce62be1d6940c15b4116cde68d862b291d4c717ec3f9b50013f63c906424ddd28fed7f5fd70687;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb97936c5e7814ef9d16b8353d1ad166bd251d975344a168ee05690dd3e6607ab39648a443c5f95f491a3df56a0eedbe6793c1d2a8de22e1533539d5957d1ca8d23265e51aa96c7bdbd0ced44ebceb6493aad893f21f49af49e89e9168152fb59702058243ad5cddad651f1e596dab88d88552cfb6eac66d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h126dd24f2cb33a6b57f4dc94853aca40487fc454d73f073bc7af4c6495d5fb9a91872b4a47515844427897f03bafe972e86ba6f6b2f38983aa5c6474c4b517b911d749b24cac1d70687ac4f2211d9a60ea4fe6ffd6bab71d7c8375cd0eeaaffa658971cf5ce5716f4e94e01f0fbbaa446f4702b7102a31c8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6ef94215846610988f21cf72467948a61f35a4d90c2e80a39015b9336329f766c4876d7d8999cc27533c794d614aac556c9e5ea1820dc0985443719ffa5d3a855edebc44b320d68436d40f2d18e9b80cfe01f5aa9c9ca9d15164f57584b5eea88dd0f7a58e2b60284d5c48ba5c13d64f4ca756471c8d274c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a37a4f993ce95735dbffae213f39dafee1fef737e65357b11c3bdb6dff7ebec2f83d45acdcd28902c106a43785d6a5c1f6108f480450ffeff43016beb7d4c09a6cad270a47213574ac6210bcc83b8a68a4422ceba01c3b931d6e5a8d6c54370c31288c90a6f69ed7bc3dc631c00e5a363217d2e7f5340f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c7d940adb41f14dcb412377b492efdedb9a668c9193d6ab99aaf7aaebc61120755e2b9918371232fb83ce1a7838a01439d2a05e151256891b885674ba336aa199d067d77787b4770b63f7894f11ef17deb8dca597603e5ceac4aa190ca71547d4bac2d5b369143348d415091d06679c1943c4a3353832b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182d15ba6de2a24315538af63ca04b4b45109a844358eb91b07a376607e92b56d3bd27b10a33fa4a2a2cb4ede817534297bf2bb1801dd4eea70c6b902642c7515a7705c6aea790ed8c056fd6048fef6f51d65023c71e68a5a14c9d25bd775941fef47cd3d3254c33995986993dba51db09fca9773e33d96ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc351e5c212bd5490fc57d6d5358b12821fc837343e302f84b88febc07bae0c1c191d5a0f30d2a31b24cf18ad7955205eec5b0af9c3f4440bf12242610e5f3c222a4b04c60361d1f558aa2b7afa076b02d0f7d300df4dfb96df68ebdd416532ceaad6db77857037a803f49917ba49eb100ce9432f866590e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10645825acde3a0e428f164811dc45c13b82d380c3aac9506311fbd12037d49939b29ce164c5c6cac41ad8539808a12d4296cda73236ecfcd0de7de9c87fa3aeac090ea6ef9922aac1699de67270f510d6fa2ea1be91c8e679ea1d4a074a000b23560395664cbda5422ba09c7b946ba8ee0d8a178eab3ab43;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcdb2fb37835127d731dce7a4d1dfb3b3f6e4114b87fe0281799d6227eba990b425c06a4bf530d320189e152c494f00bcd82ce55a836ea82158632396c3749be24d7d18f68524e6d20eaa1e6fdbfd2988e5319505929d347c8b210812229838ea6cafdf5c9e2943e4893666e4b5bd35bacf952fec4c622093;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1106c2c1158cab16379720e0ea09906b435473dd206b8510cece2dcdc4c657b761a693fdf47bda849dbc21af787a1576b19be898a54f9f4750c93398d01d2dfff8c1169acb7071fd1a18f8369d40601a07bd82790808a5baf217d8a22a7ea3726b48803a099008f6894800458ac00260657366923552e63aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3374a3d1cea380191efb2c7a3b42b0964780c5ee7e44a1bb8993e2a50ae53079db6333824a6519d7ae33cbafb0a6d8ebf7f3b389d0656d740d6317a6faef7d2d08a764635f8690234ed21379c04eb83a0966e6dcbd658eb27d44ac4b3e9901f1ca4880480ba14af8491bc28d6241ff0d2747f84b3f07e89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2b55a91e5a0c540267f1cd55f34603dab47b3be6030731c525f58748e9aadeec0740ab4560e6393872b7b3015f1fdc3c64937f661d03153d6690aad91df9b871977388619d1682bee815ee87867677764a2f41ca0fe9656e443d64ea6a0e192e3a9f3fa9d8b2a3b558e364b5cb092c5801564a0078b144b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165b193c5aecca6f342dc75db80e94508d60c66ef4868caf42908aff26086a69af4cfa0f6410451e96877ab88f13b41ef12729ed0e6bb365cbfd02c7f6fa7f84d181e95f8448ba11cb1f07ebd629dedde2d69a33dd5944bf4546f1c5ac7d84676ccd0b291a209b888ed6d194876fd4013f8988003c7476099;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19621a87da78f1ea50b89c9b2fa9cae7eddb071c91fcfea885261dd4bbd6c62252d767802dc3c124671cf3f99b3c754dd27fa5fa1e77b90ae692156fb6da45a3619060d6f4dc748d595d3f1ebbe67fa7eec786216ac3605220019e72b3eb37d2bdd94ea0df738055306c0985f0493edc81eddfcd780582793;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1879fedd64239f0eefeaf8e9ca060f2c6934780f6e8ac1b9d8f2865192995713ae18ebdcdc96a5458327181018504f4e4d89fd5caca62dfc810e55b660bf4dfd62037fa7d3dda7ea418acd73bde8c3ff35cfd5ba2fe6c281c55797d03a3c8e57a0dd619ec0e6f43fe8c7821146d19c76cb348030a0fbb3c7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f36a9fb84c9fa541aca5948a5e3c7ef45ef9b92a2b120347a6440712f40eedda5deae446e77bcc78643c95a1e4b8af84de637e057134220302b6c3130600dbcabf0982a1a58a89ad639d7285c98236d1e2ec467d8879ab35efb376d96e75931323fdec0f9ae321d2a603f3025e70bdd37fbdfc7176f36124;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f3a7ee33c74283631f7e2d514146bb68348c0a25e7e32a2555008b571f854ebae974e1a90376fcc5c7f786dfa6d3226641499e8d81035d31dc8c19dec74b20566bd1c77f9500cecb956781ca1c402092afbaaa0c44a396bbf069c5a253a21034a26970fe2ed612f7c0034f07228436032fb7dea37bc56c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb4400c05d41b2c4518f90ed2ec798c569a788fb67fd92f9feff597c47ea4fbaea7893b2663435a9b3b15f80198cbce7e47ca069b5aa1a614c08b2ea59f96b7896843865316ab9cc1d581e671c01d01479131df6daefec9581ec4fdd1645bf2ee0e6cf039e7ec0959ff510a184b4d16013a233f58d7c87c74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11eea8930a81a0c5e0e1a575316c368dec1aed206bdbc1d17d15aa64917d6c3039fab419b52b9609754f5f4e505b61c2d4485e5b51d2e7eb72aaff58ceff7f1b102981d78ebfeba066ddf7756ef2f7f4141006409a1f77f7198feca72642bb29f60b30b6e766ca3fa4406f3bbefd07dacf0a6bec191d6715d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7568dbe44a034b03a5a0cf87589a07c627914090c15cd950533dbfa993ae455eb715c4e22e3d5a5243ae579ac7ab1396f8eea7cb35b73b855087ba8af07f019b2421b1f9a91a321e885a6ce83c1ea800ed4e12eb1feed15ebd98ff9a636020c28e4b34051d211bba6e6bcd00c8c2f261c4d032f6bb6f6b1a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10763390c6fde8f51acb8ada4374eacc53f804554c78c554cf9de65532ec3f8ce9a68843d19fbde4e0f9dbbccc60b7959c8187b549ecf5e64517a286f9d150a9f590fd34ee0543e80e206792f0bcf1187d333729785740a9771968a0a3af0a05da79debf09a4296d8e52ff16c8634b6d7d3249b70f5794d6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c30252c901eadf29aab54e43238d59a0a5bd8365b8914d6a125d395eb6e6e4404911715d867b94c5deffc2c5484462c80c1fcb35180cffeae1090630976baa33fb7823c6c1e9bd32892644a041102c01e40b04609f155f387b939bf931cbd7d0c2fe4a85dbff587c07ba39984b856c21c902c23d6e1eb788;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa38524e18eefe66e7772991ee83445cec94c8e34ea8dc70f05e5aa57366b3585ae45e4bebdd048cd568d624881b2c8b667dc72f0a450b945f7f4c78677e5850551f000bbce5019ac2fd375b749565cd0829fab84512952f79d0287c327fc4ca1de2b6594552350a7918ab4e39cb37e63ac8163a5c8b5328;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h42ca9850a179de406564334d298127fbb5471e791b4ba8baadaee84cd7db0f80676fe178bd0683c9a3bd58a1e8eb3afe339e5a14e1ba924f1bd51bca336084bff39ef392885a40a8cd469afbec4a7a34d5450dcabecf61047fd0d97713a0e19abb8379ad07f43bc87d2f9b188f04eb43a4896f1cc88dfc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbec8ee74e0c67652c43e3ba3019b74e5af45c90324a511ad95a6743e4ca530ab0193466907f88b5e36317ad067a3065ba510d93df36be038c1bcbfc9117574a55a0839710489b025242e99399b2a279151326e5a5a5386500f896cb799554d9048ef98277e2eedf1575ff400e0690505cd9bedcdf2ef4c6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d5f9157dc6f01461d12a5c9e34001f2704746740a101ab33ef270ceb7367411b893e16aa9d3741636a1d5dd7e7310b59845b7991b3d9713c0be0d270ce649758e5ae4dbaa2c002877c9b4d03343fddf6ff98e94609ee3d7bc659d95b60c2587d447cfd8d8cc05e58e14a4551f120a932e590d9c47e7c25e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1397d3bd29459961ef9acdf2b95276b37b4ffd961e794ea2189f501b85f6392c3859543594711aa0611b4609e5ad63259ef997e95f95f758e0b9c8c99e128a48ab8f0237abd751b09f3e40c0ae5551d466b5af8dbc58aa69fc6db5aac80c96da32550ab9d218609f620d4eb2420f64291639e7b81c790397a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h121e4159eb826727c4193f16838e67085222cbfe23481af310cea93fb6679b6022630cbeb8cabc3e9a29ae9f5e964051f186f0cb06feabdaa27fae0b6c786692bc03795e7736ccca72eb78b198134586061492b8dc222c8cb5482d8435292c91987621ad8d8b1d546e5661203cb5ab444452c04caecbf9a85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58dbd33e3b690ce9f8352f2d164546ab9bca35e9ba60faa313d46b52f9e6521378e70895e9e9897903a1ff034cd0c673b55a3a28574bcc0f5ccb614c8cd9447c549d11a9f640e49562e995ec8239221868a3b006b0e4410d607c8e2df992176868df0f6fd76a51e65ed3ef596fdeebb0f85478b0240d3dae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c5b9270885c2aa63e2dee3dea4096d791341f50ec19a263f37e84945fad84731ad6a492e21cbd24e1c8be421af88d626557dfc4062c67d088efe97361a41b6a3f4833671ec57bf7c89cd389cc76a78ba96614e1c0fcf9b675afe99ed3fdba05dadbbd4daeb119a68e0e73b08c50b7a0c67bb7685dacd235;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ced28a1eb7d4533631391d0e318ccb990b4defc29ac57ffcb4b2c43a4a4c9a2ce5d8c1fb11f9760cdb4f1a6e8973a64a8f33ed9957c07935dd61d2b489b626fed793acebd506bbf30107aec4bf0d2d29a827e81ebebb290b2dc8e5fea16a069b96230f5c2834cc052c118efcf33525c15141094037b9c8a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h91e217ba3809cd1cb4a6920b3de68785cb37f28e51684cf77bdc648162fee7e00160aa2cf99c54cf2e0b1437a64199a7cd4e25f17c53ba8bc7dc3f079260fd54eef899815ca55f47a1361d8d4f5e3fd3a6cc24b98389776333ab961cc4444823601684a534c78890919dde5d2edaaaa5b39e38823f35b6c4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d43504e88a57949c3390fb58118a33ce11362acdb49901405ebd8fa7dad1805cd82fdc7aaa7690e3b4cde0ff22eae83b1aa608d22bb60078f01283c8092705322013e2afb573837420d88b16a9cafd0f47c3f392156371fe6e0e2b30a10b58ab706132a8cd7b3614b36c833b0034df8a02d9e2abc42df70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19772b3e04d9d52984f5270c39a41c27738d4cfd1a2617b04ebe21bee3b0b6ede3ba7b63c443e82d0b0c7ed9eaa36027b37566725419fa0d6c681777effc7bd60f2cf186f78eceaf5b2f1c8ce857a26ff3d82342bfaf0d0d64866d5dd22507761a446cd88ab54afba301c779d3b8ce9b64126d4d4f14efc75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8215c4658dacaa4ac278dbf07aface2747c14a9ca99c7c6ec1722d1fdda4c3485e5c09c9157172034e21b8e47d3f364039d02b06bc57d961b6fa9b80f0634c86836d67b1b7192d76f8c117b62d3e72c670f23f066d50f9df3e14010e41c971692ece826b68279285bdd87c100ea3db782b61930421e63a4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d2da72e69550e2b2e07d0b2ec00f69ecb06cc341913144e5829eaab4934eae470fe0193a41640d5038ba91409b27276b019b84087560110cdf33024a05b61f3f72a0dc1edc50f530788b31d2a1bcf0fdbbfa26f38dda9985b2f90decfe09912c0a161cb0b29aaba64df6055de25218ec2fb0ae1f9c23a6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5648e4eb3f077efd439e7e20af3e403af9d76a4c542e9030aed9c3c74f55e0afceae536f4790e4437c2f162b9da0cb1de77bb113911146fea34381c2d84bf4814e6b4edbfbf0bf70b46ac5be6bdd77a7f7e70efa2d7bbc39ff2bd515f4636802897953c5ca6908fefd939136100e8c3f587990429463ed9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf91f2d4cd1f6020fb9e539ef935978bf0c5903975c6cadacbe6108836c557a8913ae5a7aa1bb71b3ba4634fae28ff5a568fdd2dcca2c9a24f7cea3daf70a255beabd517f74313ae5bfdda74542f0ba041b456dd6568270b3aee7778ce146acdeeb9788ccd4dde8e1be7a77d2693d789ff5c8100bd83fcde7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0b67538984430bc317cf69fd08e69817e64561c83689280115edf4cd551f7ea0df951d1f4adfc98f069beea10ddf8c0b07be452173cc47e50f072f0663a7558d316293e478d5a6d1d2a0f9310c6e85b204705c5eabc13becf912e9b0ed3fb1c57ae37e069b1ecd014f9fb78dd8aa4c800daf322d36cfa4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha126d1b2d00f71b86d02376db60ee321f9a0560307052106fa4ba30fa3f1ae4efef8c0afd88db2f4ecb0b9c9abd7b76957cde45ba4f8204542d22ca663470e959fe22de0bfa1c1633143b357ae8b7954acc4be0cad3f77b41612b4b378cbc47f771ed75e3097a996d36e010b3b79870f53215b56d1e8becc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113e4c473106b066df1b908426c066abe38f04a4e888a675229fe202786598da6ceca016c311f7de100889b90b2e458f8859c0ee12ce9ba6ca08ac14a2ea613ea6f613ed0b3b9061035d6f90e9013ac66e2b08529dd80768ee7e496b8183358117b8a8747dea2821384809f683dd01d81f815a3dc10467784;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c71343df761aadc8d3f180d7be420fc9876e5628ec94e0ee7f062eeec670463afd11b90b6d32abe008df79c8431a4da1bbc601af7ddfa1babf279630240c15237826ed5174b985968bf127dfdb46713773dc93e761b1ab0d15dc5001a866563a37574973d5ffff76864fdc0808e147de5651af735ac37014;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0b2eb0e7e80d159016c390ad6b7c81d04f477942c90d5d0e469f4897b0b16dd678028ec6beea3f2870a1e69dcc3809cdb22fcfa9877d027a8e77cc23983dae5a7642ac45ca9689df7a227af827fddcda57c60b14c5c7b7e3f430ab1910e5ac4c5ace601878298b3aba2363b7d2144307c79d229ad47b9da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8a9ad5ca8411b3a89e41f7d9be8db2c6fa866b9ce1928700df923fb520a6f30e576fe9e97df1b309f669da3800fdb356e49c7fb927ecc6fbc7e9eebc9436caaac29fdfda67bc505ebb5c6bc704df9e45158370081b7bfc6537b0ebc822d28729d97dd8e11698a0af3a5a0ea95c3c4c0ee8f946b09d9439d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9bae0bcfe0bfc3a3f0f08d43b249f1c2d323e1519462bd36fc1dd33d17d87e6be7d82b8bcca89f24be62c118a1f0b717873e2c3a78104e1d2cf72e082a3a5043e56d8fd8e0b1a0093a76073b680b97d4cfd944f6102625da874c6c38fdb324c2f2a498ff2f7fe140fa67f7099126a362750ca5351ea914a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ca0e3876f4c923d7d6c7f5c0a4a149b742d4dab99a711230c47d7422b399a7799bbf6fb807df676839d35e218b46089452f118553054581e9a25e9373f90d9c6298098370e59f00f6206949afcee6ac78fb5bac8d071c36a8e612ac57da51b25c7a1ef9628e8df4823cd333a69b1b723e5820693737db1d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haba463494cc6467405e9371bf06e92c8d51aa551fffe554559c28f39972f0825db9488056c3ae939e241a58eefb957f458e3a55d60309eab9af1490f5ce1739a9b04e6fcb8b20b34c761e7b5f558c62dca00a43631a0ab0b13226581fed63282f3c63c51d41653ba88cda2abcf6ed8ba9caf7016e4d006b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h537c9231d73876d4e17b2c6179834372e58ae8808deaed508899ef54e70d1f8be6eed6bb944c433186755b00b45bc6a95e9f8f0946774166b68383dba806b358ea108f9a0603d2ace91653be59b0562b6276cc6b47758663179250ec9ddb3627b49dd51600561b41a7f2c66dc83ba53364fbfdcf31a27718;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea5dca3e0539413ebaa2d259ee62382fa1b49013aedd07a31383a077b4316f4879671d2e9165f78f2e8cbd5638caf2ec71fe338cd7caf1f5d69605b99ef4b32ac67429b028fd1a0e3c85e34869b36b8811dd79b01c5bc4868f0f2439f3cf237615dc154058c0844220a4563be6258cf7c39e27c1016c1d87;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59830db47882b48e0f2448cd5c0367ad8e1d44dcc266b7b1c7c80aee011bdbc8583df64bb65316f78ef2070b4de8c7aa12f69afbf324ef73c37f730fd649471e5e99a69939937dc31c5133143fb5d93dcb783b933b9a5229d8aeaf7b6e04806462a851234de7fa2ff4b48ac3249968ded5750ea5d63bb4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ae60705f7ac97664d2e0caf800873b9fec86ed59e439bcf5a64ef1e05fb66f838a1a969444575e48bf5d95b68815b290d1d1e3cb608bc7e7991f97b0cb6ff09c9fc17dc965c0946040b3379f95ee484635c397d3232507ac2d34e2f69c719cd7ec801a69615defd81ac6d158d8c3f280df9afcb1c130561;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7cca60fadf7c70ea8a2b91e77937f3739c5c44636cdfb25c219758de43283c01baf009873c3d43e47e687b05f88b96f0a6fda3ccf683d6a63046e80dfcbb1aa856a5089d791868eff0eb071c921f2dbef943cd5f4b3542c2deecb87584848387817050ccca0353e23f616716eb079f5a94e3bc144e6d3fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71bf9ec297bbfe0a06ee4504709b592f9ff58943d278db4f7fd1501c9303d545d57e36dd6d4688aa51da91fbc6eb18325852ded0466e58e8529b3f31e396814eeed528675a10a0a630ce9805faa211e449fdab2adcc081db964103633ab62d0f732ddbdfc08d3a6af2dab7096b19ecb8014d9d1d181877b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef70812765f61899d4cb97947a8a059d2fc1b26bab4e4c8ed3a7aec2ec2baf60dd6e5ccf2c8acdb7274526fa8d5b64373051942c8f493e442fc912447b42b7041280b22ff3e85f90e1e3f6fd5c81f7487c78dca027288b104b309b6a39c55f37853a217aa4b21f5f65025d2f8f7f7541a0b8cc2bf33a4c0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b87d4bf6487820a948d171b220569e7705cc143cba41f8a730442b387abf4862be16b4234334618c75485c3d38fb41a3479119cf9ee3368a84ec9c5e8d3b4f1ecf413243041f685b359ebcfda1aee41011eb94e20b545482991a72a1702ea9d110bf931a795e6cd84f49fa01c139cbca73bb7c709eb894b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8748fe18205dfb6eaa9adfb19bc51313a6c09cfcc5d8eafc186387a4a3c4e41f5a4573999772bd209830c980a4b8202da84087d2a16006485082ea68a5bd384697e632f4c04c2fd0a386f0edc53f91585b94ed5f72e6c152f1ed1f9b5faffdb30d787e200bc6777735c77800bc8f65271421f81bd98e978a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47ca59995f1af322141c2ddbf92274b367ef3ee32a376abdce6ecceb8bc4d0263d61e5b84ab8d1004aba88af8f116f3ead36ad054601b911f3f4d579ad5ce729d612517a48c6e10a26c84a7c32995bd2f661d46c64dc3d12cc0b1c18ba6f04ce3c7bc3058e1164f85faa05ee437cc48e73979c0c2a790f3e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12a9f0ec6316d7a867988762773da97ea08efaa6551f281057ada134bc9cf3c9d88c8af97934945c28052b4136416686fa61c6b867c64897a4a004060c3135fddec491555b05a3c9d36106446b51a3c8754e112aa4091bc0d85f436bb41df0a556f1f181376897f29a3cf426d36b3cd9e5396e95bc8583139;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63f11bafa633f180665f0cd5150d7a5975f544dbac3a1b0b23edf06eca8d87a212fdd9d72880166d9b6d8cecc31209efbca39af036d9d7fc3d116707437199d4b5452bee7be92588cd3e366e299525f187e4b648a4d91f24ca9a426ad700e230b1205128a4a328c2a86894172fa3a52c91a25623742020d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1998fa30720e9a01bff92e233afd08be53ff20f85f09800ed177a2715bcbac722ceed53f22394c002310152fd9fe9aaa361c25b9c726aaaa7d076fc431a5d6bc64a58c808b494997066912279eda7cfe23e2acc55eb75269855796c80d2a821a6ce13b29f0e003dcc900f90b561c8fdbb9e65f01361e94ea2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e63d2c07171d0a8edf628f21fd0d901668044ca4df78cab6791fada9a5ad4ae7060845346cb7e950f4890e7962caffc1e9226884aba7012d177e418cadc9d89450d715b8c6b475c6aecdc708c6cda41d2c525103fdbdf6217dabee45e1eb5f0d85d6c01343dccafc34b437fbb5f6939719efd35cfc7a4a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c496eed843b13be2b091e8c420fe4172380ad3e55344dfd470a91431a1612c8f414fb50d289a74bab990fbc7e05928d04dc4d4c345356bdb968855afe09e6392639bef11ddac285c23dae010ed674bb3829fde922612fdf691e9bb00975517b79f83334cee185cf70bf977f40f83a9d1ec7ab27d1f23f03d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde4535f3ebe5da1fec055fc24f30cbcba82b91b44a72ca2da10c4cd404490dde4b9618f7edf05a8d1aa992731d35d6f6542fbcbd0c237cf76e52dcd4b5e7881df2c4b74373cc6c2d269ef20bcea9799f2e69213b0af81e715d42562a76a8fb86532135cf0a4d0e2816fc1391f6b3b5c3b59cc10c77ff0b80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5cea7f715f09204596c0f5a4f4eb0aaccfeae681e809b987e1bfaae79630f980deb073f9f440035bfd4d1ad8ef893e698bc27d405d9bf2c625ef4af60d97862fd3a47a8e4558607b10d8eef74832e194b509f28a1a4aa30c9551bd4caed6924ba7d8541e606665fa85e2a18a9e357edc1d2f7464c7003da4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1daa258ed7b9ea440c3eaf4f0bc8e74204249b23f1e443921ee1adef571a71afd2e29343aa08d3abc8d4460852712115397d7ed16f493f8d430eef282ac041d894b5ea3f3c5edbd6850683310780ce8a16d975b4ad99fbe198afb782fa84d397afa8a107ccb10b4b60db41684f2020bebd4ec15212ab3fe17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c62b8d37ec7d96fa450db52389703084e0accf06ebe327d16019af6ff10b6cbe94f715d8f7ee8d0429d38279ff793f5c6006290a236bf208356826ede4d896c1ef00edbdf2d57fc064f4d5ba27b0046c0a49de00888a8450f7b9469d099e151ed9394dad5fef25c95b8b20ca33272448ccbeef762ae4132;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52cfdcb61b37ebb7b183cb070389ef10950e2959a9d548ee240c47902e987c9b6023447221a8062eaaccc026bfc053806682f44c9f642b33b45c0e7069ea782e9a125ddbb06d1dbc3ee55897f1e4e6b7616b4683cb967ebb49463b7b10edbf56abee41436c203417eaa37a07f8f53bdf4964049e052ee51f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154596d3b28d9d94858a003868ba27eafc0724ebe06c2bced0c4e55ff132b195469787b0f949a3c3768f035dcb59ef123049b3be3a2d3142ed9ae02316640454cb3a5cc7d061bd55a9ee3f08183ab30d1412e982764dad14fb9acfbdb5bcdda114a6405bc1f41020362483947a8bf626d4deb9b403f765f9d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1300f2906be19eba29c8f4e6f4e51ad8a326c24a868f890e68c8b4c8497803f0e9203ae7472a33b39564bb9ab0dfd62d84a5e5943353ec71bc08290049e0c1e0123c7d0a31239ba96f755b0aeee8b4da5b21785f3eae019791bd95795da9a17e3449525bbee2f936adf0787270e307dbd91f1e10cde05a3a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1de928a46dd569e3af54675022351212169ddcf324d05f039b9a7a6c8cc299da397bc61d1fc3dd3582a77107c26bf11d5e45d7c90c626c2dcdcd5f117d2aea5e3101256d27953f4e6ba3bc493b7cb0ebd2dc5c497051075c273cedab4105a8866ac80b6007d3111f9719ec69107335234b0789f2b6aac2599;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h297980bcfa6b7511de283dcffc2494c4119359242a6d0c15ee37f94a4853c608d91dfebe3dda0a3ba509cec3c2a0436b8fe84b820c20344cac2b8d3629b447e9abbc5a21f96bd764a30c57df3c1647944903ffacb8e3719d7d10cf8b12906a18630391341bd6ef56177294cecbe9e42c972577c9c144ca57;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8cc8e3f61b70fa3c303b68b48130040b277915bc1a09cd7552e646983c0ae8c9daadc23fd4c267b30ceb0fefde59316d698d4a098e2ed3f34454fc308b67e961dac92cac9d8d27e5fc8a4aac2e146ef80e666e78b4969094c1279cc93a1eb7bc754a8b1512db5aff9403f7b768169ba09ac037fa12cb654d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14e6588ae594fb771229e7868f0305df29f0a25b599dc71a5e321f078a2e4a98930f92192fcaeef1d1cb7d0b86ac82dc73ac6514ab1f5f9e85e9d65b68dcbb606dba684da233f00b0805fc73ab2c481c3e8feb4f3d6ab4a38d58549f3e2c8af5e787b713d4cc1e2e7be6d3658f993c584098bfe0e3430f385;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c185e10f6938b001b2236ba93dde304b6dca2bd56f50ac56292bb4bcfd5ed5fd04ce5807ed4c393101f5e9091907f3cd6e2c7c351bd41641ac99d1aaa17601ae45063f9f600213513d70a186f29d3414e69919b8f55ca07de4bd0b752c6edd4673abd87c13a8e07f178b000f020d30387fad5d90bf0a05b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59c87e3e746058cd1041405688f5488158301b228421be4582209f70705f506e5f36ba7190ace988896360bbbf261cbb58c374dc2f081b94a825f2b143d6c1940ad8bf4ef5c88928af51a67e37110721f4140502b22dd61522740affa615eb09a1b280e8f65efc38e5ff76041602153937a62c3e56bfea9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1feebb06bd3896fec20265e6be91a73cf87fe417475206f42536b2e5d0e74470454376bebaca8aaca33b9ed93c8c308de226fbf6118e8649de12e38995e191709a7b38994429102ea4b13f4ac72533718f0b8b5cb4b454a8a302909bc9a3ba7c377efb677416348d14e9ced9e5c05cb66158ebe37b4c5c6dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a8ffb9e575229c1887b6c16e37f5d32e48665a4515b1c9e6e54d55f61c42d4f653d7448b81c73258de86e55a91d6a591ae7b74bb2df8676deb4ff1de4b1aa04f02d5e99061e4fa5d1625e67cdf89948ec760557aee9e4972633ed3c371e53776139a7a985f3d38c48c3edda71135fbf7409a455fd833608c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc7eb0ffec8172c53407081634c2c2c5d83f423b4631629e6c262c85409a30fb8d00c4f5d2b371e613979e8d74703536227166622a3a091c29b836f7facf3bc2b6e915ee8da3813261f6203548a7a81e5cb91d69501f16911db8446c25ef745321fd767e11de64190d7f238c1c0cc02bff223159f7a8c488f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec7eb103ace3be3ae711d25767eef8c8b4982adf62f9475f4b9f321d4ddaf0acc129bf1f3d34688e1220cd740b19560883ae6f838c42ac64dcca2295096a99bb7df85db1470e9700ba78073c74c9477f19b1d39d8221118c156200ffeb12eec8ee61e0af91740011ed6190a12ae9168ed21b826bce9844c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d54d3660878f449c43c4bbb8d8fc353b7d4059605551ad2a7f3f436e613eb15f7940354789e6eff2d7c440760e6f7b510570856cc9882650294e6e7638654e4c903ef0223dd923c041d55030c624e48ffd3c95c3424238358d56c52349e5d380a277333821a3729978e43f247c665b7bfbad167af520276d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h89b18a112ff98ae4d827eb1a157e96dcbf57c3e55cc644103385d589fb928b1b46f8832d36bc30047382c05c14e80f59d53f9183072310c2f7013ac70ff9d4b40aa3dbc0be01e84d744f81c4ddd1ca23336283577dc59a5a4ab55c6d299612fb01ea74d864d43b9345c641076bdb16055f51f914015c60fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1054a663e250c1cbd2ff22ef1eb8869cf3e8ad5ce63772cabf64893aefc44006c54244b0479bf7b29d5ef0c41e20088f050dea6be69d33fca3c7f274a064fc689cf1d46b5717036f8980b520a7ec0b4a24c048cd9ba28b447f9bb29394295a7614200c0a2591cd86d159764cee0fc67e849d9d6d80a9997a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h164a4a6b17cc1f1e6b8a6ebfe4b05cb8ad24a264c03b791e053b993c241f05dc86601589ebfafa2ee916bec179e3a0236e698426caddd0cb1b99a420c499e5d4623d8454d2eb760d4f77dfafa91c404f36bd5be011e0188d7ab41428c7223682a1bc5b6486bc1017b9f00f8723defb8d149947239e5879fd8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d5615197eba25c3415645a9f7d15b9891fd7779f3802fe86aee5a2b4793a6991a226d3572d24e9870b25df9e19ce1a1c7d837e94b11ee54463995223a2c318f48d2fe0ffd13569dccf47b5d8977990fbab32e89b149b2df2b67d0dd8e91e6551f4d0b2f822a286bddf9554a560690a21f3c50649da4824cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc57474a5989099ba2cb0fbb7a3f80fcd85c270d98ddb22abc6455081a3d52b92be46fbcf77f703847d77b3880d98baf4366bb3b3a57fe419dd28b1624a7a676529f432d2c97affcc387633a85a44599cb5416fd011c4b24bf9cbbdb9f843bc533c27c725578db4e608ce31e12d5a434ad5ac36679638446;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f72616d18376bdcfdc1c935c07c9d4b882d00ec99190f185934421ab19ea405d122f7af6461a76a9926bbdf10e7187865d70245330483240f038d34a85412f95813c7fdae3e5c4201ed20e083e8582faf8d9a927270de9439cdc5bf0f93979dd906800b4c2ad36b522b82737335dc20e1eef6726b25da54;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h533645f192f5372ebe24a4132ca77db04242dd7cfb5f56e9b634c1fdec583971a07cac5e6429d3663c150ad24114ba9f2a6f4f30c7392de1ef05493b76d529f96d404bf2f8915cdb552e3b41ceca8efea1ce92a4007a111fa61aab1a8ad27bc174b062da2be1ba05b3c1bbf6299ed717275ecb0f8322a628;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e321655add61b52f88a54b70f31f6157967607cd8d6947c470bbb32e5a63a5bc822ba3a15a1b030f135c40ffc65b189ad0c280c3b81a9b5823732d1e8f3c393428714e5c06860e7597d7de542f50b99d5afba06726d058186486b9909997d8a181902caaa3341a6d34a703ae6375f9eeb1e01b02cbf07338;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1970eb46469a9e53697d918e4fa64840949fe54f0e5b59f130b1a096e69fce99a10d468eb98e96ab73e0a4a6cc7846ab0c97622e4047ea4c8a6ddc77d436b9cdc77a03458e782ad19e84a6eab0d88c2381c1cf4f8b4fa115ec47f492b9982da37025ea55b33d13826eb44facba6cb1697358055e955ba28bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6d94927e5b5e2441654aeed55f2a028f4aca74c5a69ba69cb4267e992c084ebbabbd80247283cd9c2820e79e694a23572a963c12df0b1717bf3091990f505fa67f78b97d4d31576f8dda123e2d27858555c9cff24f53d5b7d38325af4ae81c2083e9987dc96e09f6d15a815a60c60c2216bb36dcc48e37aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe105c49b6451958291ae4d2d72605befa110603407c4b7b2a81ac51de76414ef8415ae63f874d988f7f243b3e5ab0c8cf464dc3249f23ec116401ee90ca503f3d99be7f14d953c943e622742345f3c8350c49725aa4185edac80d1709b0b5053ed01d63838d0ea91422eaab69c2465e6b39b8d230122e21;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1200e118de47ccc792029ba110a9d673c3824799e3b7e887996aa16299d865c60635c78738c1834b75e40b7fd36698ac14d2d846791c898e98cf70f6a253010a9bb39f0e78f5a481e0c47184bd5ed2dc14ed1f40e95ba0ecdfa1b8538af7f542644073f4fb6a9cd7bb6cb93573452a3423c968e8b7bd0536a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176bccc4cc670e2c16c056e4dbba8e8ed01dde074b654926c5d5075116c82babe7b95bce8435339ccbe739fdcbbf66403f7b90835b9be46b46e9479f94ed7b077a4c40cb5c6f0a4c95b623cb0b239d6b8dca073f1a2a6bd07ff055823784be046a3d3b1955d259fe400d44c59b667ce368fc8619b3e72d495;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h803ffb404dfe4f7daae2eeae861ba9326359195111a888664f5c77b7e6d160c6a920e164c9d4a7d9339e31f3e74a50b41e9c60df93210bb027fc712785ff40b21a625102167dfe9c753ed49b0270e3577431778d227ef9a96aca5f3233eac9fdb06deca03c5b824eba17f6f19e7a2cf9a91b30dd4cd32eae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d9491b845d17c9bc792df2b384620d8d080247c1f3f034ce2278a145ca79909fc79d959c3e1e8ffd2b2343db8ac6a4d898dc922cbfc1e16ffa5376da4b948599db8e01314f7480a86ac3b7eb47b743ff11453346a79d890c0bd9334035b1b905a801dfa75232b858efd53366e4065adf1217be8991a033e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h80a01c2094b99e9a50d0ff975d35214067bfab2b216df4b1865d587c37d366134271a05302c3556f7b461b08233ad891aa56defbc8e527dd66d2fe066c3e710cf359b2f284a56005dce904ff2c6fe7ab1f19e969c761434021c7f1bd05d4ecb8a709aae008ce1f9a6e339ff4ecd63fb2318366ffb4b111ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18277ee7047b7e1cf44cf99057b8afd9bffb7e0ae750c3f6c1d2eafe2a42d762e5d5c4f0fbb8e3510f89799ce3f75b05adf6ed03400dadb3db0a22abf71646c2cc37e339a5b4fd2e9d1df739d97385f4af54229cf6ce39a5fbf1bed878bf4634a60ecd95831c29d9d349ad16fe12dba355992b72dc9105d62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b17beda12feb784510f587ee0a83e264ab2e8b64ac73083a930aa4dcdb68d59abdeaf60600e7c72e633743d26db77899387ecaaf8f8f52b4ae01ed50a717a7eb91f085a417012cb201c1e8c8af682942f5c244147f7c08541f3f0aa730325334bc5c50e594a94036cb0faa1c2a3cda66ec8ed0f04b6f41a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e467f608c112307ab1874fc0618d4f4e49ddb01ef64c2b8c6bfc5e5f7384a290054fe710b85d5157e0f9d9be76208d7105a83c52676b937edefdc6777bb7b6d4aeabc6b6bcb031ce57ca3ebb1f7667472cb1296f649d49fce8b06e5a0996e9a6ca7acb8fd8b57c1bbe9a5193826e76fdb3506d1a2db67812;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96a01549a6e77b59d646b1931def82eb3d8dbe64e5952d36401f1c64058060b5308770c89eda387302ccce4970162c18cbaa52588c02848da4dca2d3582445dc4903112cea91fa99eae9166395f39aa5a15786372bb13fdc2f013a6305f4d9fca81242a2fefb3e763629c3089f4290f528b4e860dd6a6717;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had8e701ffa22e239a7f0c9776fe7e46e7ba3be4cc42c46de06ae751c4126b795e036f68cd2e138c1f28ea4ce396217cadc97a9842795109ed15d20994049c2bc776227cbc93bdbcbe3f9ce31178de8cc35c0411f885a339ad9a3922a4939a5cfa907ee8ef01e0c1093241b1884748b66a382a6a00b5af87b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1925e0337d94412067bc2ec0d542b4dfe78e265e54018ba0c09f822c4234e462d389f4fcda8a9fa4f7656ad0215f6ed68a5d82c3ab921b984f1d91cd8ace33b1a7cd625db12f7d3d12ee909a51aaf1426a3a6e42d0b9e5100a5f80dfa67d18d78e881a453ce9194bfd3d51a20c63d6015b11e0584d4603f74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13eb926b5301e2e32f92799def0928a3b8c5aa934465dffa279e3b425ba98895f5d47c7ec37bf6367e1e9b68cf1f47d3718a2e505cc6889bb3b4f113a75058cb442ae481015483a710cd7c6d8bb2c951b5b494f2af319f494bd7ca33f797d4aa5a57541259a2b9f68e94794a3fb17c9c7874e3af52a246c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4dab08f87e050fb916e322041bb83d9b70d52af98550a830b8242ba1e51f38dc16fe1f876656126f02ad4eeaef48d38c7585cb02aee789d59ed5dfe4e92078d582025f8f6441cccb94c2a93abc961fc5abe529d495c0dadc98a4c246ef703d75b8259d9058914b85f77f994ced284649154a5f4476e51def;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49240f97961dc745b65d142c97f2cd727f7778b5aed3bcf5e1efddfb7d4f0eb9bab2587d4f0645e9dbff7cc71b05307f77174f8eac49f5ee5591cdf2947a6332e671c0ad52f3bae9cd0f620cce90aac7f6f435d30996c700b1dfe8961d4237ba2f86c59b7c20246619019648659685417a5ef58517a87d22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ed340f8f72e8deeca916eb89f9804a1d80241f84cefb0be9b988cb8b2581d3faf55dd3f47df7dd1a565a6f6e793b854a3e534e334626b27b45c927b92116cf9dca9c0da9829fe12a16002e1d80ddbc0e58dca2af72a54801a29131c1d54663da52707a5f2caaba1bfa6c1a6bd5c79add99480ffcd93312f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4eb19413dc7ae36ed28bc9416be663c9564b6038405d5208351eeed548eba03d4059f9cd5b56195d04b8a95dd44fe0eb0a26a215608203a199a0d9148d5b5c43af2860ad4771da5d23345be2f2772e32a9bc4dff4bdb2191be8028132020a7cf672d35053840552e9ec1a8c8f684725db09a92c8e647f8ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1131c4b868b0287519d4b45ff036b3f563d37d6cc15d1c92451fbe93f4fd8b61948aa6d1d64f59fb9297cfdc7efb8643d726e05d57bce6420405b9cc3889f1090cca95c689c89f309afe3b8b9894f2248f12ec75aa4175fbfc7b84952e97883cada5a3815d860a2cb78a0068e2d7080d23de6bfb106bcb0d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c86bcadc0008f8400155db79a2b1649fff36a6d2925eeeed7253620ca7d7dfc29d7423aea55fb05fb6fae16410b5e087b4e818af0f4c0ea80fd0184d577c7fb46202b082b2737c1f8ec0688ca13dbf55fc83845d1c22ec7d493305320435eef29c756feca98f6d22203d6f58060f3f00216bf00e237d27ba;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd53a245231563f7e7e065fc7bde86b90df1f6ce9f9f0c34d48b9f34f467105ec41e2e1a0b81007892f93bb8558dc41a9a2d3fff6ab832ee93b18d1f18b092dcdade4bcce379debb3b13873976b2714d324d53bc75928f64c024d27506d7ee222dbb280a96b90eb383af779a1767801e9a3b366cef25bdbed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12bdb044d9d679eab0b27c9f50c5fa667395d94812e3507e5cdee26bea3ce6dc6a93d916723d1d3cb523c61990f39d9127faf64f22b207db9fddf0bae0912db56b4b629f9b4cdad7ecb4e5aa549a7034424a46efeb6d604a4222d3a39b5482b5fce90750bfac09412e9cf1b42ae993d05c96da451f3d3d40a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68af4fa65d2156e13ed34f0fcaf6917eebf65debf7909b33666238c0dccd6cbc37045cfee628f3b3e7ac4d2cc79c741e5650de9370019e38c5d6b7ef561d049b8b331fc71af67d01db38ea5adc4623127760324f6d68d15aa5196b414bf6999709741fe81ceeb05931c712bbcc5e8f5bd39b86d10e8a7b09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h48793aaf7a7d710a07c87ea08e00f93aa9e8d81aa6308db36de7626ec183895c818023df8a5c7ee2991f0c349e5228378c179708f1bb3c5c66a1830116de9a6cd2aa7480e82f2bf982a6a2a71aef028f4be7b53ddceee5dfc63aae1d1a6fa6e412ef1cdd64de9d6b439f8925f594df70bc9a62f7ff942eeb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f2cc3651407cbcdb1cde5f2fbe19c973a46fc99f83927969418848c5eef72d01d38aac425722d296c321570596e4cdfbe4b6f350d5e2e68db95377e84b892879444c19a5eb25b939159f5bae8f18f599142957a2a25b814a1a6eef12d6c97bbc51821a30baa676801e59412535b527cf1653d5b7b415376;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h758ef90f43f7a28feb5ec10224a842860d08f82d4322c4e6845c21f8bcb427a2758df116dedda075b9ba2616074b91145e0b70e87447eaa211c52521b8e920573439a439b7c96c33275befefab16f1799b299f1d6e0cf966c3f561d291cbe61ec60d6c6dcbedf8bd49cbf375e7c81c2b97be946805f247f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0af60551caea803aa301e3afc67ad3324757d7808bf53767306fabe7d303f47e72a5a546c471a8bc64eec189bf5ff82dffc28b74433a063248a29ee93df3a3a2616fa989554555f1e0a6eb74b3d62ce9522386f299671144f619865bf890520e19378ac45be4ca95efc2ae3b3e25b3747592f3392cab871;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4ba97d3b9e61f2761ce179efeccad41f6f65761cb3b823d21b96b50864e997dafceca6b853369d4bb5b8e25336917f5b7014d0c38eeebd5d2b61be8840fa971cdad9ed895a5dacbfd6fbc31447c2f68077344dd5b70528b3498944e5056f2121e37be6c7c2716585d1035ee66d1669cc632652c146f056b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h126b2b14e1bb677b16de5dc442d4b1be88d1e3d880eedc4387925f3fcda7c541c9b6976fc3a820697e92dc2afda427b7c7fb11ac796a1cc394d2a76c13ebcd04a84d6bdd77c89bd8b5e0c2037f8148d8ec7fd028598fe23169c16469781b80ee0ad48422a049cfd929219c742176f09150ab475465c2f621d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ff4515fbe90d0823f1d8250723f6a3168eb0da32f9467dd32ea02a9fac815326c1e2bc8eceba871ac51cdb72fabe3b6420f349e8d62a5245eb69fef35b587719ebe2975f7e2fc05dbd8c73399f33f18330261a629570a9f662864bbbafde5668954dc48bc741605045bf64acd3d0df9b1e9f264c21fcad2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19afa6696d50113ca20282e1bd78ac6e6b3272496bb95872de51e01c3b51b0338ede8a8ec6409518a9232ed2994c495abc1bc4cc7d5d2e6a0c789eb9f5ed4d44ab5659f714181c25e7047334252b409c28669e887067b917247bd7cec13a0158a3cde5f6eac70861fc0589fe05a416820d27a30d40274879;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c63b2213211f5111f43a86d7202f913f9db1f2a8b19b13cb7607709f6d836e6f2cf4416ca31af0839e4b19a813b353a3cbf7590f93538569e346fc5c1268c7b767ca408570dbbef7f4a384b7263b7ce1e0e86b9c26b532d8d36019c073f50cea88b41e791d47d2617ce00626f5e903b37d91fa10252c64a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104880a5db9f7e2f44e47a51a659eca1d67cf3d11eb4287bd0aac1398de96adcdf923012c144b168cfc34a5bcd72ad36cc3ed2e516ad694cd707122b78b7361d311a5d889ba2ed7b9aa5bbb99e39fc75c1288c9e758e3210d457dab616ee8cca70ad07c0b47cb7908e75ea7742c4b1389d9c1d0e8466a4b0a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108201b03df7f64c3895db127bda3c70282ba5b2c7ecc5b2591b69f87d0fd76c2109686d2381946c4f7d4cd38d230700e6c23ccd3c10d7fe86a3de455c61924a61bb49026c9929e0c5c0949a2afd029c44220327d2099985167c768c02ab52789b9ae63605de6b35c9c6401fa9daf9d82608a2b5336ec5743;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be9469da753daa0eaa665ff3ffa18c74be12180caa0bbeecf174607b6fb954e3faf802b542585b10781718351ed202162e76ca77adf4eb8df5b34a7bfd826965d4f1f7f68f2e9737ec284f5fc1c97cc47d7642b6f28bb160ab828677593dec4180babf246c2485981ee5c0fb4fc54f4cfd6f8e91fbd22fd8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18bd6e8efd778f58d4deead7d52bceeaba45fd1e1ea45926fb643144bf2fb8b62ee3a2d09d65dcaeeb6b0a7e18fa326bdff4010f12538171f0a1bfe12a91c3f689b30d4ef886f6b37902421b58ca3240b23b9958300bcc94cd1c864ed2bb70af9c529aa787817cdb592d5879df4353b3ad056d6ef6be3aa3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16424608b0e2446680f1be69ecefaa7580af15daa8df638c1646825485cb270dfad091d70867a11fc0b9b2f86217b133734902c679baac1515658905b4b4f2583f7abf8114452ab0c0497f7fa80de4d00efaa512b41100a7ee9fd6e3bc79daf75e832b463b4ebc44d41b4fbf75a6a89ec2b1094ff2dfa3ff9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1acf33906def0d558ca1322d93e9b89a73e2ca249847328b0d31fe0eb1b54f3fb1192206f2eaae1b4199d721510fd43b46c04cb2f39c17b7e8755b6ac2957fb6009250319855c12a390fdc5a2792c22bd86e370a703e541d5dff2764e937bb3f6f5358ca5e25fe7ad5b699bdd2e4d93265a504b6c40839bbb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2abe1d359bcc708863ac8f83791323db4230f4b1c2a7250f2c5a16cf5155ce27e9402ee8db63bc7d230871fc098af10acc97b168906b83d5ed0be7c2afb23705aee9ba3f9a0e299b3941c265af2642ac4c487010d51ba3113a76d601e606d4d5b2e6d37f21e25dc61b1ffde8d8365a61e52cc2ec4c180f97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18489a65aa0b43437360b63e2a0a29e6b3d9f9b39bea594345a6f46ab34ce1c455393437de277ea546f5de49d74201e3f318ae893318d136490f9256703103c90383aa2881e61e713a22b71ec6a74c7529a1a324d81626db86855f27edaddf5c358eb4a18996a9234f2ad501f0a87adeb2cdeb86090879b41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb08ad1623bd118a76ee3dfa738604c37a4d66e32db4fb208fcd4517927ae761af3748e17522660d1b6db98fcbfc950f7422d841f63dfe4ba9b5ebb315e61f4b32f1822e3ef3baa5ead7ef4f58263efb03deb03c1a9aab55386aaac235d46aa20ec46ac40769a644af9c3b095d0b36d941f5c3b96f464b470;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc48225cb70d833d460be23da0ef1f745a19a844ccfd3801cc9635884d37764ee0c9a5cd584b755923d8ba397e2b9f700111992842a8d33695948cc3fb3a6fa91b117c70bca4e458a372b44de29abce92ece096cea7df0f8645f7ca26377809771db8d34e47814936984b655be7377f0a815e92e87c9be665;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1977ade7cdbc027e9783264f19774bbbdd84e375a6bb445184609ed0ea921fef413b37019b070f114a261e5bae177743761c558e8bd86ab4d7e3a7875eb227c5d29bddd789c9c10bd554306ef26b4d8e799af0e50d7cfb9d8b89d9b41f39fbcd9884cc21aa022f9dab3c13f4f6203b7a1076df85caf384c98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e5fd83ee968f7d8a7f0d173f2d68e6d17ef7aa053bbefe582b7e0390d766b89885b7a17892b24c73887ac0276b67bd286800ba6b4f328c24486b376b3b71e2b6d5140cad7cd379735e5fcf1d797f146b293f1eea8aa42b17eae6883a6de42928dc827f9b878b2ad0c622524939b81ca11ef2a6307dd6b45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3ffa4f5380c7413b22257bd2cffddfd092a6bea2cce5070bf4a44d0f02f9bf3b62dd98c2e1c2d529a707ddd782f3b47fb58f6676a21ccc6c5af9cc0cc5f9ab7f7635a03759f7bb91e16b4463d4880d02a4ec896518949aad5acf0f4c9a66c690a407d5e748ad9422cc68deb31d43c354ed05b352bfab2956;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf27939201ec6dcaddff39d881142f5b707a0756bd052e8ef4180ad9b99252536e4f85289d38e5a8231629ac6a95dd76cc9bf5f2a5c1797347c1c26b18531c30d42556dc41cd0f605f96a90943d950ee05dc09bd270347bf9a92e03a60507dbf4cb8203e58ecef0172b6dced3b8903dcaf5a900524d4caaa8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d0073a80af1ed0f1784f48003ca90410081be366031fb1a78d178a6ea24a9bde006ac4b63b5047b51184f8245af2ac5bc93026754fc3bb160913ef687d0bfabc7264ca7661145e8f6ecfb6ed9426e4dd40ae858f0d7a8ea66e90142eff472908015552a4a32893cf0af3a2bfd322dc0d56a04e4af4220ca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d5acd7bef7099d0936c33e9e44087b0731ee61246c1c8ae4083d2993d5123a5edc588d4e51b894bb58664fa10853e784464069bb087ba5d46767eee58694b19491b3f9ac8d50a9d59e8b6772b88d3f976f7c334f58fef86f555b67c33de7f9a7bcac1e5b791f7330c83c7176eb9eff6b50969dd87f2af28d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1707a1ab4defffd3dc666bd0ac392bcd1c926029860ba4f4c9c4d036213847e2beb5ba59adaa360fd5d0db32d1dadee2752b65fc27b9ce05bdeab405ed9a1c7190ca85edc6220814504fc5fcb417cd23e98d94d618f78275d0e7c8942159469bdb3c9645575b5836c5c0e3349658182738cdfa68a960d5970;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h199b2fac2e9369a28c94114f129c6ca8dc62d21b0be992064aed852b717a001f5a863a8e378cedbb3984534e78cb174accaa741e2ca3420c2aea3e906b452df794b2f5adf929f6692a2637263f50922bee660cd095ed0e5ace4d0fbee90eb9d4699b13e64402f4388b38d0fccdd98cd405d127a68777b328b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cddbb7936e8f0983bfb26ab7ba14bbbfa4fcaa5db7600f7a9b7b2712bc7f2767a72694a3794df3076e586cbcf916a2ea59cbff85afdeea31529545808179b64325bf1acc69ab85de2b7c9e22489fbebbd5949e2652dcf4aae9f8c3f697459c1c2c8885dda722458b58883172c1e80b5e1a43e3462dda128f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78985b2161fe1d3729ea2cb054f6d8105e38371a53c8cc16c208c3692a28b7107a62640f54ed227fac6619054cfa2b827faac2b95736ce12428c3964f80c7eb6cef5379b36bad79584f89058462760f1bf0e9c18fd5c6c5de0ddb557909a6e7086042a3466d3ac5d9bcf9324ec2c6ebd47c70005d66f4a71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167f7332dc5dc0dc4508cf270e070138e3f5a68631cddeb287fc538bb27fffe4f318695d46f3cac84c1ba3614b38a6f93c44a7eeb4e47a39cb71b2e16098aaffa251446fed6a93c12642314f280fba06914394ec61afe6c97412b8156a06831472f6a8982237451280e05c70bb98f6d4c0a8dac66e6526317;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e527220f7bfcc855e62bdbf4cdde362beeae01dab2a41ad8967e65f63d578ca1a5a9d8366d775e3c4caf0c45471e19120a9c9abd7093e52197ff21f618633378759c7dfbd64849bc113bbd6e952f292e33c0c3c2b820f28d5c964c84ae29ae09ca977609eecd8dce6a5cbc59cb3291bca86cd235088d7bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0b3dca20b684b7c1140c30b6b1d05a14c427de299b93935af0e0ca9a944408ada3eb3cfd4a591baad0833042eef1e5a587f515f9a78644899bc0c213f220d6144fe0bbebf1ddcfa58b107879be395bcc57ad425bc14076bde69256852ab66bca5ba196accb1b79bf4881fbdff8b65cc88a4d60eb502b566;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d45a6327f0c99005c4572e4ae7c0f558d5133897a0ce310561ce0a2ed81dbd61a366aa4d1c510a41e81e7d58f17dd8f8e74e57ee18cbdeae2f925ede1343616cbe987141a113c95263815c0ca376f7b64c7c1fdf06a1b873c8ef2a7b3017d7f950a9f25c79402cd44190416eecc896f3b0bbddb99a8da48;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1516132060f5dad4d32ecc1d9ae1f0096b4549296c40e389a3a245f8557b05a42fa5d193953d2a41098eb36841ec5376c9e3c1bfeb7c9f944c1ae7ede9fa5d321cc2bb64ea9339afb2f0e791f18e8109340320177c3f9e7799f6af5c66de62933e0df02710ca3f13a78b1f01f2547c55ca9e955bee86d13da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8a4aea109ac8772049737c593f0a6e56f2d1d8c02ec23198cb6c7e43a3b11b7dff4a2e60456d5ff72e0c5e5018d1835ca49235e057dfd44b8fc276695236b92e01638970908a734964d725479a4881b44eb706297ba5673443bc4bcdf8cfcaeeb58b09e11dfc91de868e1a6f1b131ea1a32dae9b2aca596;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h32f2688ec2ce5715a1c746310d3463a25c0fc45accce038f0e1bf6141d6521ceb984bbaec20cbb783b9ff6a2d07a460608af3e04632d7e61a05a4bd0771c3019c85fbe6472b024cdbf28dbe0418c0717c74f32c44e936018c4acc9bec13bf72c2d4b41bb982a96592ef4f21f7e4936f459a16528ab301bc6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0a865536480e5eb69ddcd3a6e86b2e7c8a1fdbb460df3ab3dd68ba0f219d359c990644b447a271953747236f98ad679d6866547e5194649e1f5f6f9c0f38adc1ab406f6f441458ffe362a6b0247b597895c1b37b79a70c52ade693c6a8f5d427b9ffd4aea17658cf787c96e4812d750ced39a068d17abc4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbe7d44eddbe61e5f07ced5a3e297534d4d870591c6ebbe496769472ee797cf5f8e523cff58ad5815fd25310f60960556d1b1a120082d3c4b5ba83cb026bfbf3b3b3463884b21153a5cbf5b9519e195564adbea93910558c6b2d4476d61be6ba861f6a74dd2fdd989ff2a28742911ff99307c25543b2005b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1db9e296c7a10ab677088e55e6d57a0955f5fc55ccb547f6f3f02319048d0e265a619c255f7599e402096e26496d3d9bb8e9727e3e412dc7ac602f73e6361e0ec1bff5aa5e11b0882e0a0b4d664c76a8e247bb6a2e3fd9157cd069b3abaaca46175e862f9cfb00b047e4546b4448affb5eef139cf96b07c19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1329182b550dfc5db1b24de6f54115150fbb2a8e97a02482d1ca9ec57d06d0e3e3648f622e2d4b316e4d7740dcdb84f91ec08c20a456c8e2e85c9cd40a2189fef2dda180148b2206cb94f774e7ecda8366a132bf93809641cef6ea45e7c014554c2e7255a34867d7b00ff2f3ccb3997b73c804018ee5480e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3239c9eae81ae699f96919afb4a40dc0d0107f02510424a834f9e538042899447c3725c8fce770560a25077811b3065242bd7944ea22a2b4a355ed1f5e0cc1618b61760c9eae889d2bd2e131c8986a0f2b2c3b12d69a8dd87f4d1445b4503e4f1028d9c0c567aa52bae8fe3cca147a3680c1b4950cd846a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e45fbc682a550ffd9193fd41b33ffd174e5f5977ec3f2e4a2a8020579b405df6f70a7001dffce316d068fa7b635bc2c8163f7e5590cc82867f173d30a0b4c2d71ec9519e717707c2029e94d348c66086d5bc5f0e928a4076854c765e18b4fa8489c0da8086d27b63621ac2f8ebaf5b49c3555f380ba0971;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16433a578343405151ef6d760634546eb8ab7d664243d8b64bb5431650468b0c22a63fb6986748ef2b18ff8655e28dac3d5e57be8602b01317424bf79a095a356a20838b12151c02d2ab21f52415b066754eaf15bab4f31978a156fb37a51159615860aae056a355629ce294e4c64eb2519d54caaa9303be8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cd2ccd681d50af39a706be33f2c1f3e929d8848ab7ed476b80eeecef4374843be4a3f9a7ebce18fde29d0915dd64439e990c56aebfa867705f5a6c405b2db096d0d2c8bad5914ee8b633652f0d675c9bf61cc5785c227f9480d687bd7a9d8197ad6d4abb8f37a2d2aa1d7c83b7c163796c15372af36602b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf59952bbfca20bb041cf063b2bd4531bc5dbd5d63481a41db8826f34a940002397a1461998303f71e8d509ccc8bc771150aab842beacd68842f9bc155546afe50f0bffba5846bb47538fd81c5898b298d286b48226d84faca1647f60fc73ef16a107d278a920743775a1b33cbcc7473e361c9b05752082c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fccca38c9a93fe7656860676dfbd43a0294356f204c0eca1cdf15d2d6b035755d0ff4bc6934c68df2969b0224193e0d9433bd4c66cf14ad69dbcfe0d714465849395902c142a68b085350e3f09f7cb527d120bccd21d61dc6c234f7a86551dad53344c8c4c7981e8de0e51f8021665652db78b39128eacb2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b00915f57ff0cecfbf7517b36ee7d09d21b7eb8591f43a5029f99cfe093b64f5f2c3ca747fac3e8de974bff8cbaacf6d770bee50791b6cfa021cebd0088c565436444e2e59b65fc7700fb49c76de6c38c92b59161f1945c9ecc36b80dbd9a1e804399ca6e75b988edb1f307cfa66e9edc50ad37c9e0cf0f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1978cdbb8bff5a23ec9d1d87ddab3caa3d24950c0280c38185251d8b004fb99a636381f0c81deec28e446d9fec4732248c1b27d469cf4b9ddd6dc16133046bef18b8c4a40ff287417e024fd0cbcd6a97e3e0e348797a60faa4379cb8403e1db52c81cbe042ef2bb29cac538586c7ad4280ef34047316b5d6e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10a361a85d1e5c376f366a5234a800162a53918c91ca534d3ac840d6d6f44f08ea25777a289458c58d19170d5d49233f1e803357c288ebf4f44be12e90f39b34a6ad27157083491d244c4b7250aa0037fad09d1f29922e4d181211122394e0b5050942a7996b17e82c5ef7cf2b7971c761a3463fef20d994;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc3d2cdf84a42d3dbdd585bd01d8babbf6250bfab4449310561bdef9bd9573a9fcf1a91d77c5cfd3b4ad756d68342f949d24c95395df03acf9e92c627cb5ce87069163da8be5b9f75a779a27d3979b1d63574e9e64d9049ab5daae1561d65cc961a25d1f612b35572a33aed3997e69979c0686e6e0fca90e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2276f35c39b8376db43c5c9433933c6ff91765b0a814398bb66d02f6b69d2a12bef897e17025cab681da467aa2430b7168c6510da4a4e14ea4a769790bd63b42da9e99aede5e2cf62261301ba9e55262af54bef22d871d4822a01dead84dc6e58ec6a137d549f8c9c29071cb6a9662a76b81e617bf8bdb17;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h199dc0ec23d0bfc7573f21ade93a30776dad4dcc3beb7b7b134df7035683475c0d7318d61d450de071b9c42d8f2fdb782b721f421242179dee64290d28276be467e0bb008658e6174c0913419859aa947dc4adcf73d2fcca942bd0c580ec83f1c55830896cb76924da4c42406d55fba21a8d7d7364de9a43;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbbedb92d9e82f9e9fa7126d7038b6d25d563c58849c1dc89ac7bde9ebdbd91d1317a58dba86e9d0e6a1b597056ac7cba242ea7644c5b0ad6a71067144d5080d01c6f5c9b01ac3102c88fb0d6e4e2e5367bd33200f4601fa0157cf39f1d00121f520bf08dd2f210d5542f2aa71ee20ba775cb8577250f7ce1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc76142ee84d91829a6eb1592b63a94cf6c65b06ebfeccb01456d1c0b72b945cbd88ca34f1dc994275223dfab39ee528779d25f44e46cf7408ac386a35700729e79cbd3aaf6e020f496570f2f740c9d83fb5594343d4e92d056bf5aac0bad0d94319041847b583208f939422a02af261005e5f6e6cf86a8b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h154788c541283fe0578c52a0f78b98041ac0627f4785e3e2a561b481b0ecfbd3eb5fa64b655376aefb0f1ed027d7a1fca05464dc2f730578b5fd851cf9e5f24dcefe028cde08c0cf6dfc69bacf897acb5915ee4a337bed9b67dd4067b9b84cd75fc46dc9738de8afc5bc0a30b88ba29d509eb24e0bd89f104;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hce7b6a1ecfa80590ebd1e2b6843d2c8b9065ee80f0fd3bc66186c30987c6303b0fecb13895528b743d444b50a57172d05d15aaa29a4fa5542bdfdbdf98b532ab364e3b341f2fb08a8864dc67e530b424f280df5bda0448de90b27b5e293ab27d48065ba8abdb944a1543e32f6b09e3cfddf894a810d96cec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c78b3fe06fe6fcf26ff9f2a72dd23ed713e1b1ced7c61e29c6f0d90c5d8a6029adcad753a8b27a9061c5a4f6db221e7a1dd166c943816166ad202d5caae03bf0a8bd94c586c9c28d0ecac99e2b005b1dca91a287a4184e1b33141cb6416fdb446e759e44d389f25748bd457ac68d9b16e017b202300118e5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc8364f5b134b9d5f65706a9d54781bf7b8e945f3ecf0c8fe6b357e3bab93dad4eb8026a68153ebee265c3416c7a1a1d55e1fe47c338edae08e899f61aed07e50f4464160a4094a204f0e0428699af504a55a90d695a2f88ecaf85cfd58500eed01dce2e7fa76919610fc581ca169d741d473edeb75e7f59;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h647c8054e3e3badb27baf6671b9f7d49c5390217e0884b998596085b7b4889cfb670492ae2860e2856fa0f4bea9f2ff1b81c2dc978dee07cc54c8744a539a08b6e1870340d4f9cbc649aa37840f0b856e9ba885310cf90b1b84d4d021dda5522131f1d7c5bd7460bd1a6664c79c0f0c8448a9f7b15cd45c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb156065f56aaf83a99ba65cd37c2405f7967b270288172e4467283d36302b5cd91727f460d933ffffe46dadb5b7db50c4c0b0bef1f680c5068845837fc5856dfb19a765c1c3c49e7808a8d35a531513653ca41a2df2f11e8773189b08086d26d3c1c23e547f8d2ce6f55f9ffd2718a23165a3f89e07ca26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f28780c788e4835091966fda3b31b8360e57e7f675e70897cc7461c692bdff3fa7289085e60f8a7554a451fad921d6fd56f3b42f0deaa3eba532b93c77d7b8328933eec4dffccdd42fc239552b905bbd840f8498411d71a27d6cb8270b9a8119febcb47e73dee4637c1e51a43ffa36bdf8130772879230f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5fad81d5ea8a5173d5779f3022141bc59137b0472b61a8659d6be4d7ec274b37eb8a19ae21ce79f05cefe39c7f0683ff9ae824f7e90cad65a0b290d16525010220a9101c46f366ba4d44bfe888b328f31a6a2a6a225f684e9cd287e107f5701280b8d5c516c6b26797525838c4ee7ade65edb78bde0042e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f37cea310ded00103c951556583cc32b21c0cbd52731b2e4f5d0445b69321dac8fd02d09a50fd573a7e866c257f681e6503ddb68e6f6e3d1f0f73a5bafdcaa50700fda8aa11b04dce6cf8c024decbe19a1c2ce4512a8b214624d6f472cb524c04d5326e4d02f121cea5dc5aaf8abcfbe2d34f44f131df475;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37e10445b7cbba429f14a6bfcdb5d8d850eff5b24c92c70d207346ce87f55edb9ed4603498de14131b75acf18acdf3e29c32c464119a33a20b608aac93a7edb36a3d19509b64bf1d99b24fa630496a4365f257ebb165807c20dc2eb225ad91a07b15244b0756527b8ac714a5ce4a77a1d595e147de518542;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f7790891cfaf301c3d01d4e1b751e4078d61016e166f5ce771bb43be69266248f2c758c533fc0be5ddced64262f72f9ca3b286ba7eb1f65031f1283d4b4d7af69681e42203f0eae31f9602a9c5911178528abd9ffff7c1a6c25afe4bf818215cdc562a6a9c8d96f89eedb2a3b5e706c866daa49eea5db94b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfc643b192ff25207767aab23d40b2b3efc25d4703123824d549b5557edb21442fcc623aed94a9e194af1ab733e44bc25c5bfe14f3676d871b4902a801f0df464fb60900a0a98f60dbf02e60434c73b3f711858fc4088e0e209d9323977c5331088d122dcf09749a2af68bbae021f6c19e4db8be6e6f6c675;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h47e8b81b2651487f79265b6435282bd03adfdd28d4c40b62927a68c9ab6060069ab0c3a3ed384d37e60accee9d55b0c612cc1b710c54f020881d92f633aeb98e0e15a55c503c312f0660b5b784272e89596d4c0ac671360a5c1b9d81c8608d87eb6aa3597324fa3463567d3521ee4537b3d410248a1c1c03;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a0ad70b2faa789b80ffba0d4bca2196be45bfbfbf6c2160d67c57cd62552c331c94bb19f5ea0715205dd891d858c82b98b27caa2419def638e0ac92976db257c7e5e662498320d2bdfbbf94e230cbec43797dcf1a38129c1b3d9392fbc2724c307a19ff969aab7a2753a48e300220f9ce4834caa4c89461;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0bcb86a67651eb902174110a594e4b465d7c52c72ddd9a78c80706d3501056c4e00dccf6d74eaa8ecd1af2af5d271fb101be33bdb93db253c478542d91d70c06243e10f999d8a0e2261c3f457f1aaa82c288d5d1985db4ba0f93bbe7d3a1ac67827e952edd56661ae01bcb8d1322c989e3ddea6e6a6c09f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b3f94d1e7f74e394efde81642053f4b128ed0d8ef7f9c1c098dbd974144bddb654a58f65326f3463e91c4c4ca92917b2af7e4e9120f7424d74434b4a98bd95eb99f0ed642801a5712dd85d0750c2ae17fd84521dd6d7971c68289201a43a2e14ada97d64bf10edda93684f6513488d2b191b80ae400c79d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12670fbb54d05bad16b3207c6f263d91e4bcfef839f219c34463ed2876324b61dae484631e449ea3917167c527abd542bdc4615073edb0cb0e30bff5b53a82bbc718d88efd91f44cb02dbad9427fad9a3fe93d80b76df16d9af08d8fe84badeecd476d47260fbbcefb50dab1eaf9b2d5fc5c21dd00966c8ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4303db1702393930bdd76c0f9d3e0dd33ecf490dabd606a077807ab65a4d06175211749a28b9a06debeb7a927731765f1390f0a36bb612d56b2a70c8382f9d369544ca60ad2069058d5abf8a5cc4fb0ac341ee21f4f18f0b6e12a341823cb7a99b5f02b0248c0f4cd572b2218585b59abf516dc3108f60a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc4729257895cc561caeb1e74b9793f4e95dbd0abc9b323a503afab74b0464326437b5b3aecaa931f5e5f58cb124a5a8c8acb6459155a5ada78cad0978da5a12e1c4e3323c58e88c8cf281526eb1ff0994cc241da14d75394183b5304bea319d86d38f4d6d9c0e2003a039c261a633a8873e1417676ed9ff5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d2bec257153dca85fd96b26e47f2fb65ce042483f1d35a8f5abe71405073c27fe3553d825eff87db60f65abddd5d80484158a69d1bc0a67bb2469cee94d7a8b933a82fb185dd1fa4725f50a5045f0f15410eb89e66704fbcdc8ebf392c92cd0f4fc8754f28b7aa2937bf39356ea07a683bba93df897b9f79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195a72c7e201897df3a90b9fdf47c3b7acaba5a76307aea40b23cc45e9a3b2eb1fbab2225c0b321cf930931b387da6e9df1be227abab6878a21badf446b6e84a3a6e395f0665eefdc9ac18a9634b4eb65651dc0f4db05e449b7a5842284adf06342cf0da57ffea10267c5ac2384d86230eead31c771b655d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef8c0d8b30733c6231965f114008c75c626706fd32018e3a3f3cf2c57e6685b4113398a97d463189a454fa579d9ab9f5810f7290e7656017c5b63964c563ee2d5c1ea135bd68d16930340e940ac9a08008b0cca678ac20f4fa9880ff50cadd2fb8b8b1f50cfc792ac5c7e1d4271e8b9c70b6a489276feeaf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13fd4d25eec1db8584a97cceba927ea1f79d5677076f2af7f4c42c1224afa1396560cd5649b7ba1dc2bdcf7c52ff9b0f64650c491a8923a512898432a3cc9926cd2bbe6fa44546732ee8d014635e444d249371632d616f22e3fec7bae9fe53c24265bb0f49f286ad6096d9bf9e51c72fa437a350191cb7aa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb32ff2a807e6947c053dc0ed3b93e3445c62a6a6a463748d61ed98b53af3b1796899deb660485a0c6e8cebeca9c8d5b9f4af7748da8cc01fabfd873a63437be5b90b9390c1a3964e19f6711245b94f5f6ae849606275b783b5f028869920959a436f3c93cf6fd42443b41cf541e73c4d61f8c4a054522df5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h143a96ad4f46573111b3664bf0fcbcde6901c6a3bd48fea56b89189389a2881014377277086f917c08696dfd8bfce7219621a43f77ba7721dccf892182ba97ec2f5ff993b111df09d24c890ac229a8fab5f8786a998be9d4a1367979545da102e08d442fffe9ff13f6f82ee7bad6a6ed5aec56fac3aacada5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdcb2dbd5ee1a203e70a53a6a94ef4b6444a6aac37d9cef8df6302c26c8b40ed8691dd9a7736ab7f316f9396bb2f29fc8ceb14fd775f6dccb1c0a2fc79ede0f6483af525e68d553b23ed50691d661232cc3880f110160261abcfc4cd9e4a484fccb12adce2e08819a1c0feadc0165092627378566d991c4be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6b7c79d3289157578928c8d78f2bf4f24870ddb3091d1f63ac4f1794dc403d746283eb8d8ec0bc433ddb49e6f264340b81fcbae70b688f07d9de573077e064169bec778d157f937ca754293c3ae302c700bca39d370ed91f267399a2a6b3d4c5294e4519ae11b9986696c3fd9b869b05e72ef01390037fca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104ece45ceac723be561a61b9e16f3688b4a11795722c079108cc601246ff37ee7f3c12ea81856538cee12614e58cbc9ddaaac9e11a896faadf3a3191451dc6699991da248d76a63f94703c1eb7acd3eeb2e537610f8564d2e7f458aff2e136dbbd349781ad10642a8a3f64bde63e0512a0ebc6ab34057959;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8207197d60f532b4fe28153f7d6b1dcf9ae747ba42d2f70f9995d9b35230ee0b3248e4823e52034813db1bc2d829636a6b44c04842b4fade0174994eb9cf0960dca2c7fdde4a310496caa8c7264f0524b9e09f971fd7d63850edb58dcc3a6f82934d3c7a8df1e98ba9f6b303d8419e50c67c7e2bf470e25f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h155181d5e07cf97998fc2f30007d0bf11a2b773dc1cdb79e0a32ac1977698ff231fec438a747dd324058fe73763e75286eeb79e2ef7be4f00b909d0a8e1c001700528069a184477f35dc61b637f642afb72479b0c0d28bb0e006eef03e23c436295e332d789bb78ad6bbbad65ae7b0dbf5f7d0a4fbc5907a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d592709ff26ae31c0efa293885b5ea817ed6a86508f78a9718503a620cc53828bb19c9b75e0159546383826a2be6c30113a5483999b4de890841fe0fea3fad60d20d01b6c93d79c7a5f549483a571cf6da1543856ee5600cd5e165c3f172522a47de473d4d24eb5d916d60789ba1623ea71f78c793196d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h517fd5e5b6bb59b0cbd494f2f3acbaf2afdd76c336b8ae7ebdbef34dca232dbce773e8cbd7140ad5088f7c4f84235b164a689668679d4792189b15414bbe4ba33e220fcc4a44581533c32cf37f541e3fa44ebcebd0e5acf792e32acdcaa20897c5a9c1ee6c5b30f86fa33ac6b7f459609fe138dea8139b66;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdf9526d7263bc5c18e6fee6ffae5541119d8cc9f78cb97f36d62afcc67e1bcdb997d971b24452ade4b100fe48f5d5396b5def54fb8edeca0c0cae1f276820a03d271de404da0a40ead53c565a9a58066e2e632e6a32da6f7ec3ad61257811255fbac1b143293d973f3584630fde6c1c45828d29a3f002a97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h124bfe3515bf1c3e711449a10193b2aa4562d3ec679358136a3d581b553ac8826287686dccc5522ece011b8f5f6e5b6e2de8395de024a998e3baf205a6639e2c71a15e00dc18aea3940b2b784f0c556996eed34014e3900ba7aa47178449f75e77f63403b73b3da518a2262e574b765d37bf46cafa2888b8f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf05a8025a5684af7b29262a6cad6f817efe4d76d8ffd7bc45ef446cf841e5a3d5979e18dc137f533bc0ae628586523934762fbac330da60fe9e7eec206c40b611d3b8e28b53f289ec721db55b33d6c8c80b9d1426ebe5f3c22402a017746cabd82b0157220a09892c1cc2af8fb5873ee5a7bb6dfe0c088fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd3995f2d93e68192dccc1902229559275e1d08a44fd4303fa57c77047e121d6a880319150d2023e4f550a24ac0be45d593e6b6d8dbd84a8a6e3ef9615861dcb0c69174a7c7309b1f7bd7358454b24d317a966cb319468bf19b48897fdfbaa7090a4c1e4097a7185217c9589a71917db62695671774e48e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1990c62d8a3520ecc944f8b8cd3a19e5804bccffc1ed58dd554b4808c744d47fc99a9c2307fc11206c9134bec28683512f108bb5754ce635d649230745ba91cce7bfdfdb597e43553f6e914517801e6667d2a8e16561c69d3f0775b2c18ac644628caaedd143b3ceff2d51b58ef416224c6d13158767b7ea3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h422a0a5650a08ebe0b77d5398b3e64042d70662d79e8aa557ed10ad81cede81e4c7aec8c0c978877d60fbf8f257589bd0376979a233277b164b7917f26a61cb0f98a73ab8f88769255ce6952d8b6e7f8953bbe666e6dea50b8215b5bee6a0cb95bacef52a01f49217d96262f5121b8fd74137d5cef969de9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h141da753dddde46743945ddc4972e628bde7938c380c181855b018bd915dbe470a7a13c069c438aab9f32d3d9124fee786c4d9dec21eddfbba8eb31d42df949397c6e1099352c813778afc9f144810bf6d63f81b702b5a8c8c8ff3657bc9465b6b2da3fec8e94d1744701faaf663ef92c2449183c184895c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h593a7587e70cd9f898f45ffc45e226a5b872b6d0b890a3f3b0f131e1b7095dd4e6da9abe6d4e60201514aa96fdcfd9061c051f0abb884b20bb51cd7c1bbe4b964993347b54079602387b3ff82c44cd6331e79ec0a601d2ad728147382d34c573a8727e8352b278f78e9cbc03b2313ad8581608c12ddcfd7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h180f50d27ccc8a527939249ed105f67c2edf585c124fb02ff0aabe0103e761ce8a967b7bf32faa3b31656bdcff70530f738639885ff3111e5f58b632ad4310832841fd2caf539aac49d4e90e52f74541478fba12a5bf2ef5fde4207ab8120b64683cd953106fd71b50389ab68eb067aca3ad012395f845455;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf00aec457044afc2b9dd86fa4ac102a49f3cfa7eb4f50e2de32d866679188050dcd3fdc96363111a30b17efdc62563251971f7385ba236a9df281871190e4f3fe1cf5475908ee0581cc0f851147bf021378ae0c36b34b6d2bc547aea8217141d2727c98b44da147476a625d49ed83d276b59cde41329e1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d73027af5c23fe38fe9888c5e40f6f2b11b4581030f1b9aff0a18287c03403b46e84478c2e03a758265bbae9bef9387b1b7fa1196a1ed9b125109e6f7ecbf3d134bd36b50a62c695b0fcc9dc82f72e1ca93450ac791a39ee192a7791d4218faee92fd1bd840c1ad46235da26cec60eb1a13d10e8e15bdf2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b680618e46fb22e0044c318c580be39f4cdc72fb4466a4f5c795bece55157825f0c5a30897a15ad326657eb834aeaa5ad89ff781cc9d946a4fe4a55d1e561347fc0f1d25c63f6a5cc7b091a3e178c706abb973d7c4c658d98b16bfd8bcdd2e26ad162a4f58d1ed2b33ca59033164213ad23bef54e1780cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0ac1425e27b8bfb1859a5bd0fc1ec76cc966e05ffddb0bfbd2f94c287bb24421b9f065f8186cc135f31a63dc621556b75e3f0a7e3a5c0ebd0ddb6b91304cc3198b88cdb7c00dd1290a13298863284ccd7abe41486f19182363269be0ebbc0ba2d67b5d029bb0f3a7c75ca860c677ecb9f019a9aa076cc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb03730df71a648f1d623b348fe266f11d2f51dcd60d474332d34714cb0d7f95ced69c1b85eaec04141a1f67ce31ffbc0dd4627a67d9cf1ff4580c62f9f5fcbb9887386399dab070988a8e0dd2e0eefec3db0bb29836c6111ce75999b1a2563ba8a514645de26653cfe96e2daa68a3986c3b1aa380fb0b74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h163c95631a426fd0163d7b0cd4f34758b7cf016ee8e786eeafeda6ce5210d8bf1559ead5f5b74780fe93c9a2653fceaf07100da235237a85ba5729a302ce1c9fd58c623a261bc47244aa7cbb2fd13fda0c40a56a8a11aa7208a91f5abc559063a8293771c33f5b2d588af36fe555923129b94d843fa5f50c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab0039ead693a1cf84b1022b18ebef37bd17345b4643aac1b8e7b9bae87c678fd6b5c2d3714c84ee7aa5add5a0dff4f70f147e84d6c08ac1c982d8cff8ee891f0ded3a475ae8958f438f3f1400fec874534544c1bdd120d6e5da78689123fe459506c1b5e8405ae8438bb6cc3aed3494de904a17929f3d46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9553c0b6b4ecc2b13ac43dd9f58f0c153506e910f8669b40951c06bbc5b21dd25f5b9c7398351ba30f5350db8db98137eb38918719eac7fcc259b943807a3633330453717a8cb16c5b425fb5055ad1210781b48cd436f6f5aba7e1348552159c5b8188db183716ee8257f69c982eb6b3cc0fde5912ac27e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9cf86bcf049d1caaa03fa5b1ba6c242426a8ff1631cebecdcf80c25f67c9e78f99c95f465e010571145d64873874a674f2d46242f866628e9a32d304ed3d94541cb5e08908cab4d79ddcdd2ad2b6c54e2f3b28b634919e22f3fa9060c04f1b75d1e4c504174f2251636dad4893d319e31763321cfde01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15491c49f9a03a4d8c2ba9b4f916bdf7572848ef792e3d39c3a04fa460eb1f23f1dcdacd8993f538e873adb5df5a2610b9d4b31752cc2dd309c2d58dafabc692b1bb34bb9fe316c42e3a979f7771e126ac18cb14620126094edb0f022d59a61602f10a1193127fd88f413f949626b9dce33ca9c0f8f92bdf8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h54029069c8ab77fd7a06452350d34a696a8e7664d1c325a1c459e280fddfce98fe2e7b9e4093250186a47888a6f4d6469c58d8655d88176ab81f05cc6ab6a4d7d2a7916f8112dc7a9097a6b508ec709d52ce05c66bedc722a26ec22189775efaf12049269b34f4c2908090804532f25a516648652752bf41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb399b4ee22459a4ba97c555a867a79d2f50505937b3e0836f55af22bc46b221cf9564007c59d48b6616024234d4a5d5f317931c24d92a93dccac80e13c1768e0e2d499856fbc72adc80f7cb7018492f6a4e0836317dd4c633d8aa815021214d47a30aade3ccbc572a301e2f7d5fb6e9b4b51a2a91e29ea2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1614ba00578c0ecd8c9f27872b896e0bcbf6b76690c9bbfbcb7b15b867bae78556f1065889db5798757efb2a314acfd480c0318ad2984148f0d8b367571999070d2188c68f6057477656cfca82fdcc7f25f06ddcd3b935852a202e94afd47d644f4a2d09f77a82f52422434d5bbdc82ff295f65532ca2f4fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1346f76994d6d4980707b98d708215f6925525a8f334037ff13e4779f0b2b43c9ca9d3bb91493f93a6b0ae05cf26a34bcd298fb777667ea7e78bc3424cf8169a25a17af1ef4485018169792e36be4f3624011f9436d5558d4bba7b05f5f55754f54f1edbe5487caeafb4da348107d8491f43cae5713d6874b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79ae49549dc628829312542bad02014750e2d6a23dd11e1c085796398a858f47818d26ce93ca02e089c06d3a743e83d23d5e5847a2c1b470ccf710cfb555b7793f75f2c31cd591752db4722e1c8be7794c1251506193073ea9a763c2562a94bfac6914d9d42ffe9c5cb107048962b5f99341629eba8500b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d14d1b9c36c0b1afd98b65366fd83ad26e4cd5a99efd8973f4cb297b69b377521fff8b1a7be5922147a16f87d5e5664a474ad3c6f856d7c7331d4e7df793bc164785846dbb61ce5c8b5cd9fd539ea73ff23cdcb12c00c7f5d789aeab9b39717ce1652eac5fe380dc0fe561980b5b16011a6988ba7444968;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c762f22e5c9371f735e9eb9841938efef7de3a7d25bfd306eca537146c72d44479a94e57ae86bcd04b78246c71dded5791a7809b9c885100f6f1cbe2f14e9dc9cfeb761f3f47b7f97bfa4dade2e37e15d12fd5788d950085859336aee69eeaba5d04a363ecdd126b14ce87dc6aa19ef9718314083d7a8ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcda67ff364b7331ff440b8d116dd41a2e573e8d1d1c9fcc79810bca7d566297a47a04d542f20025376e1adfba98247562ab00793c122b7ef7030b7dc460c10b99f504d90ac33d2da13744b38ed7a28684413ac0a07036cff13827ff97f9dc8360edd2ba622a69b35fa712afbf17ebc08573e3549d42e90e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hddd0af667551df0c138ed05987b49e2246045776d3a067a29379a35441c2191d685de106b50172232f4fb20e7374a0bf61c58e170f62d530927fa2c014801cf9c6945a004e54ae9e6a76b96fa176a7d116154427de70c38a8d8fedad03b194c85dabdf3d2fc9ff84784a5bb19e3e05e8dbbf71a72b66eca3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12ff0c4b532f8c7fa5cff3f6d183e8de3b7b0a3c015f9078e873c81d3c99c55fa9002be469af18ac61a816a81d308db19c6dbd87e68513df8914ab8da6b45599af2910f7035d0fec2c5fb4c2feaa60af77beedd747932ad4029dc616c3f58c5ee14bef673913a8bf482cb218d68af4a184858f95cc84f821c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haff379fd516ac2e3de5627992718503c351ed7ca082ae2ef186dbedeb5f936d0cd4c83a41f9afbe83e73ae05767a51c3a217aa1c215f0705a0c1db09cda4c4bf0088ebbc2d251ee2a93da9f764dc1348feee49569c85f5723076f26ce9d7c8fb35ca4e0a17adad0b0fe9a80871b5e5883c1a5a46fa7b8120;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65082313aa35a46062cffc9870e841f4f15fbc353e5564c09d691796cd6cc9309fcd4cb89b45f2df0497a62a2ce6ddedb9ce92c892afed0b8579948617c60c5f3cb5e0956e1245ecb8d3e11d190d97151d197cb44df1184d75b5416f9002e4f88c72b694c343123be7007ceb1fd124377750f084906d6366;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193a322eec3c1bddf7623ea7a8fa207faf9955e231900fc155ce8ea8b89ff894c0f4808c625470bb849aa99935184535c90b649f604c2b31619b8f7045dd37f98912ba226f5d10c6cf68d4eb75670755d153c3938d14c4f5c47b8c845044c3ca91f2a941b5627f2a70bca6c72e642f23d97f92d3e748408f8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3939235c6c2760f5db75fbbfa6dac0d58889fa291db737bdab82bbcce9298dd6d056b83146bd3a58f9b97134a3e94462bd90905d102b33c80c8a56bb59818ff086f3329fdc4ea21f55de2d4c74363048f11fffa127595078a578aa149664cee4ddb4d7e563e4ed43a9671b0905ca6ea148c21ebb3b1df1b;
        #1
        $finish();
    end
endmodule
