module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [15:0] src17;
    reg [14:0] src18;
    reg [13:0] src19;
    reg [12:0] src20;
    reg [11:0] src21;
    reg [10:0] src22;
    reg [9:0] src23;
    reg [8:0] src24;
    reg [7:0] src25;
    reg [6:0] src26;
    reg [5:0] src27;
    reg [4:0] src28;
    reg [3:0] src29;
    reg [2:0] src30;
    reg [1:0] src31;
    reg [0:0] src32;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [33:0] srcsum;
    wire [33:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3])<<29) + ((src30[0] + src30[1] + src30[2])<<30) + ((src31[0] + src31[1])<<31) + ((src32[0])<<32);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf7cdba49a782493e8419c4f57142939de694b640c3891ab5a30c41686e3b64488e797700;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13563c98dc11587e643a4b0bb83563a7e0b8e463ccf9b51b5161329710f0c2963d11a636c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6e3057572775412f33e51b76b0791364bab6472cc6f5e2f9cab9541d4680bf470c04970;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfdeb407aafea22ebca7bb7ee0ec9feba4e3e7a2961b7cfbcb2b5aa39b35b366e7dd1cdf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf3a658fe447b613e88ce76b66085b8aae6f0f532e7f1dac56d4780cb430bfb48083a800;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85319cfedac379815920dd635b63a27f8a90e8b0ab9b63955492cdc9d1ee764be922f7db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5cc791c66555bf74ea2dfe56791378344754f8e519c13c7ebab88b45f55ab018e6ae417;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60881e12ed2309b362d12ea23bf5590a9fb0f0715b35abb1c273b304240ef50a7fde057b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd430487402b77b1c28d192ba38f1631f7d49d9cd5264d096f219d9473686cfa225618ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b2bad8a2f128415beaa3104c26e0f2934b1d57bf78b2a7a076a89fc5e86d43abe33663a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4ac3fad7e5ef94febaa431a2d91e7de25263592bff41d4774ef47236975a49e9408eace0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h708daef4e868dfadc84596785827a376af99a1e0ffe8eda6e75b8234aa55b191cc536149;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91bf4bfddc9cd29632da1a21176b2749d1ac638b48dd690ea9b2eb5c1cd9849215aad50a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5b84bfac66ce1985afcd3bb3ee9f62f2415f9c1f12913b4fec43ecdb552b4bbbad9b665;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85a7720c4b899300365b186d82e653d54bcbab7898fe370b90cc7f5e3f80cfa07db4f2df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdf52827f6df35924ee0e87ff901b20c77f0a37d91506535b2dc9822767f7cc051a5c45bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1d3e59e3bcdd90a4d32b041e934ed4a08cffb71ee10c9e0acb150576bfdca94be7a8872;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h102a37242ba7a9ef81198e0c4575c4d51274d860045fd785cd9915634547e4b4e3b9bee30;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca4b0013ae46a18ee1cf3078522e5a00743603432fed6026a1be20c4d272a0436d29e14e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19453ba26511623e22fd316a1f95bb978964d2a71a31e55ded3ce595731f0d5e60bd7457e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h95cc159047bc420b044e8949225f7337119632bf600f40b8b333fabf2782a9bf5c84f193;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c82ccbee7e6b630fe4b4e6ba8887d74b8f2d306012b8ade2ac0f2323edc75f6dfcc274c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e12b8ee2299cf8f2b168eb3d5a56eb56c02eca879dd7ccdff868d4814e55bafaec8e634;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb60d62f9d0d84d932527686995ff2269fff550b8e9165e5d20df46673ee5c9066c003f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa09be873a16071de52763247f70592bf31cc2fb4f0df37cecf51f9d77d2917c3079e449;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha11641395b916c8084b3817385d6df2a2f332f68a0ceb9f2e18852120571398468c5e4af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ee290a1c8e19bc03b40f2c791257037e6acd53fbd8fce869c052ed8f216843148cb7f2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haec5d9f6b180f99f06d54bc66ed1750098871aae7d0f4bcd260bafe3c883daabf5384f1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ff470254fc9ad9efe99dab5ffe2a4320c0cd3efc3c57f0815bb7bfaa117a163c3df838b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19fe53b06b80a3df7e29b6a36ee768c44336ad37ec61399e6d203ca44d02d2000e2445f47;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36ad2f526399f2d5e30c2ae376a1d4a67a8f2beab6fa2f12c8a0645656ec6ef965a5bff7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1174ff9598b392f23fb87d24be5b257687a854e6d3604ce736e422570ea24e59691f46c34;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he523fc70a835fb800b32e83912bfbc38661d20b5eab32b7128e6b54c6823151a6e748629;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d203d00584e1bffe85bfb891a6fe0cd20bd29b22527cca9cbf5fcaf852ce7240f816794;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f3a88a136f5a369f2f57ca3ed63803e043e8e93eff82ad7ae238f127f091d994f664a1e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f78d11df4a384626fd3a6a5431f562eddc0059b41b13ed8b40d1ed264c248a8e0eb48bb0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcfc56cdd4401f052113b2a96d5a6623935b56368a6c91b4f0a16cf98669f332181dac835;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c661533c99221a5e6efcc4954362398ae386d5955db9f81d3e64a4ef703d69c49c475cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187ab97bf1f8934439976c6551f2242c4705cb2edbaeda90f57203edeae6c2761d6ff6c39;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1364ea8819d8c16187835e950d892d48f32ec6c7f8969fb75d0c062d3a958c3eeec4f98b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he41edcafa017dfc69b585f103c4e522286c0cd7180495423d5f9d8c5614996844b7f58c0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4146be0dc8590334e9cb92f2dc490065ae396f734aa1ff69b9d5af5d020969f3c3454fc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2297576d31dbf726afad7961a11a5dd8789935b4b3459abe03b081eb0a34abe3ee2622f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd815812a9d3d0fcbb2289052bd901023e9135628c58bfb2dcb273e844cc3a3dcacd63061;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b3ba6be5e242cc4153ef903aff20158c60ad9363071d549ecbb264153cf6c43c5a16015;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h35d8a6f703b646ab40922cde2682603a3f4a5bfa68d9f657c0f35a9b4cd45886741247a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe870ffd967b479a1390c0bd923d373ad0a7d7f6e54563525781554e31faaea6e19f424f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b25cf957614b15db1661bf7bdd89debbe9d2a83f4967867054767627801d5609c7674d14;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5deffbfdf0f4265fb1df2c4f1f74e8a9ee8a22500422aa87c4bada673b7298a95f3da2fc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b0324b9778526f2e0b6f002b973b71b162879c605111f349b3df3d606b1ee65ac180c049;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h868511164f6778e54bf61ff0b55aac5d2d686a658cf1e62797f416140705e8bba74a30db;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1201c2fe91c627c5d9ed4293a77c620454f1ce647b9a4a4fd7280d6ff7a093ea7bfc8503b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c77aa9fdc38ca8032eaae3c02d1ba74708f97c808a774f5d997b908bbc5455ca513a202;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a587831250cf38aa7e3a5b8d93167b9b93fa4d20f6a30f39102452c6b2eab31a77d5bfe0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4ba63192d63f1e3a82fa7cf59cae4aa05572554070c450214ad43d202017c3f00c1113a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13d7466e68105c927cbfe43fb871597634ef4ce4e7332d1b38411213bf91d31027c83c0e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170f1689c7fc5e1a36873615b868a31d967808ca9c4c97ada184ae853dfc6a97288348748;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d94fabafd949edc8570a7a0a47c58bfdd397e5ec3454ddee49b9392ffc40b5746d082145;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8c71360dad66a0bcc352be0fdd5d6a02c87ebaccd0a4fc2b833680c249905703866fd7ff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b4758834296aded3bdaed019602608efd222229762d404f9a567661857cee0e5aa15f94c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4658871454c8db734d55c4dccdb6da1ad23576d5e61595f7ffaebda6994f14764fcb41c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdcb63056e085c806391c74827342219bf7438af23acaa713160d95d55422dcd61c6c11f2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c76282b1eee6ba48a0957d3bcb3763e9f77621c69d77062b052b63d8088aea04f55b2970;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h56d81f876ab64f8b917e02a07638d49e38aa277644fbebf451dcd532575a2fddfbb58218;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13986dfc4b7b4133e8d8b17e4f8dcdd036b13d787e8942922f06f834da84c805c6a71182;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cea9ea0b14fabd71c87307be856132d3f6fe187b7687de692bba1c8b585fdac0370fc8b2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc19ab72eb7000eccf1379e58f359d0d63bf7eab60e0c23dc28a868999a401e06e00fe0c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111460746421097cc7b5f7eadcad26362dd1862f81a9f5e04e229940b47b5323aa467567e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19be52cc162934c8fb3c1e9e45a42d6eb1cc44763c98a483d1f4689c487a6e37e5378f436;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8094a8e1e97983702c5f33fd7c1f2cf0e0c5dab1f50ee6bc269c6be27cbc570c6ab20a0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71c6ae3bbcbbed605a443966ea4b95f5aae884c70f85327655e599930f7830585cfe1b54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0993c602355e3b1b9957b8c5b0e6d288678b39d4257ea8ebf13369156f6ddeda4f8a214;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141cc00571e95258b3521d9094c4b467229b5f153b0424d2a76ea0f7f9c13aaa1add1d19a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0a74dead0661c5eb3fd6f0f8212439916b141651042f29a4128e925c28cc7c7e7fab2bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ec15fd8e338fe444170ed84eb623ed7891642c2ca713f28ec57c6744a45dd747c6963bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97f92ecf1c9dc3c8da3a67cafacde5403e7de4e6deb6725990eace5ed16cec08b878abef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175a93ad8d6918a1ceac4ecfbe575dc0dfb0bc28a52851dac701a1a7aa20442daed7af845;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbbffc0c744c9ce884475d20e0bcae22b7c41ee14a1e9be0bae10713799acdb155d360a8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12de159148511bd2d2966d0cfb6d95c4308a500e1f87ba49ac670defc6f38bb2409b4a4ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4ed3f603c0e8d79520198cb7dff7f2313e17ab27b096a8bdcee4c32003917c4036ef113a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h496ba8ac78c1e6ef3fa86e846fac045388d3b9402354f8d1d0ba9657934f5a12e744a5d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b8760ea38ac6bbd56c0d696a496a14edad70cf32ae747be235ec29b1fb590b35ee74a2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11bb39d4ef399b004aa883a09ec4108601b8869fd87aabbd00fc751e32efa4d82ea7c5500;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1220d7dd6e71494b5fa95892647bdf537fddfdc40a27ae210443c8440f59dd8692b3d5180;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f1ea355ee3b007356d3c96b28dada4f544dbbe1e8d94a3645c58947f10e1f2d91e6fb7a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c9a2359c17fd6aecca5d6e7bc24bdb43db6a45381bb58ac44671f76dc8084c1eaa59581;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d85e3b0204f8812d01bff650de607fe28baa0bf6aa688d55c8d28c5b752e443806a3c3a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h440bc8c35f873b423873fd0a01a26cf7e33db0adcd714d5a98c1acffec483992fb77e925;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66c5a9a34605be064eb1a1a1b1cbb4fca371f1b2637bd3d81d33ce93f9373a40606dc9a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d754b1a02e314855c9ef9a2ade8541b62a7c9fb2293c9dd19544bfd5919f9dc71f65b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ff96b12ac48d01c7d282bfe67aaf447988a1b4e3bdb88acf049898c364aa943c28e301f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1826cae97990912ccdd9d83a139264f7060fe71aada00854a81ead894606e84784f06ca2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h760770f5def46aade6f48445ac444f505b7a3c85819348dfdfe6ea751f97e9b6b50e9700;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab59ea5bd817eddeefe1f7149f21536a8621ae5ce9da40f4d576fa053cd4d56aec146c98;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h165971df93fc7ab3a30f1b063cedff9d1ef1aca165dc030e93deb500dd996c60ad42f8cb5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8ac8eb9c6b5975154fad015cc70e534278c4282701e965a12376d6e2b4b7127a403c23f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f4bdf3a8b1050dda80e6f72dd5d4eea79fd2e0051a3ecb8c71d1d0a64803a034f8fcd93;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h54c04423048df381fedb59cae0afbce7a4e0a7d3143efc4a201b32fc41ea67a124ce9f31;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbbec900c02750fefc5ed0867ddfbca0eca4676ae70d815f0093f11576d1e79e234eeae99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef7565f2624acb10236d43c8617dceb91f37f0f4ac0e304591b557098c7efa29a770c0dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b798f78b676c652ffa300712ea2cf2a2a7757d526578bdc8984c56acaea5a0bb20ae88b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e3ba76b6c924935c708652a579aedb910e68faf3d9381b09fc2bf7ea8b597959acd1c921;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hecc61846ca0211da5d38997d59dd243078bd8e4436a1a2ed6d68066418bfaa87324635cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1807b610889fd8b538ee6abe2203652d1728214584d67772c4c6dbf948396cfc62fd150f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1b8ba740d008185528c9c6382ee2a4f1c3fe6c77cdfcc45a71de76a9c7f4590bdf39cc6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab04ec7f0e40f9592141b6452e212eadce930275e1a70176836c949a3fb2a53250ca2a5b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1697e7bb81ebed9a5b8aabee45ce4ec8fea3cfe1e0dbfa33f8fa176a0810aad3e593d1afa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b79e2108735e7b935c1972383fc8fa8e66287d71fdd4234f5a0fb5b9a2dc57780cff7379;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6df3068b198346e65c82a3bafc397bab55d2f7fc15b12f8b109d88c36a793db223e0495e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h858e00185eaa6fe396e5418999ed25217464c26bf1e4d44bbed2b63bae1ba95c97ae2a99;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8840e188f46fa7cc2ccec514e6602e8f0b3a2be25216bf3f29b2a50a3ae502a56b4e9bed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51e4be9ee3fb0f547e284f91f0590314714487796a6a484ad1aeca8c69d3a59098eab674;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ec520fa4e71e370ccad257ade44be8db29605f4e964eb4cc13dc93af645dcff5446e226;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1857ed98b20a90fc68bb6309b573f9a0cd162dd7aa400bd8c42747d5a7d1aafe19d47b201;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15dfcebac20a68cf6a6026d1fe6e44fbf5718ece6de11edbbe4b2e3e5cb025ced42ee4a4c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h321560a52417985418b885322c6f56b9a55c2d81e8f862bd640e95301b4ec1326b773381;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d1bb5166909911c4103126b9bff6667172e5bca0cf9d12a174e32597854040834e106dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179755c3486abce57bdb7b72f1ea9c0832ae789164dbc32c5d84911df9a0a1e9384795b4b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1042563474e3a87b80dbe5878338a383240f2aaa4f4e4a75e4df684cbbadfab5820c28e59;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b0cfab593c3b832525ebc1dea5475f787899c10ad0dd8746867cf6e03683e1e478331dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf89b25699f6e59237f90a21dc152bd1d89d1c14ad28a95ce0bd19b6b069a739d0aadfb67;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bef9923a5f16732f323070a36aa703be294a536cb6b38e6a3d0afe5e5800e9aafddbb304;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a08d48806af09261229b5f9d1dacafb129053477f63517efcf3c226804f85c825063119;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ea5c583286e72aa31c5145e63b06d4c37e8154b00fd5bc31c027c393f71441b4955a429;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6e0c2c12fc0f05b4720fd41976825a388c446639b6581d7fe138506e7ac220f0b09d9bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59fd24b28ff8463741b456bcf1dda7189c5070af558bfe54134215a2e75243c4ba64e141;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb159d4fe86db5b1c3ab32adef74176c61f338a9f0058327878869ba63e67f707dfcc3b18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcd905088f5fe5ce19c468ce45521db1f0af47c05c382ca15fe637ce3f15d899d6a18a44f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9299e92c116e0128d21fcaccef8f334861008cdd4b2c8f6de53d90ee93265f2be9569fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195be802764cdd2d65497e0e32e43538186c5ce913677eb076e0d2c87d226cfc1e8e873e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77285f05320b97325587b94bd46f5609ed30b113436ebf7a90f47ac5baa1a351e6bd2906;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf316c15c95c39cdffb267de91a7f5f2edbd07e3bfff3c4c2b6cba96803f5e749f42e85b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1961aa52729a909e10f00c68a2d50c45be7de9728f078182ae1c60227051948b12002ebac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d01d0be2a03870be68c2f90e7d95eb333cb9364149c835675d58de20c965727d6c90149;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18eaa0cc2bab6ab56d8855b30334564cb32b53a7dfa359deb6ee54bc2e024ae508417a329;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37ff20a6f27bf2795e22db24dbfa6cb5fc53b0a0dae3693248d4a484aaf2f7c12ec1427b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h986419158bb15df77ac977833a52e4247cb3bfb58a20ba1979252daf4d75e5ed918b4ee3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf8a852742008e53a897ec47f84e97713b6662e7e58d13be050921905f1054004ab91fc1e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be102c0e2af6e9b89a972baef3d8095bd34753317bf81ed9d67a55ec705e68dd02381e5f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6727e79613e8c13f357e3c107a5128711d9294224c3a85427f371782afc6e6c960b72bd3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d53f4ef7222f39d502a153c31f705ef65a9196df091cfa8d08dcabe4b89bdd82aa87d33;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2cbb7e37dfd6d1e70607bffa1d7babd0bdd18b2fadbe8f91854435e51c66394d8d54495;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c9f8b97ddb4907bd3abfce40868112fb464c61a3e00b71a6127c9fad94f28e2fc088ccbd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9d7548d81ebae748040121c9f786573fa02138d65575a811454739cdd72e479ce914680;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6afd2f5ddc5cb3fc6bc30f78b83ce8ad776462611b9b191f25c4fbe51d2fd3d88011945;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6f7f14e511c3d643544b5ac7d8ba554d8a4c334d79424b18ea43decf89fd4e7860fd1d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8ad7a0633143a90b5c6ed4129e901070444bdba44e6bcf876632a3833c2965c4da8bd1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h417bdf01357024516dad6fe9960cefa0c3a1a6ae1b6da5d2b0baec93babcf191167c7bd2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1704dfa19ead15d71a8c265502c78f62d57755618801725694c8abd22098783da1a64ccf5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181223b647d9ae7c02be8be1b617b4e6c68e2c1abc8fe33cbecb6f1a56e2e1761f96b9cc8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h191c3985271735c2ec175554268412f688b02bbabf5d868ae700440ab61fba9f1eeeb4ee7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4895e18c03c07d10e10acaab52059af87de5aa6facca33afe51f171305a5098e061d02cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c59da56935cf0f50584f2d952b6f71a3955caca06eca7f988d0036c603e8befd6af7dc91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7333c58da6f30d834b6e651215e35f5991a3b1a04e943441fa199c1a225af1420abacc7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d04a662aba92cffb5df3ffedf7f06d1413d7244572508430761e2aa4ab40816f3f7aae5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf06c625afaecf7ee8a85e17f44b14205a74c5551ed4f6f5832766d2ed8fcb4616059974e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6cc977bec921603fd3107a3bea6bff2a9e2c2e9a7f45aebd02ab6af41604e4458eb53981;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha24b17a7f61bf1a2cec49896f8a9288ef38207421546d0f362dd27421bfadd38bd980ad6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13c785c4ebea723d0596dcb2c578607c3ad86a809b234c262bf3357f27f9888bdb87dcd8a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18dc3cffec3b3fa21c6d9525b1f2dc6659dac2720a7ebec3427a475dbddf5d5cb4b0f9b95;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e55a72480d5ee995f4c1d8b3f8084415eeb2342b6003fd0b1ac05c96e375a3127badf781;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h920d5866ae5292bae3839bd3ed17cf1c4085a14946b26e96b01d1728e6c4618636150855;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0a67570bc4b9be2b434139ab7c5869c93ec34edd47b1dfdef18d72670febe5217254e24;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ab7f66fe510ee4ddbd582702fda8cc0c6aaf078ce9de4de1037ea1fc8e33d0def0b021b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1810c740e2e53ffbdc968e827f2b4ad37cf8081aa769a122f6c3a3d1f4737102374fd74fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb16fbe6de3e8e952354369ed63edb48bf0568cc52fae8b8ee8d442c0a33f634c426ce017;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa46fe08aae9ed2d292290b05e708f85121fd5ca8c3f51cfbe2fb2aa27c1c612eae42c04;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135cabac67964418c07613fa6463b6b8546c26087ce256475314d98ec75d09710bde294a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61dc9220c51edbfbd42f7203cc86a788301af6acbd61c3e452e49a4baf4fce656542329f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1529ec06384af4f8db4536013d706e114bb567ca4788d47e81079f1978621212281a7b2f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1eb46455f1f9d795da3838b06216cd8d1de4fa8ff860596b89ee09f9801ff759c74a7be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1711246cc3260229e9467f47804a91de197e504d263da3981cd509d2988b3ece0fef6fc5c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d85d184ac60c5e09cdfb907376f457e10359572c06f2a7598b70c5d46ddfffa5d530b279;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe475f8266b8fd2fe1b59d462b61c71e41d8c133ed490b6147980318c1faa85d224ecd11;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1881c1d99200448a1088331dcbc88bd8ae44a80ee3cda5f97a9549e45ad946a055847885c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h157a2b4d0541d17676ef41f1b8e10e5f67ed141b58d055e0bda3e6d5d4a2d527876466e49;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h161a4bfba7682f0ebc317f98fca01c05a49f9a143ea8c1443df8d91df7f48ffc6fb5ec85c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7750fe441a00d9dc04edaeaab7ceec589f156281b9151d5258b51be3a022ba8e82596d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d77a91d2db85d581aaebef3c3e14e8cc97a83800a08db404a03442c198621fa19c07cc66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h280fdae60647a81afd1ed08726651cb3ecdae2e0802dcb594ceb3b475f4b4f9dfd853765;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb9a2db9acdc8ddf487941661d5e30a763671e04f06595095d06702a8b6234b89d3a1ca2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha89837da95386f9483cf2b20f785e99c21fcd3bf4cb4ba7c1f055f94aa55ae75767f2da4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb83d0c06657cd3beee515c7c10ac30ef79139a9a65ae4bc5ebd5222fcbf23204b8b81d59;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1827bf7a0700f7e31add6dbe4f0733c518c60b7c8dff3737d549d3a832c61ad6fb83bdd1f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea160596ee9ca5795fcf9140fb74da5f50709190193ae870de546f5f74bb1bc14844f39b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a53e93a161d806e5fd27db7e089a8a5a6c98b5b9e3d776ea4858d8a5c65516c89b43b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb555a2b5e640552b00c33364c613bdef9e1cd0317204b33e6fe4367f37f508c52af491d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h656ee5ac173fa137b2b512aff9f07d6f33ec410cce571d8785e4d5aa62da570efdffaa16;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38c3702f395732381b6bb3f5b002a0d1c902a1edbd7d51ae2cf156081cb28081578c3641;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b4153565ef4caea3c6f51df1f6bf65565e48f26462a37723124ab4c07c27c6d323cdd9c7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb507fc5207c892809e90b0536497683a88518361c8746e87e61bd708994671694711ab00;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9b3859c0725cddee59140750ab1d099a61610653bd196e128648dce49406d6d24bd55d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10c904d86983cb8390b125b65663cf90c0b09d61d9e2966e23beafe7d5f2121931bdb1075;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1507c91bc19741df44203d69eeca3fbf231aa052ef5579910468385a2018d3a1a74acbb57;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109169e6e8e5280e5a9f84fb4b7a11a24f22d06443a4a2496507557e447d215a7e7b8b191;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d5338010f054b63e55706e36e2e5d30727ffbe31739532ea6f28d967386a72e224e316a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h595555f0c6fc423fdfbe0b952d431590feffb30e9ff84414c1853a651b4b54d5533db476;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h149ebfcc877c9d5942a62c4c0b2a7fb361cee33dff17cf5505230a112a2a75551fc3625cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a80337ca082663373629a244752e3e22ffb5894d737fcfefb057512dd1bc86596c823443;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h485f674435492c9af993ec7e1a6aed0f710bf3bcc2c9f432c6c7633821daff81f2f8c797;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121311da0f68bb8d6e2a27f4e6f2b6d4089afba437fcb28a9ba96f2f962a15d5c1d810eae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11395a677a89cb7105ec376a3a57837a834c285f67af0c51cabdaf84028758b0bb560ddc7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbe30c4935454edc0e9404a756611f2e0a87cbe30244d1fb71158e8033c8a901f6e55ba3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de7bf046cb6002cd0b6311abd16c539e1b7a9c2d14b70e2aef793e705f6273dbe1f528f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h326cc5557d1aad1df424dd0386fd5ac669049b6d4fea6cfa16a590c06ef1e1630d44dfda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda15528915b0e4fecee75a43f2ebffc2bd3aea4b3967726c385da4f926a4496004a14801;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b561ac2729a5525c2091d31bebc91712d3fe5a1cec6684877708f094d4816bcf860430b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1150fcf5f4641f3b2abd5eb001cdeaa6db3d27848b3b9edacde1107533c47b8daf1653a9f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cf143e5d2fbcc5bcbaae8d86575910282b1b050abcffeb46189268540de12fb4bf1f54f4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3b1a901685d22e2721eed487a0ffd75eb63c7befb977bba11232d518d2427d60a323625;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf363369bb1a4553010834e2ec66a1d23c5465fa9115aeb15b23f5e7887cf91cae5e09639;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6c27866c0fefd82b008c201cb4297b8a5d79c1c6b8cdd0ab3be9bf8f72d6d10bdacd8ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19211676e5ad5192b0bb4c76edb12a04f21fc11f13f2e8b2a1cfc34538f5201bd0e33a2bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c50820a37d0858188d4eb4d6bea273f54fb62f354e9ba48232e20bf4a72872d2b7c1346;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h194a3784d4c77c45930a9a455546ceee046f63033554c39acf9e12f9056069259b09e76a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h146700db6b4f7a5dfd296b0eea3373f83eeb81291cd48e2369a863c7baa84437bcd36b0f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b43ffac81f8f6d0ae53fabb2e789923dc7cc28ea935635310b58e717cd11fd2f8de7f476;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ad3ecbd6773a9307bec2ae84b42d16e2df76bf4778382e06ae179ccdcdc1098b1dfa183;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fcf7c02b263858d5d7e072c8e85658ae4d87a2ff518b731168cdc11d9280df78dbfcc081;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff416845b79ca8ecdc93acc3b8199bff64ebe3cfb07a9c5f50649eef9f82de4963de46bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee11e963a6d47020d233d0915704b2792e0cd5dde94b4a95a97181a6dfa110aaf143ecff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1778798e807d0c003db15488091ac1dea1c149cb37803cd036803a93887824a21d65b8cdf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8849fd8801e6ac6e2885917e15cf8e445cf2ad4f5b5925eab76908a1128f06111f78b2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f21211d43b38e0b6b58572e9d6673188fe181ba6e74fa1764ed1a80313c827f5c4cefd5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9beb944719bde7b9f17c4f079e3e8f96caabcb9f5e4618e479cd80082aa99c7dfa1736bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6872596a43e675c1aee8e4e0292ddc2df24a126b593b9f1bd4245c929eeae9bf7a08c927;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed992ef41a2d8a341c2f67d410de387badb67da4388b6c925007ac2b57f351121c074621;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f36a2e0a3e741692812ce04da77689ade7053cc92795607e2cfbdcdb2495ffbc612434c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181b96a78a2c5a9b823b1030381d4c02852f14757eba364f587b5fc6c77a25fda4175f153;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64f3c644ee5e886825b3c6c6a8f354099b1c739481969e7f12c1c0c4a6346042834f57c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d182ce1c563d631afcde4c01cf7a0f5626a3183847976bc86ad13828ecdd546f8565298b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153ce6c948e524af70661a7ba8cc269d384dc29aa3710518b089f25145f43ddcdc67d16fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h600e19eb6fa268b9e206d470b047afbd6fb8cab825a131697b55120681a5cb9428abf63c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ca6410ddc319b2e6435c8c55955795ab12d2f403fbc4cca0a180af23918a82ba65da354;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9e00a70947ead702b45cc396658805b87e57f4f003c786cebd358cf88d48140e63d2f765;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a2e319d8a135743b68d4377368b94b6747edcd062155c04c561870863f44abedd1fbccaa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154ad3e847db5e7d9f27913998477bc0afaad63f29c2500478ed25343159d5afab9521c6e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11505789c288b7da6aa7090e4413d39941f42e2e251a31e772583af347326ac9576c8a2ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6563efa87c14d0497e309ad0a601bce5fcde8aaea1a694805b5f991a01f930d6667eb637;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152caf32979b62cb88d9cf4ef584c3bb885e248def64158fa564d067a6091ed9455af8fd1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91a3dbdf2a94316ccf64092313c645084f94454a7f9b3f41a1e2a25e925271c4a4caff12;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15502a78c48e7c748a332a5e45b9644362c22e69b14707855857ac0c57d626fc061b6173f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168048a26aa5bd4a2e09e34f683da89a9835a20a2c985771e592135442a732f968162c0b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10030d412e59bc5b85a5f78d00ccacd53e0a32ad746a7f70c9d17317b8d6554f07428a06f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d482c69530fa4a88a79922d19d1f73e7d7723d966c484036da7cda751f3c82e6ac5c43ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b5301765da833f14fb5ec01134ca3a1d028c3a1e9ea566b5d16857bf5e78b64560f550e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbec4c7454dd9da3cb957d370d782c62e6e9e7ee5c4bfb123002e0d9ffc10dd6ebf8705ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdd0a47e22bbd1d16c018451b20373ba8004417c7c82391acfb3fd40ad9a8dbfc60b082ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143f694b636762a022ea92812f72bfc5e8a3d9c5c0ab6d7a24389486cd4804837dee88796;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1087c68642bc3ccf2418e6447001812448b999a3f1be8d06e9ac572b3500353402b649b27;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1203fe175b781add6f9d205dab49b73ca4d66f88f5feb094f9f02d5a6c30f8ab7f953c42;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cbc73cf78d39cbc59b05860c7ad64a3abde83010b48cf415ed433caad02803a5e24d1a5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d595099252a2de4d87990bcf2f80be11bdace703f85e38dfe205005f82d03a3c1289bada;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b52cd38c32006d2c011136f4c305925e47aea168b263fed5c8dcfff576ec676e486d56f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h861a59af93e1c6e490976c424be620846a0cc3d84282870b5b85401f7a9e73cbfcbae885;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc74c588b47a248111d6977eb7a1285332bf427241966519c99d7db3f803cec7ead81643;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h103eddba9fe852059199af95a5e3a2c51f56e2766364f889b1c03b3c7ae2d68331a951f2c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e3e6f291f0075cb7ae3f6111b4ed31191834349a3ccae2489bd7a1402d0bb39355f4027;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2b0a0cad55137ddc87f42e29397b2d2908a06b567580dc09b67b255a46fdde70f883e4e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf96bc6822599718143c86f1b4d286313c3f6eb6ae215f12ddd440dcbd14039fede1853de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f10ce0ef859de1b7fc77aa0465b8edd5ad1cb9eb7108bc9050ae226a7676626e8c1cba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he153325c9bf2413b3251ff49a10e5e6ffda26d25f8c114e3959e0997cefa8e2c2d67bc01;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177fbadec8751a7152c097515bce67a0b25ac0d21433d46cc0f0fb5765e7f4d0bddf64011;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18c6bcf7396796892fc00fa8229c1da94db8e9a8e81bec41d53481b9b295f2d19032c10ce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6eb6c4d08b573fe2a688902e1fb9aed8efa447d89ac40769fc65d10274cbf2c3d559c29a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8506de6b877c921518cb6396c0f1f02006de8b8a0300b39b6b75b462d31e02a6da295b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he1b50899e4b16fd315e9439978dc1db559a8d7dca2f8593cccce116e10a995c6c87a6598;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10091a6ac869be47c487c9c861cad64e618ff0b8d4aa97d3b11e772c40fec3495930a5626;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc51148df774ef19a020feb48690724b398af13e234048d4f28a327deaa5cf85e16c81d40;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df33334d1e7bf8e852a4c29656f353400350f1a0c652043c00bf83f93d4ec22de55b9d4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2bbd70230cc09be9bb2aba6c3bde031e4bfda95b451eb03f056dfdf36b57f5ede90ba5e3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187223271ee55b03b9e44de07340b4cac0df63d2055935225f3fd47099154f256b2c03082;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc568b8afda66bfaaf0851d1225c0a3fb3aab27b1d36b4c3b2d424ae094c1d2db1c2d3dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6000315b1e00e123f6f670ae221b9371ba19fbff325b99cbb7f5afcbdbb721d72170032;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0f47fa10b3e665ca4966c22e03e23621e311efef83a3d522739d5a440b9cc176ea83644;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d2bf27b2bfa60ea10afafa116a921dd876b5af8291aa9540892a5b0d4f917d91148635d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1413374ce4b2ed63ddde1a454f3fcf9b022573c32a3f1f2cc702633f5b942f893a3efd7ba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec4945d1982ae49430cc7799addb060f87cd7ed8ec7a65cd41e663ad92ac1b62bb3ffe83;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a6b7d773ec563b552631939320b7814e66eac4271f35247dc0eec7a38aa336f96fc0689;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h41ef6570d54bf3ee0073d523b33fc00eef0fef9942ac2373907b33596140f12d5b8aa064;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1afb139987279f12b8f13b4add3afdff0b0e13bf8789372ff015d946f153c5e9eb22a699f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b98e5bc4351b6308cd9d9d53a72d37339c204d94f8b7733b05da73ea1370e8b08d3b68b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d839fd48676b9e164c9b50f1d13c6b36e60891b2d87dc72b1b2d4ae458532bc2ee97ec66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a84e8f5a411d229febffde5e1e5295be47fe97b96424f14aff430ad1272ab6cfd4cbf6c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d531c4ee3ee888b18776a5be95c15ea12180a01ed786ac7042eb86f79cbd00f135897375;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4cc1513e19edf98d81e5d09333f07f5a5b5731bac884338599b6a945834bd068efc3ba4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c632dc2549c9dbad404bb9aef0f554953ff16584a3c6288d9f3b34dbcf759d0365d59fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16590c49ef6ca564814187fecfd2afa99775af8c286903ea376968beaddc068bd997a6f87;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15ff6ec3f846c6e1f9c1f0f7849bfb577bb7af053da86558a4f41e4ab4b22ecc2384c8c32;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d61205cc0425df21b63137b5980e79a81a64c66e77e463cf64446f201e875621dd1b3e76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf6b432fe0d3bed57353c7160f43069b7ea1e1719ec4c1a5c5ca48a6fca40dda8aa6c0df0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h142e2f0aebc9a4772140385532e6a06b77cf49292826ad127d2ed35a54645014cf264c5c8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16295ff44828bf7af336c9d9a2cf7070446bb59aa3dbd50a97ddb358853b2ff481fb6064a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c3f4ffe5b03fcf36f9d82ec89cefbe99a8ce060682694b6122d94ff575f510358e54eb6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed7b3457e64d534702656f65e8c6ed97c9b2e3beba6b07aeab563e75084b926d74da20b4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d83e82cc29eada7baa368d3da1a2be7c8aa1365c392d9af2584ef1136f12e088f48f6fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hadf45bb48c3b97f3d485fe6e3138149c955a2634512f1ca9162e6cdd4b074e682575a531;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6916a28585d7a58dcdc312d714ffc83a9ea7aefe51a71ea297716b48134bf4537588d3e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a6d0a94576fb7f55a16e93d96af7806fcd5660133b2c022de3079be697ca0df5e65b81a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a146fa18ac7fd9f00f477bf0bd0fb04772d06ff074351ed2b3865140e2b34f58f20f6ee4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9e103ae94f2207761e6bf189362c56342919628a8aaa9a8e7debb2d071fab734fc945d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117bb71b25cf165c8fd57ce8a419d44adc899e8913a9d17b76f1db915dd667f18a6959392;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1ef3cb9936669a6074d88d334f5db20ab2e55a2ea9038ad8ea727c774ae11254bfe22e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1deecac5435f1649929874e623a2805bf80020cbba689b3978c3da3a0ff5f5338bbf8a4dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134a8c42f4c831e76dc3e1f71efe5dd8691c41cb54884d3d9e24e9aad28061172f1f9ad76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h256e7c81c6b4c0f9dd7872e081f7a14909c2511b7f1269db8c9b73d572ee4f223f4e36d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f63587592d5e8d488a000a056bb3c8f6fabb9b249850e7480ac63694b982e464577fe822;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b806e0cac1a86c73ca9e8e8a6f144429c71e6068d605fe53d1b4285f5b7e1af2b379ef8f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8f33176f7b6d6d9907953d973ef3e92fa1eccc508f17a7248dc433e30d9664829375794;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca695e3f2bcb1b8f6cb21471a0de0fff4190de92b8fb18bb692e13cfc8c22c16212a47da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb45db27b2f45780d5e13e0da401ffd1c3c4459117906c83ea1378acc8ff55dddc7378f1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119fb6903261eedec15dcf3763f57d7068cbcd28e78587b3e828127819da064aaf6ca50cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ffd3447a1a937d5811b8c3b3ff9157b12e85f2a2bd5a7c2a441b507a19bf2359a3d40aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db5bd61ef33df31b0b49c0df4e901d8e2088cf35e6c1f1a6e26eba78ebae5f98206aaeab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9450b39fa7b32071c75965809e1f3925e01fe41bf69596d301ac36398daa6305e2f711a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141d9b708b2ddeed52802eba0353549efdd1cad1b1de089919543f388b74ba6783c853d59;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11900c2254bbeee86e13a20766d698a5f7c79d314b1af4d0ac6447d6147f9d285f2da2465;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1640e086a60553fa7046b111efe9dccd12684e2c6b4dcfbaa1de2b388a8a145d97180a063;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dacd69351283702fbe9ef2d2015e3fca50d5d1ce06a43fa4a5025ac2c2603b0c2e39014a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc88beda358a71b25999535969ba1ff5d3fd635ede2744386491e6890cc35c5f31fa15383;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b67be70a5160005d84f1d2f1eb5ddfdd6b4941a0f31b931f35d04f80fd65cc6148738c8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc60ca2b8d3cd3a69b023980b2ed21fcbd49a9acec437c78c964724473f2fad5499cb6d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eae97f0836a56db51e84d8897e1905c828ddcd112e3dca9e1810bf9861e94fc058f04813;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11a2984a4689d27c75c94a4ef2dc35e35c27ba5349ef4ed5a0027ef0c0b55c0c29f5ada60;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156c98608857e0050ece189efdb975150f2c159a8425fbbcaed28b4fcb3bf6141fc2d6491;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117cc7fc9e39c79e80e61ac01a2ca28d6e8d4e7d09416c32fbf629fd92363482b24f46ca6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8fdef5676c27626c11528b3f203dcc5c125fb44ffb6a83597b84cb8634de4de07aaf97b9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1099ff6ca69238703c95bec3c0ad67f630b5383a4139e729af904ddd4c4eb93b076cbfa66;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h53d9ef0fa24f3a2ef2d4627e43fc507e15a4d213bb6d1f69dd05fafad251e6cc704b7d26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17410c3c4456e3991393c69dd1e696c5f29879fbbe55bec94e4c0856e82cbd7e47cf7a5dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h230c6cff1e451d17b54e1fb38ee53f5f755bc76e139869b72572b94287252744218adef6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3897217a1bd3890a3832c9851a97ff028c91540ba931528d41b1e496cb56cf848e33aeda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad8a67877080d2512b53f21bb2ac59b96a0bbbb743b13f1f6d54ff54a08259e265b252ad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7c6713e08b96da4acf217285c478ff7fff4d09cd950b538bcbaaa07c6960f0dd755cc0ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ede8b89a5e300be2c70ec846bf21505b0b141632f18a64d681ab12147d6aa8eaab27322e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1efd3eee43efb3fd95203f33e0680c0e9a77932d700f0f5aac8cca4fe75f21d5f5d06b374;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb3645e158b41eb80b7cdde38927434e33af2d93ed7e7e304cf3cf11939f7ec9e79471eb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf01ca8b51178e4444608ed7651f58a4657e501d7c7ef2cf8627c06739d17251ac696edc4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15af5ff63587e680046b44661b90b21820e8e9c790e708ee568b04d1cd5801fa849233274;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h937937fa867a93edf1047a3a382e9fa1428a8ae2a54db04cacad3f63a78fe8636857d30d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e1e88bc393fae95053999c49ee472cee6b95b30acf6cbdcb8e8935989636feb9149537e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1583c9f54e20acff758607d9ffc544f23aa480a452e3d28446880968b740c6302e015bd3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h110c323bd148d5b779014edd529704c3e8d6a0e2809b91e43af1061c9757d71917cd6d3ee;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a6d1dab8d39bde8f0ef686148769ebdb1d056c05739238d6d3ffcbfb43533c86c37454a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c5356499ada764e0079075a41060def01a659855cc2c18fc35060d1a2600523509e37b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d12d2d5945c76c37204cc6ff837d1b345ca5f03eb5d4295eac5a9982bc7276921dd83d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f40db1ff1a9684db73bdfa34401421501f9a98c525f0043aa72ca4ae896c7e003e404ad1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h93f3b199944365a71430e8c2d175bc910e924340d6cf7a7130dd49085cb154cb311ca999;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e866b678a168a5edba11945b744fdaf9cd5c120e22e2aad5ac312e4c07665cf91ed674aa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h514d853cb9296c112779f3e2673bcd2822358b4feff4c028f311ae24a23dc0cfac49ee29;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf7dde2521dce0377593e0a0d5c6bf0910035f06eacca698bf075a96e13bb37bcd8f68af1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a7da064b6084731ba16ec914996828d5b545645465dad481df448be009975b188773f451;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h191850a7a5f25d8376cf13a9cda5450240490c8de0966e7682d1dacd775918e8905667039;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b1c6a52b48bc71023ff6a59b28662401977ba6e2279674a0966b9bc0d5640c3ae0625fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6719540414da0ebf082a563244e808fd900447e95ea8a918ea2c5b675667702fc7a0221f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c5a204f80d5911e1b77f13047a3bae0cce8a0d7c39176d3c5ec95c311cf5b03f1239a1e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6993c18747c45d7aa72bfc3753eccadaa95e3ac89fed3dcdc0e9cc0076c0de86b943e30b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4160d23d88196d62491203405f30bb8191493968692c43f2a7501b06d77a6f55f7ba533;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7bc4f96f735b3308530faefc5f32d1d8b5371bb321ffd98be9370b538a04550d7787f92;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124fbf11e1b66175a1cbd174d505d01c7eb004f431496bfe338cc5c3e51a00d9699737d57;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18bb63c7bc853c0ab6e2903dc21255883f5ef11ae009fb676370df2672f756025a2d4a35e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f5aac18050b15846cb14ece18cba0a49d9cfa4b1139edd7a3485ba4980db8eadd9b84d1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hddb42420a17c262ffe13883c5aecc0e44cf1095256cdddfcf5c118573a0b45554fd4d102;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12540314d67c4266160dd0b2426c902c737793c27dfd9f6a606e3f787a5783a140b0f50cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a741d8fccfe2490c64c66f12d81ddf5c8be585f911826c19ba9b09c4895b584e51413def;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8b2515b720d2324c4d54c4276374f4d342ff29378b709403b0f51906728c7cc43644c26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eacc3cbbfba8341d502bba472dcbc713b59a76548655f1a7fa8656b20dc28546945006da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10aa42a0d9ee30d9b3655915cd4946a320d2911590f1a5debe1b7d6b0f7869fb7fb03db93;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5964d8bbcd51b1ce562f41eff3cb9345ef19d915af54923384d14c54600352a18c9e6ed;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131ce0b9d012767df4fd4549690170da10bc430a1cd464bf1bb2444a34bb997ec975d269f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h53521ccee58bf1490669c227ec87f52218866668ad77f1a6716e4e7dbaff175706441868;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b95ae7db63ab5b4d9cbd2a3c30292f7b6e01665623fa9cabe15f8b1c639d3f4d4f5cedf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e61b9addc5df1795d848b8f633cee914316628d9673b7811cc77fbde5c816db53b12b828;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17ba4c1b7db600de50ad3ed6f4f93470d7efcf8a93fc54502c0313c3c5d01e8a46d03ca84;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d906c04e6f6e1d0e7c666cad61d607c8b2944f7617adb9025d275c28d34dcadfe4e032;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h967bdbf6928c78af1576c0bcc4f7bd01746cc6791f9900e4fe1e8e637389fd46e0328d7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17e8c46ff404365146dbd00dd1f63f09aa3e5ef5af291dd91fa2e9513e7da193939e12e3e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a4713699ffeee7ad16e7ac89a8377609f830db35159b556a6eb77b52376adab705c1fbb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8573d44c9a7a1c1d921b4db096973f7b36cef748b11239848b5ae05ad05561a7e001b69b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb123cc13e9fd4a9253ac446246b25910fc0e7f98f2bb029c8cb68022a4317dad4b4c0ea5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cf47099993773532fc4f9f13802de49708671f6f6a150e768bdbe63321b9bcac56067f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae79dd748ef7d0a64343709ba6ac59306b27c95e5c42f3517885480e7e51000df0a2fce6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5891f724da98d3e767a440011ab08f7a350339e831d3253daebd02e76ccd0d8897f1684;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fb53bfd076a9cab8753bdda02c7a7166880d204fb94e604dd17a8b8f80f0a486a4deb4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h605f71e10d3984c9cb884e7a2b8e713dc3f10f00ae424437a3c661fa5c22ed8db48c3a83;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6454f0824f353d2f9d90a085db986bc2a6366a690171b2eaf5061b2d4800513f6f6f397f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b4281265467a18ecc87e7a47fec59f4e3e63b9f0816b19f6b86d77fbf0b6387f2baf28a1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17467088481d1d62064352e27c6239661f0915e8d3c5b4e85dadaf6a1e67b199fc00f112a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3f3d88e33fbd51f409f188029fcb4f4baf7a0d42ddcca07188fd9734b7019de28a69412;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90f9b70f18640c0eda754271662cb3baa337f169aaa1a9bc5153b3d3ec5b2048a071d425;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150ac7cf86c5834536e3c47a2d266139924328fb0d3c9e9eba5abab5bfb0b2f001e56a324;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a838d1f85f71e709a96312edf8d1bb53174a4581cb7dbd0995e0965b7e08a2c82a49401;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1563d95396f7d84e759b9e7719d787dfd7523ad76157d73a5dbb9b0d836dfd5412891594d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150f22159a79aa0418b6a10329ae453639954c785b04beb2ee4d461519f8a0701802b38bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf730939e251fedeb1eb547fa04be3c0d542e4ae562ec4cd6f9d5d1aa55701c111ac8da41;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h148923f88dd54b2497e4f5e5a39ee302d9f06c8ea26964837cc4610229015e77adb172b26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d839ea74b88a67d943b94def0e3ce845291a5f2872d285ccda43b631bb4fce41db75f61b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d88df1a546d43c49ff4b707d5d14a31573e279867b083384f1b5fb6d2d6d7b3dc9c08bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20938d390a71b016b8f2da23e2704e49160e6b6bb3d3400409bbe4d4085e0b3655e0ad94;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he574f5419996a215dd2501cd3b4e80ce6fe110f79a7efadca4e06ca7941fe8a36d0e1b9c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c8f25bf6a370973d88667a469dd54a025f200c9e73c49c1e917d9eacbb2d054038d68be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19667f3661ad1b9397ccf30794c01e078b496ebd84da150bee7b35ece7441cebcfc7a7ab1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e28b737bd2fe666a70688c8499e9878b06c6b79c52d412c094826a8484b9af80d910d956;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16d6697f7c8feabc617606a7a1e44c2d042c81809d2a662830100f9cb0ac81437b8188053;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5c6594a83c5651ed11628bcf0f7964a5a19169eeaed2f07486401b76de9df1dcb8f08930;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1638a963d32834324d96448c772165d244c3a5a7856d1d1198346242fdc5a0b26620ab07;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bc66fa90b5a17c133b57e772aa8a98631a4a38477348cec9c2288316a4297fcff4921b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb363ad3c631011f79b031469438cebd2f5a5485542c269ccb0de3c1a25502de292b7118e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b2bc2811f94bf69ccadbd5c772c9473aa545fc40b2b13c4703507c87a4300c95730d4bac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7f0076809f1b0dc7d780655740e67e30ceaa77ca31e25fe626161651efaafa2f684ac4b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1585f8595f1388229fc9a9147bd42bc21a7f5450813c71e826dcfa9a968349b831ae3cfdf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h786637bf57c9489e3503621fd3750c7a36c4c55a715fd9e3319f5cd76d78bf8a3f3dd986;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4404fac03f095bbf370ac327b20b1e381a1545df5773dc9f5b93f90abc0035ca26fb2100;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3be2fc3f00f33bf47be21b484a415d2cddb806b773d30a372b099dede7b7cfe60ea8169;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cb8a974e19c78cdcf117f82ff42f33853b84b4e4bb16b8a6be49cedad5fc5106fca685a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7963d17d06038201a00da714d3d95b35bb1e152d6e91e08b8b5cba29d8ae5b5439a08d78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129121b4f0b1cc86cbf31a937cd59b33172a3311d8dc04b24e409443be96c0abee450a756;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2c96d22911e06bd6abf87383dd51f9dbc058f79c8e2b608b8bf24773f775408c63653da;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15788eca3184d9b2fa0a6ef29442cc39369d39fa4499c5620df86ca392f29750298acf21f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e2fa1c3b58dd08b8039b118b15cf1934fced396854f21fc53cec3d2d90a8524aa426242;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6cacff45516b68f9029186b9f994fb4272576315197d4a304b5d749fd9452f67a4187858;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18bb8ab525ca3b9ffe98a0e0cbfe9001b6369ea72f7cf7de55f8c56b848ec9aa8d9295a35;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de44fa629ed511d0000d2a93817c1a4674797ff73aacec1d69da5bee7be7d413c321d7fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155d928e70ee13a811d68ca906916f481f2b8289518a7c282207aff8715eef4c573064c8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h567f0417a71493fc22576fd61b5181a18b87d73dd7f67fa972b27a3398d671156f915306;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb099e7f05ebeb198e39b65197807cbb6cd383840946911fca056716cad5f165534c20bd3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16754239b1031851b6557bb6a975883a41e5b0de708432079bcd384ecbc345938c13659f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13239b75e023c9032f89fd711cf31b3d20bf2aa05308c387a685dd02fb2f8ab3284c60875;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c5542768a710f0ab5bcbcfc2ccbe2efe9e896d89a33243b9196c6835d0c3c9703806e9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6bfab84d037dcb8770bc048a606da54526f303ef0da4b09fe726da26fb63148c3401f71;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f1d497e8d3462c1558dea22b447d0f4027477c2c90f03444c263fbba3e43acfbc4206f9f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d02b5b4ff701bc5323454ce1ad2714de4acbe737ca35b1d8068f8fda3a2809680c775a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he609ef1a59c6ad9b02fe287281e37326333438393b9c98ce7644170f8818f35850accabb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195fbfe00bce05f126c7a7d0378e04495cb403e580f2eaa340195e9db4f66f76ae53011e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11be757972bd60d0c724a2d39e945900f473352f99fa375c200a6815ba764c131dce0b7f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e31bb3bd0930d4fd7f4109a45187160f1561dcbdca2d0d570bc0037ea08b3741e5fab1ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cfed5d4336b8eadc298d8f8d51def0dce83be313343f2e1a887c31220acbb5df3dfc8572;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h559d9c02da70213c8ae63c14f7bf5ad7bcdba67d5b5332d3942219680baa4510386ccb12;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b1958fe08126cf3d3a4b2ed34a9efa9599d260802e9b5b2cde18c89105c7b0bc70ec119;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae507ed0e57078f1cb322d29468c6a65eaeb26016f068e715c7d83c1cbc7ae9e8198c647;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5b92201c4010322657d822060c79566e61df06c16892d3def0cc80e464707e9d7063fb75;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha0df8663a1ac1acd351a8e2c41e135d03b6ee11f780c0a36e67061218f10fe231507e28f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14fec138959236a5407620280459cd24d01087e6686de7517045468047f9c4f54d680b375;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd89af71ed023be4759ef96e096ac0c4378dff3f00c58ac245a03120a0d2ce85dce18128a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c42f94e96a0053b19e84ff63544db2c1577efacfb56f5ccaedc72a88105df700cfe2fe50;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfc153476d4fc36a241f480b631bb5be9167d1278bb546c71b5c0282a28114744b72ddb8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba7f787da96af894f850ca2f5cf6ab01eb2f586cd193f0855567c67709f58c7acecec683;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h357c851596d031e9d88935d463481b0a8ef5dc9a20ab2d91f65ed6039c9f0cfe4ad9bb6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1745cc39089c1e8e7ae2a4fabef86a15036cbab8b2266cb72c346960c8b188253585a25f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12af87ad4100b9e5e8cffbde09e503d6094b44366ca400b8d13d96d5f772e9887f327b4d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb02cf302371cb82617149abdbafe0e2c3d759a80e092c909ea03b7ffd9719e7b5751a9f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a73510d0afd82592ea5f30810ba4863d65b0af946595fe4607a84928500e3570e982966;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3cfae299476146f837e31c33e10508eeba3173eeb4954c2aafa93807c0ae973160008714;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d54a868fd8bacbf3934f5d259d10d4fb6ea546677130c25192e5b4296c0df250515dadb3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14650cb1bc5436684683d395e7b939dbf9b2443197081a87357bae1a448ac9544a8b5a574;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6a651a55e8a02a5e209fa8247f1d6d580bf4253f19463145089e20d7b110b5ff530ad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c4615b5b622106d32a6ed2f8ea599be312b4582dcb12fa947b825fcb58ed4badb4722f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1602d8a16815fbdaeb35361bc0beac9a233dbbed2eddec4b1e6928cf04525da06c080b1df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cab8ed9286acbccc247b95bf3be41236da1321a32d94408a331f5ab42d1458d5cc08beb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa1ddc48f3aabe00e3f6b16514536716f4760cab3653d1122364a72cf85c822b51c027a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he8c6812125020a964d850603fdfd4837d1d0dfadd990627f0c8e5eedd1ec5847f7be36b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4463de72dd76e045e80ff27cb5e6a2f8a2b1732d4a5b84abe1fd74a0de61c677e5d1c0b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3da6ed3ff7ff7497847594fc7b230c702a1bcf89104fe73e88bb82de3bc70e03e5b7a16d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfcc433b3431263cc43773f16968011176a8f1be6cba2d335dd726d7d6577631732e31ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6eae04735b1e2c2ca27d1f21f1dbeeece325326596b3f97baa3aefceb84f29c4917a943a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf3619c6a871b24e1f2a84ec7e58109e999e7b1d6bd560f743346c78617c7c1c63ed1a012;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1999cf2b4427f24228d72ded2a3baafcd83540090fc33cd92c7313fe76e3d2400f3a5b981;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5e21f240862ecfece2d7d38bcb7baa5259d1f483fd0957924fdd229a1f5a7ecd96793e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a2963118b7c83996b806c26aa9f6d367e715cb908df7e2e8d1741fe52c73444747383b1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h110677835b9c051f0133ef18013a558ce6076036b9958d2dd3c4da1acf9667092ae4b9622;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bcc6338109de7cd88838d86c9fd110c362ccac9b10a0c00779f04de153a10884d0737e78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c5f5916a7dc943d8487d62fdbf78fe62daadc9cf510c1403ac6d7a69099ab30fdf5b274;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4010843a412d5a812f77ad19a8b8faa7a79e140ed1e8782a00ef544f5ead4e930ad1be1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b38f4df0ecbb6148d83eb513290e6caf6208c382e64a4bfe1e7767880d26227f594a0c91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfe333a923f757afaa945c04e8be8f98fc238c12dc3124f3263d19bd2fe35601745c449b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1861b67964c5526cf58c5858dad14e285bd4cafc1f335be1b0c979046f23f6300212c2b43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h99b56af691412b2f6c14fbfeacd543be5154f21209cd0948234a7c20436c65eb7dc826b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfa60f06896e5df3ce40e59eb8a05019890a18f930da18f88b584c7565f28021dbc7b2c1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9917598f859f8d21fa7cb8b98dc43bfffde4031b272a70a2dead2b65e950430dc2e6d99d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12fc2e1c51d3c944c1b734d6ee4ab287a4309309a729e958edaea7c5d815da3762318390d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd6d607abf1280e8944bd484e94adaec95cead1d37efa829f5ec5fb8492ef198c7eda611;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b223b7a72a7f0afc928ad995ee13e505a769324c4fdf83af0d9c9e3bf16347bc04f884d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8a921151e1f8eaa57c75450b3fd2cb089689db7663364efaac43f42d8a836072698e7f1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h176fd93022f12b125bbfe756611945ce79688d317dfd5f9a0ca7e229ca1f60a56bcd0026d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h43c0f4b3161f4b95b00b2ab0148118a19593f3bcb25e15bc8034d16d1081a7ba5b9cfb2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h93d43e71727c71a45af109bfd8c501ae6583df6bb9591ee51a55333ef619091d935bfdda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5d409ee7a48cad48d8bcbcbb7f8e1940d9bbe673b1e3a63b8bcd6d84bf3aa19b992e4027;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7df93c101e80c499c073e3ef992c09b3578d9d472085dcdb82acc064b028199371a6fe9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f91a9902931bd32a3ea587c6d67337446031babbad200ab47af1f7ced9fe0a3ebf2318dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h528049858a00a04693e115fcd8ff0de08dcd5c27dc34e2b40ca1d35cfade8e77271019e9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b1aadda214a9ee25c541c61e775cfeb2e5b0296bc475c1e8425626f1b30fcc11fc9603;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1828fbd7a68a2512fbf6e185232a60715c048d0f9436fd2d4d8613ee7f81fb250fecaa5a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha32f491be9f67073cb14290656709338985cabecb8c6aa82be501973e693e377014ea5b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc5f62fe2107471e0d24c23036c105f6d8fba20cb8845a50b504252c5319df0a61ca3d5b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8926136a9296d54aad09c39c03d341355cad529b6e81723a74eef500de42767193ae8819;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15a291c1186a27984dc3f90d4571d88f77c8a7bc46339530b1b488e345af497a9b93bc400;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1413469cfb87f4db71f7c9cc4ebefc19f889b0870687c3cbb8f41eb4dc5008c0b1d89197;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23353b28ff028464bad2d04e82b96faa153c6632a74def6b2c6def2d1152afa5711946f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1456398febc75318afe2366dab9a21d075693edde3914bec590be066a41a171411b14eb02;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f56c738377a32ca7cfd16d1bd8d83ea7e3f9c45c2957188ea9f40ef6d5dd6b1974eb02dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f24a918f4f378dcda1d54e308c88ee57d278623fe8797a0bbccc3724e5f126a4b398520;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6e4be84810cae9b9c3052d8bcaa9cccf1b0b9dc4b6a1665f25987141ec7c7c3755ba01f6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he23d9c0a5f2f2e3d094c57007fe54fdc4b669f18d776cbe8961e9680daf0d475e000a396;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h132e2843949f079c387a16f3c72f6530f1b23f0f222dced1417410967f2ff5cd85a16f9c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f98b98aa6145fe4ae1801837e03c85dd3a4213dcfe4357defa83d6997e1e656d23d2bad0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h973fac4ceac296f7ecb07b20adf3bbb4573ebd1de9cf2cbcdb891ff3a53494dd98e941ce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcd169f362689309fb58621689910989785cc111149d77bfb2a55f0bbf992e4dbb76fd22a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha4d5549574ecf5f0ccd26dd3119116402a760a1a7574f1029e010596789c7af56d4baed3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7045423ac3922263a2d9f158bc5dcff706ee017a698ba523f979504711511ce3e8fe98e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1920c9c2a17e59b92e712bb0b4cc56f380b5624487727d329da1f00f6b1fc18fe50fd1aa7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19286f9f4efb9282c56b1230245ea6311463589122f351d0796cf8beb8d159815ff1ed378;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8d7d39ff25cb9a2ed8bc16904aaa5bbf8b05a0b8aba26161282d4d519fe12062ffe5ff6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ad76fa24a5c2ed9b71d6c4cfcc88b57732b33d5f1f64674b4292bb993145f352219aea7f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11b5eb9cd3d0e0b41bdbdff29f95239669189ecc0caab9c9504b8e69e564cc60d7b52fce4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f00b61f63ba4d6ba451095a85fb9905e5ff20e7bc6b0fe2092f9609765d6a97ddb65578a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd3d70f57e69593be5b4941056511be1625b926d1e18fe06079d40ab748afc9c3c009202b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc948a92284b5bee111686e6b6c5d8fe675dc6520457a69bf627e3f04779389edecc2bc7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3587eba642f828502d80b914d6d2b9f0950425621bade41d32a88487bc8ae65942494643;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11facb13d4157612d65f30c64bb45203e3aa15db620921431e5c0c194b5da9668f7c00ba5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192bb4bedaca486af78acda849820854970a3577f29802c5fa7964b16da2178a8de764930;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2834304e00a8a688f2221a3b0148102aa726c332b31273d8701a37b14aabc3e4cb34c9b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f0d33469bb601c2947a9e99e63f7c75e0fd41f10d0a57891f3cf4b4ebc6555b9c8cf0032;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1289a3e9ff70e0c5ad121e79ef5757b1fa8b511674c26f06d50088574cee064905bdad5e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h74f69adc0ece61e22502b600edd6af5bd91411b92f9083db42058143e49702c976ca3e6e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1a92a20e2751efc5911f5b0a68c94d87cd098512803d2973da2768918900f35715faaa0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17aa2bf945b0ef03f3ff2021b062d302414ff1d472945d4d9ecc94aaa76d10fab7999fbc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12fd8512b4290ff970b5544a6023cac2103dba49e8786e1743015160b7c35d1d79f084257;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf6d9617dc32cf01d58412bfcca835a965c2f17b94a8d6e31f12fe6825b683005215c4d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h163fd3d541d6b75d96a8684458ac7a0dd7e818f44b0c086a21bb494985b2dcfc8bf83a558;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2fc1387218e99190d28cb1df8b55cb529bd82de5a0f968fb1c8f74618d8ec8e0f0d64e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1159b027dcee643f5da1c5e52c009b15f4e355feb687f777528684ac2edd54a2431b62f80;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d7b961950dae669daf7ff245f1e5d2a04105be0c78edc42de4cece3fc42222f85ab542ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had49110513d9dea227ea84fa716f59ca058ba55c3ec8becb125e660b27995234ff222523;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4715678c39e45c229a82825e081624a824dc5138b2ff4ae1c1fae90a2fde863761bba2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d12f4ee35ce626a060347390d48e8d4b81bf24b2a433085d819a22078d53d3d031a9f437;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183c32473363c8fe129eba46c93271a148875181b27fb96b49b93e8fa56dbcf76b2325c1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcad50e653a8b72cf46323d61b995b154196bc8a340aacc236fa0982dedc44c1b18e627d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdd65c4339821f316da3dfcf0da8a5732e4d7c4cda6538b11f89e0b22f7efe3b4400b7e56;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bd189d63102309cba26861fc87a1f2d796ba204df6e1bd16af4d964af4b8d1b0a0e7fdc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h186d4a659c1c1606a761b0fd05b3a9a80d9c9da4939f9855ad96f24ca0db8ed8c70837f02;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he58102bb590e007a47f45831631500c0b125d4df1a746ee4749a504816d5cabe8a3e10a2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd4115fae6540aab94cf1a88ac6d503cce08e3aac01b8e6c18e5d50ff6923f35c675426a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c475ad2707bbb95b5cc77e74ecd14609ae413b71bdc3824bd8c379b1396a85727323f861;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a794a8d27662315651c3abf719fdf6eaa7b76aa044c0611c4763a120601fb540312b090;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h662d7e27d9b093f2ace6abc561ca06be0ebf17a3075014f28a1a06d4e39cbd193fbbcc69;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdcf21556d071c3120069c24beab0be1c2657bd87fa9c9af5c4bd337abd990e8a52c8a7d0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9bcfbb9c1a92ce02e2b521113925d0df5d0510e1c308292a4cc908c21e9fd8488b30d89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hedb4d4017962b78e07b57bf3753d130c85602cf81bd5a1a9c447d4382710cc6d93a1af9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h142376978e89421b5f3a754effe81ce6064f28657be2a236b0588183317992ef7cb08d664;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cf3b1707121b6e6fdbf9c0392ad1fb21508219111db828a7df3f6d695b38a4bdf6b5025;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h867c67949046ed95ce845243c0ea8a3ac47cf3134f8eba53fba40215f82c004a8f868cf1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bacb740b09bd975f0eb336258908de71eb1f14a407c37abae8b1422134541d049cab0a4a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h952283fb0742cc3fea692256d3eb52bc5dbed677d120692550772a4aaf0cc98b76ede1ce;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h921cd3c771ad0538ae99e1d1f7d2102a4a7891f49456fdb23cc21e8edf4d0a486abd7ae6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f416da9e025c8169b5539f2d23d1dea1b2e6e9efab1bb9c899fbf4c9ceaf3374f416615e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h895e38b6f721eae0bad80a8b06bce7566dc356b927816beb0b3fdfebdb49ca0f88d14c0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e5cc06651ce7e46b45a44835111773edfe5e3cdaa4331ed893c697253dba9c599643b38;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190056c37db2f443d17f70bc56dea40ee1912b06ce7b55a6f79abf5f47750aa11068d0fff;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7fc7c507709422beeb6f3e080770fafa4738b2144edd86989f122881ec0089bc910808f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10fb5788fe88bdb6a978c2dcd3cd61c35d1bbd6451b70eaa94ee1304e6fe9f732163ecc08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cf767490bef825369f39ed37c684252a3fbf53dd8a273e1970124340229c3fe9cfd4c74;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107fa71489b75614762c6c09ecf6461bec3a83586a4fe006bc82b4522c97ef46a236a5eb0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139818cd40cc36d854b0fe9be9f69d2aa5b2debf2033c16e8460fc83adcd718b0a12f47af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69230f0c2456b30e739e148877c02ca846a9833ccaa223630f57d15f089d2d8d75f9c688;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b5d463a131754938946c15b9c6a371ca1d6617ee340277fe84ca6a480e8be56702bebea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd06a712febc823c717535832f1caac5d2d435d6c0f7752c41fdcbc0b7bb8e11cceb8ce91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d1e72eb8a29399a41cbd729dfa99a687bdc5f7fb84874041a1cab5d4897e15a8ebb5fa0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a92734a28f4fc58ed1988a009a6ac6d2de832321bfd80c359916c612697fac31485aa65e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc826044dfdff669676ccb3224115753fdd4d56c8ff5f2121da910713002eab1ee585a56a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h902f0b1ddbf418111838feb1141c4a981d3a82c553295e5a9c38502d298af42dc9fc2c1f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a7ad2fe279e544242fb371082abac3edb58c2b508b9b4ad8ffa7a91db09099fcd1d8603;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b4d7b63c78d7482a43d490a1e810a9d2a39e13f57a98689d9b262064b2aa42be3ab4a18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h41debe3c82df7ab571556c7cdded71c468b4223b9ac7855c8a8c823a22c7d4d6569a048a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h29fa287e7e07d97a1260dcea54d066d6ac7a551c2946f4031b13216b6d307bc14b312d2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17025c5aae1a2df0231e6ce4eab6f7acba8d69b7e207b79f62256e1f23425f391d74ef029;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae3d443cb779a60ecdfab6e26c3a18d1e5a6f91c68a4332e06c5ad855d210ba829102ab0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60160d2a25e82d8ed220ecb8663f5d3caf90b78b04aecdabfd0bd04cfd247393a61dab73;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eb7511ad1da716f240bb6d5596c1f2973515f91132d1f9aaff37ff3c8a66241614b34cd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h52ad4747aec7b3c888ca0376f9b76fbd86fd0a3924ecc980022d8ae8f5e12ea5aa10cb53;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb407aafcd692d57a8f80a7b00f74558d8126409bfc72831cc3d26ed40b44118d303c819d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de91f6af39c8580c1aa0da272801bdc2a628150b433521507b1428bbdd2bd73009d24055;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h21b01c6290a65c78267af2162af3523e33db0575a04832ceb08cde40a58742a81a84dd28;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ae7f565ae5b5af03687544b546652467acf02450fa98eb5929472eaaf4a0ec9edf1f103;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4518d9ace321371f8ddfabba20d91451a5b397c31cf2f4ac0a04d4a9d7f714a8190e240a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19ea6851c41d8ea4ca090284aa7198424701574e8779ed62a7d5da6e42a6b1bca64e24f6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15dbb8f90824b3f5902ce697d249e4db6cc4fda5a5fe7e8eed72bed991bf21d30db57c599;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfaa4c2b74094628799dab15b634991f0b69e450f5557c691c5a6e725130387e10487cc2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd04912fbb8b365b863e8f58f5a47a24a104e9774ca71ef413c63740b6d1b0e6653f4fa9f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha4fca15320cb019fc550b49aca48192166770e15292ca006b5c0c8fe828ea402120652bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121b109e3613990be0ec9fc53d39d4ae3eefbc21db3a08313313a763f1975e8341f91a4c4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19b1a25e866c5a3d0868300aece7c64b3e7a6e61ae11e61fd601afae896a001082fa49277;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ad239ff3aacf01b1453b9d9cca908a338d021bef9bfe0b03144577f1de539245b32113a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1524455b9a5ff2e30c3f306db6af404dff7829da8ecb09ba883ce8d9b32db634a7016bb72;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h550b3aeda5f9fb0f4449d2c7cf1417c3c764026ed33ba92ccaab792f1699152e7e1a0975;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h70145c2c561bb5e3f9afebf95761800fbb3324252e48f2b571a54b5ea141ad2b183abf5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h93613f14b0d26529e8b657086738d016021cf1daa61d0157a60a65b8a4d4fc347bfbe897;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha7111f88b96669569181f0b0b00a8f6c78270afc76fcb9eb04c42fa1fc4807244bdbd0a3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1578f44ef47af5c1deb87b618e6b25808a7be3e6658cdc7b093e2077fc3da11b5a50e2620;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15925ded4f78637d2adc140bfaf59c5051aeeae874269f7c04c3772650b8d95f4080c986b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1294831b3e322fb091b2799317ff54a95ce16f19e0f183adfbd1ff06075df776632761c26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf222393f5f0cd832954fadb33176b2c2716f8183576dbcc78ad0e895414aed21e322cb65;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150b44b5b2d265e15325fe691fcfb6abdc626bbc3c60d8ff46639599e8fecd7c953f1b4be;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4007cf6e2d7b6c40807fa45ae3233b4506896e36a81b525d031bc59ec81a9a37ff15f647;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6943fdebf3a43cdbe5968a8d09b970565da4a8f9d9f062c8b41883678f9537c65c4708;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a7ae1576a0c661aa955893b315d97985751e6c709699ce2e67d3f89c449b0cc1df06ce82;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160a6932a414a2f643976a1c11c752a00628df2f4575f0dff58d3d6a40ad213e46e53ebda;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1970bc85fbf2300a47683357f7c55feb34e92a4ce549e5de4f290a5ba4eea6e073260af5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e1dcac898d1b215deff3ec13595c3a6a16d893e2ea7cfd19d6f44d8a65c38d09544887e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1618ff796edbdf2bce5c266c1817a2baf3fa252d1301575de48574d09a2add88db30dbe1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d75c8731dad4de1e44bfa2e07bfdb24ff6c421957c50a87743aae108062f0666789d379;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13fe58867e17b3332181ee2e5441064ca158fd805b8e64ade01fed94e16480b354f08b254;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12cfdd96ed862883060c461235d6c3275b3d53a0e054df26dc3a50f0bf1619fa9bf48491f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd228005d9aac1691303c9392e505f28f60c87d8322981a6d35a5b976ea4efebfba91442e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8c48f9dc16777895ca98fd26e79ab1ceaac74911c677bfb271a619b8ef5a35d4ab4dcba;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b5a11e748f9905b74c4c270cc86006c77c118909ef981b0c88e089ca50105634d895491;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17fc0d237197d0cedcff273c9b400d9ed03dce8c18bc45f45398f46b66c08c2dfefc808b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h292dd63560c78342a2df640a30740b9b74a6d398f5f2c4d6fc872e4c9457169b848928e4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36ab004fb50de4997fb930cc2b1b0a1da2e475081bbd26f657570d68d6aa889a177ef1c0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb4b366cbf6ef8d226f0dfd86e6b0ff951e18d7eda03e1cbc8337abca2bc17721dc5bd363;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5ddd6b5c4db939c49bfdf43d19a7693ecfa1f1cfe69c9828cda54886546e94a69c57756;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2df1c366e9441d794c1b124f6b03672f652ac021e79bb7ad7db5a55f9de275cc6e3c626;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h590a73ae47af046c846bc164d066fa4f68aa4a9d45ab4bc6db107b2aceb980f930e19173;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80d8b02c187e5b54a9bbbf43b4b6370d0e8ce7d67a93d309800d5271f03e206ed76ca944;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11188af5ef1c5f8b0fae23a57e579510d77856c76b51eacdaa21b76574e353013c0871751;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1204920681fd0a402051ea57f1a89ca0f3b42507d7a35ae6f04969272081d247e32f53a62;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73f1a6f2146cc8be77847aed4a1e6f149db3827f6b1386b546dc82726ab240efac72dfbd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he7cdaea274d593063aaaa613626d22f84ff13c71135d60786578f047d94268a0b12dcfcb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h150e62760d885225d34724bcda34113f83c024a133a7443fd7258d19d813ef333c399a29;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f05b512b15e739abcff9dbfb09e7f048004fc309c1e4dc2f682e2e43985b6245db278399;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5ec88288ce4c6bdbf875c1aa2c988fbed09d77227db374c0ef5df14e5e9865e9e825445;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h58779b51bb04be23aaab7b62df3288f3d651ce43bf6fa013f23b5bc73ff57fc9e46c7290;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h625e97e14eca680415ad0c71788cd290e9d116257ce8fc029aca513a7e923d6d4a254c26;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10046afbeae564db5a5e0e3ff4ab3a07e266a17e9718159a0e4bd62f8217399ad4a3a6220;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h24232007021db396f9b9c4be0aee66b3b29abb836cd54ded6e23f9615607f9baac9af6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124b5ff268cd5ed7f8276fc8a7917c180fe2721ad5891809d691dc0f3a21e6b80d09d8624;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h106b0bac3bbc837fca601e4efa8aced538d374e43c6691eebc3a6c1f1b1b734206e49a21d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1267ceea8e712021e23e9307e58e4bdbf5b8d6bba3d6e4c248b4f3f65270309af82ec99bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdbbe5adf5d366e91935c31b3d75696e747980492242a95e19041f41e76d6a1353d153683;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86e4316820c969f87279b3a4f2cd967ef83b2c0d97dfdb3d2a457f33a5023efbad29321c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f014c7dad9b60ab82b9b63d2c46052b26621fdab5cbebc8eebb6121231cee864ddcbb9e2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3f6954b0003843e308c15557fb6467602aaff738113e62513d2a32b323844f1ebff9079;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c17bb79c918d0aeca0cdb3271ef9bc85fc0dab10c7b36375750296d9181dd40c65f0218;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16004160fd0ffd79c0659ed6f34e2304ac81d734539d9046950c36f5f695c69d4c01f3344;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c40bdf18aac70340f11efeffa86947562b672761bae9307a32589cb319514e93d01ffa74;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h83ea80d34dcdeec037a0d40137f665faece1187f67a7e79c20b3e412340de3392bbe97c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1067892c9fa394a1094ef6bfc9238e6b3d25e7b76893662786ba6473394274645e15b52e6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he743f57dd8410f1ba01299b6c7ab18c5b02b5ac7f48e1790f660b8e621e2c596a475cf00;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc70e0322729325bfe105e666f7613478c0e555898b244b47b7c4584214d4a24c6c27164c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b6a9e18a1a0f3f6e8ebef29864ff1c12df5cdc25e0097533611761d5c869cc9adb82df4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd3de95d954f05876355a1e6c71472b183ccf181cb69c524281ce9be83ec57590eaed0b9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5df73234576a7d3495633250a33d031d951dd98f76f722c5325a92a17c5e85041703bc0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f193755371cbde5e8399cb2999e63ad7f33043c48d4b15ef690a729d8ebff4df682c021;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h905f3e69314c382c34ee1c34da7398316983d60f83ff8cd86d1cc277e1e0aad196beb467;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3f1e9e65675e9ca8c43b9890876edf4fe44e76290ba37420465e0003c74ec8b101c7d7d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h969aa98e2ab4998a5080433245981af75505270b28d48e05102b0aaee9f3a715e3cef40f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10bb88f2f99a5ef24a026aa2795596ef5d84229915de79e4e8108a74758d4a532e8dfeff4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1127b6adcd98bb92f9c716a81ba1c6e2797f613e5dac326ea6b636ef4f49dd3b738c2d72c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17337ac06407d9845f2e76a1d3e5c1337c8402b98e0f90150372a88c16a79c8aba63604fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'had1e65bf97c51e27e0e2f7a513bb05a8f6da195c542403e239893ea2b641d3e0db333004;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118ad671c5658413493db4f5b9dda359329cad59116fcde62e45c5c55af98554d7dfe3952;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0bd895d285b40c5db4c2b58df1118049d7c830e1d039d727c78a1640f23a9b74b2c3252;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8cf4e8cdca3126f2624f8cf7c7b791ad0ca12334e2ae7969528a80bc6bce1505fe59f613;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19148663b7de8e04c9fa516d4b460a4c1158eb46fb27b3113d9eae722317fb78214b99e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3a159bf5f3292a2c7bf95219cbaa1085ca2aef4aa0e86bb1f295dc41acd2ec248c11312;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11f1ef2e1aadd471c83c7cdbcfb31735781f47c3a7f87b1476c225ada0cd7b029d1b08fa2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3eb93cc670a257209ae6583b8a888bf0138f47019df90ff1d93b612c1672813d67f7ac0b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2dbd5abd6f5a4c00e3b4cff35bccb456f9d0df9e2a9eb3b5d3fb1bc6b456a15553ce1996;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h754e730a0d7e5f4ece86409d66c175467af8245214096201fad7627b7895cccf7c75add6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcab43becbdb7781648615ebfaa165301f951234c0aa829206979ee91a9bd475f7a0744d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86d2d1dc434ee2cf639ddc3122ccfa2db51f044a0d15fcffc5276131d29249ff25e700bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h684a55ce78393db024e74a42aee558de41e9d8df33ae2ebb253a0290e664d99149573f08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e16ce933bc2d225e89a3e4dff70b7463ab56c711a0250a7f55297cc12532934df1bc95dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff07debf54a05bb83dbcebc9ab29bbd2449f1e9cb8ba6915b083b37b5f991dee5608b849;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10def34d502322f220cd87fce08fa5e1525b6bf2774a4c61874f619cc79ea832e22362ba5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7362f423cae0d3f9a050f18edf453bbe8140b559651991219e2ffc53754dc7eddcdc6325;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d43a568215b71661cb2acb8c3b9c35dd65b87ca6d223dc57c786a18d44e7d0b134be130e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73775f7d7a06e9ab5194ab62aead9dc41736886b32848b799632db594ad29291c1923fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105f30e0877861302cc49a3fab8351c13aac5aaac57477260df8da83a3035a21625275953;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bec9bbae833408ec4ad6a380838042a5cd6a0e27c5cd2ae9eed5a795e8c28dfaf24739e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h608687d80fecf0c9c124210bd1cdf456d12923a7bbf83d6e642850c187e8c6cf81757698;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16996ebef9d4c3c0fd133a02a42f30ac4cd095b47da6a8996d6010d41d4c1afe24510278a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c96132a9d78d9c1e28bac5d5db54f79271f7f2caee6c44e216e640118223d4f29d9f1f86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1934d23e9a0830f1784e2dc037819e86249f6293f52ed8e5b79020498bd9354523fa5422a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b9985b6c4772dffcb4a358ade4db17d4b4964d026375ac4c4c0fc00135b575377a7587d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4c45c76b9215e9ba86988201deeeb629e627132733ac8de0a254f6f3e3feba58ec00be5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18ab155463f1a9fb1ac1870092f534b2fd6099453847e1475a51cbec60d3d4c5f8d831c5f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7979dcc1c43649db5a6967b3bfbc978bcb966c60a0497718017af7d83b90575426764918;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b57b453fbae79d520ecad501a18c0c72e251e7a64c8e49e0e3bfb532ba417b4c3f0a4cc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13380a08dd97d0a911fc0baa7c8c9330032b1fef86b1a834f1f014529b0d51410130d1af4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc846c5737cf4bcefd20cc1cebc9450f49410c5788a9b2ade3ef3c45b4a299b3059fadcf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba05fa6d8859174aefbacd10f3f6da15a4716343865a140eed6e29cd4acb00dc9fdf4e2b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h711ca4a2bfd4f26695a75e92b79e0e8b19f850f18fdc0587ba0ac21786012362bcb77e50;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73d82909464cfc00d8d7c4404a96bf6f0470897498dcc71f130a80976624fa5e62bf65f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13b0e81a03864dc34822d7ee804f3b2cfb31c828bf93f78b42ef0b574696e8dafa8650312;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a40a0e0d7b87f8b3781936b7f03135e2476c72a765fa31c39dbc602440e8e3800d375f0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bb19a467f0d1d44651b2b853e3c06a38de0647c7f2bd7888ac40157f475323d3154af4e8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17716f6b456b82ef1f5cffa36154f4d0e7527632985ddeda501310c72291dbb33e3543afa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca838decb9c9ca735ca8273cce7d339d6f42ac3615152fb21ffa126987175fecd26a0e18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe3cb08aee591368ca3220dfe60851eeb2889d25724dacf83893a64dc7f4d4be5b6909bd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he6452ddb4c102c8129c7d0f7d2fa35523bb979b52e04b16db6a382cd0ffaa9630914afc5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1ef26bce01a257b3fb0e715519264bfabf645fb86a01242f07517356408465b59f0a600;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1242de4a63e690f216792f71d44aa8aaf448e883773f07f11caafc72f0c82a8db8b8f16ae;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3dc600ea1304e7bc6f7b718fb1d552400df64a8334136b0f1b2dd5a18ff335653a8914e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd05de778223a98cc234ee2a7fe8c1c5080617dc480634e891de485d8a03be7762d722ce9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144070ae65d9be8637b78acff10529e1d1f35c15c6dfd410cb1f75107f1c67afa6c6e0340;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d7f21c8a1b3dff05643dfd3fc3ea080f229cd1adcb811bcf87921b674517523fde6e17b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc6fcb9e7f597123e2fc27aa27fab69ddfe28f7b676cea0bce05e1b21acaa5924b17f2ef;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d169989be00a549f06a04558b527a240f7b4d30173c85c206ee973e85a0f4b57663b4e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee436bed58d425becca6ea6c42fb96dd9256dc1d9d05609bb9904c3c140caaabfb11bc24;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c973b8334a8ffc812650f78d25a93b217d402ae43121058c5246337896bbd96029fd999e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30116ae9073e42ced760c9f7d71b4d9d59d8bd2a56c5737f4e244850fd6791fe4bc4b76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153f2f8f4d1a1186a020f5b9869bc0b151cdbcb68a81edf58f2dda6f683d7b2d3b51ad55e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1bbee63e2939fa1563497cac517bf9390a5fbe8253313e99e096efa6422d5934c7d0a17;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14849a88a6ba3d43e6e64d72957d702a6c53ec682871bd9a12e31ec71abef84d66ac12513;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10744345efe1976fbca4560d6fa901ba71087da978d925bb6283e5137c88b61883210419d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcdb13967fe20b7e085e024073b2c02d7e1dd52a08dae3d3c21e523108f89e19614350824;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h119ec4ea56ff7d9bcf8320d8d79f7a3b676eb453c84f387f743eab6ee1748c60f8f19a0b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc49330e726ee5311e99a965fa7893985518cdda7d76e75a58838302bf7efaaedb3a3935b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a90bf7e0705560444f961a51984cf4e984883faa52fe27c86800b89b7a7015b35c55dab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dece13e0f2d7606a5b42638f8c2cf3341bf0d452e17114884cdd5c429f52502f1331546f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1afde2eefc73e0ebf3e87e44114030ab3a60ae18706e5b88955e4ef5eda617f56f1ab939a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e1fc82d874d50ee53c6fb08134a677c45c10d9d7057e3fb1b24ee3443db361b922ec2d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bdb706ecd367600020fb9ebd77ec72b354278c9e86d572d3f9e1dbd64b3c83b683d0d59f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e04fa1f649066ef7c3cdb54614219a6b4a9a1d9d4dd7f4a35c20767329a6c6d10c53f08;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c68316b29ddc66a6fc6f053428d8bf072e730469d61e2afb6c1cd4e2e2bb626ca2735bf6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15de9e38f786f831a279c7d98fb0c8e5b9e747e1ad96c8c0bc4f46efdb1decd364e90594b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4aeff8da264d807426c1c5bafbe12dff86cf7b85f00fccb8efaeba326fb81b289447486c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6fcac8f67cc20bb621fdf78ec2587eba446217a6206fc8e5618719ea5418162330630574;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb51b53b6a95460b2f1dc9db5609aa58f251cf3aca861718810d9e3fce73ccb99c34bf21;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d62069b1c1c1efddc75a0a685134cbe8721ae8906bc5003601c45b75b76881fe4536400;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9a239cc8589ab385408197ff10f0c13831648101f13ff294f627cfebf7433eb2aa17d123;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170cf96f1b72fdf2cd127ee7cad49b89ed9f613b8100456f1cfadaf7907b6bcf16aaf34bc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187d1c44cd70bea85ba97c30d361ea5afaa6786da8670ef88bcb800d9b1cfd6dfe61a0dd8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d79f20a922deef4fc6c10660c62e3db10ce44ca3baea3c90cbc837c3f5a65af3b402506;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10ded01e293218aa21f80a21b7b942b3cb26a551251dffcf647894f925cbb628e4b46d9ac;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h77954da5629a2b45156399301332f26a3a46892289eeddc6c92418216bdd3d56613403a4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h112e1b3317a181716cdd1fefcf9b3a4a41c3f2d711de0c918fe9b64874eec06ae795489d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141d5d4c490a8f332a24adad33ec0e9f85faa13f5451ead67b1351d38d431af6363fc79a0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf86758e9b5b23bf1ef96a4979342647e89a1e017d764b716d075b9b235ccbc87361dd6e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6aab0f1df3dafdf9836f19169d41647680e941d471d782b8005dde297dfa5f610a846e23;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1df35563ee00bdf48d6a1abd6b47448cff81994643c6b20a2440e55677cf3a6d99f3fd520;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7fa1a990a027dd0956a409939289591a21c9f341fbb81bbffd6c501016366d2a1dd4f736;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca10b2a97ec77bfb2a4a3d19300dd0d0548732db9ebbaba94d2637c0c043d5c606332cc3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha53ea71ea7706baccf1133c456edba1b1b19d046303c9e8d1c0593f9db04b40e57fa43f1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66d4eb5a2bdac94d2e7f13f3fac99d63eb003e433a9480aa2032fd460ec6ef47e94a5e9f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e38f36881afe9da2ffe98c0430ceacc2c275868ddc7a8cb3f05534d22cafe645af6b98f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13dc62c8e3016ca64c9275f1922e00456c142d76c9a8018ad14683c2cb2ef78a67acfc69f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ee159429c47a1640855dc06051bb469783619a93887244575b09136f462fe848c61ed91;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ad1dcf969cb4a0b809253e9ca69c204501fb50db65d8053a7d1121f90a48a3d2b8cde8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4bc45838dd8301f24dbd5b029e2d001ea2c49d34133bed83b3436756a4da4446a64bf129;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h887d2e272d38ea856117aa04a7a7bd011286b8a9ca21eaa688b77ad5931f4a030638ff56;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e99f5f97b0e0f68f86d2cc7a93162d412d1a86686f8fd2436f7c6c6db80ae9ff5e067ed1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bb4a7fea4d1bff3c1a0feab351a5da2ded638afdae8666442a978b82c638668ac8bbbd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4853fca7c3aecc0866d8c923eebf642cb0144a0e475bbd85df963229dc37cb82076622f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184fffa89d5f55ce574bde0984bc0659fe86583cf2fe5edcb767cef0746dc2fb5baa74c54;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebe2c7e0038eb5cc7506ac4ac148b490a5b1b2916c4d4113289892750bf863e7513f0e03;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbc3152f0bd16ce6ee7a5ff1369d3af4e32c1a00d81c45e068c9136e4134c50228924fa0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bc03c519dd5d9560089aca51facaa84da8c511df2ee7081c4831db5fe374274003eab7ad;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb6dd0f350c195d1c161e1387582a094fe7a556b61ed200567cbd7fcc70841f00e135fd86;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hffd63413151eb4fd9a8525c9cffacd39078c96f78bea9190a48b2e5f257df48cbde409dd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1823356d8afc7b7652c6929d7ed9cdeb2a4d013ae6ace7ca6329488b85fee929b35d5c63c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9d01569283ef95f8c5bdedaa5231075bfcaed6a0832ed104504b243b38aff9013d27fb4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b2874b111c814f057354e3fe4637ba63136e62097dad223af754f4d7c62bc2a85eae932;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e893c36e81962eb6a93de95234fcfda7b129f9fcc0d1c55e2d09fb5e50ceca1804f6ec5f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6757fd69af97bf4706b2bdb7f75ea178a8c047ec241e01af5e3965182440be985ac59d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h73df214d857a5fe5cdee2fd7b658ba80903f8637375a898c92e5bfd8069bbf08f1a2261a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2c38b13d606f6ada52d11fd75bac0b47c0aef3071c6382182f8a0caa1bd3057b9fc1cbb1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h458c1b5a78dae4d8b3acb77e3f39479f4e858ac6bc30ced631208dabcabaf39273e0dc39;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'heae6f02b1dff3d6a130f81523fb8c53a2d224f3c8e5a6f85480577a7cf5f7d4ef33a2e3d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137c4d7ef0b45dae57ebf83c05ba8c4052302b5807b189c00361fa6842936d62499217755;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18191e9cf76f1cbfd6fb693d2cf6d21cb716dc30a6d02e6716d95965c7d42700aaf5eb973;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b65745c02d2baa3ae697d7deacc1576efcf3b10c4ab6bf301db3809b6f1782c0b6e1321c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f02fabcd6d8729fd889589b41a529837ca608d32a3e1ea18ba797d1d5b8af25539b6ca3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1057010562c67d943d1628234af142a3a76551f0fb9da681cc8de15bac4bd50b7ec7be391;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e0605a7560625ec8ae70f95f487c87de1fc78c3efe40aa02d1e1576518c422cd6c63d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cadb9e7808365f3706368bbadcc166834ed3e1721aab9c9fa08d7ef3fd3f0d94cafebf67;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd4c741f5b5f321d72980061c3b43421bf13a78beb03dc641aa18ac58ea1834cde758cf07;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b132b9ddfba60f6dca64e843ef0d8d7a43551f41c1eea35a2fc1617043a30bd85889cb8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dfb6e9d35f1c39163d9cd79c2c029f5584f5e754ded3cb0aa14eaceaac702fc10d1d4a41;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbcbe733ff469a61834d73d6003de2b317539a570805df38276a7f3eb80ba90661e789d5b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde703e4a485f91b982361bd9c21b23d1ff729f9ea6e956ab6423f1a66cc26417744b34f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7bdf895648cddc0b5604e1a49c8dd73a9fae6a4e88a85a6f6e4f15d211fdd15b1ac14fe7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3175078d94a2f518af7bb7c83372807ce2dda85cf2a54f07fdc87b84a2fb209bd844b2c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30fcb8dd63d36febc3961b35c913f2e0c80b2e769b1d0620193fc739ab1a12d06c7bbb6a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h454b5d5f23985a3c03c4b6fd292c551e6e4ebbe4318b2313744c1afeef5615ff77329baa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b453a7d6e626b02ff754b34356e90bef80217b3d8140da33503ea72895714d1f3730cf71;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbea890af8f68a686ce51e8bb75460c495508b6f5ea44a5c591bc26f4238c507443db855;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1589872656b39cb156d6ce8f34d3273ccad37646a8272d64fa77f1a17e00f039aed671ea7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h163284c6ebe2c96acbbe0d7c9bb6aff381c09711bebad21c366056cbf3d31a699da4e40b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha34ff2f0f4ce90ac60dc2d3e083bca0a249dbf8c63bb48a7e8c557a858edb625e9c08f1e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h633d1eda113bfca67ec8455df367b8639860e0a9861213d0492b303e05c2d42072fb33e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe423c4765a948c0e4c39cf55008aa1ef66f2832faf6248eedc8b79b486dad6d262e1590;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1422b1eecdc72a357914adc6b80942bb2a36b86dfd3f49969f41d159a5f08dedf497d3013;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d0caf366a9626683ce52361a879ae5e31a52dde2a659ce9a8d58592fb12046f996eb6e62;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d57dfd0a3daf4f5c0298a3fd5ab50c60feb86493f3e8d7dbf2227acd6d3d2b277679b98f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd0c50c9b4826d4c0239126a87184aba4475f990c7073c664c0a716cbc2a443229c41c74;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61ad5822816a653a45f7ef6c5629f1a6f14c09a794ccb8ffea448820258ee616b3d7e612;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4571e2a500dbd369ad36d2abe83093dbf4fa88cb263cb82785079dbfde93dc205b5fe1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164b5bc134c896191f4730b28c1ae0fe8ef1fe415f456ab04646ea9591903c9f56bb78d8d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h185a5c526911881cfebecd2b78deb304baa628cdc5949a645fcf7236fcfc5f5455d31aba3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h116c0fdefc1cfcbbc4e779520f4dcc34fe253e29e2fd69296c8dd15515034eeefca039194;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1341a3b423a38a93c47728c25f464150a29263cd02c49e50b9647df65aed6dd895dd35894;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cbbe33d783d94c041fc8e6c30ceb33c50ffef1ebaa8b4befcaf7afa6136ba3091cd86bd2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131bb845a56acf20e1a6bd83ca3bb431d46f9666c9dbf3e55f1711b85239161777eb243d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5453f7b850f72b345591751b0f0b3130086cb487330b223eb480b2b6a12bb1f4665fa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18648e0c8da61d169fac5a572cfc88ed1e55029826aff799435cd3e19cca662e2783b52de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4fd42439ef4312e2be21d08bd076ad726538d81c52c1fa47391c337ba44a038c68d14899;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he197ac9b8db357c8b6a0bf8d14e05a4afbad4bff00c1e88bfb780f4d0be20e693302fc5d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haefcbbf12d753d46a08736108879955022d45442d0e7b038f356da300789aa8ecf6bce0f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3903e341a2eca3ccb81ea9fab8d48e798ee06383a9c033a84d97ead1149fbe1e5d7ed2f9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hae479cc7a819cf0a9e29200468c66ba2c4d4cf88ced9cb644bc5195669fb3792c200bfe0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h88952311938a7c6deffc0b98ebb91e58350661d2bacfe3803b2bbc7710c9203bd1128110;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h129b31745a7bc7b051cbd5e130a01c7ac6c077d1cb5e104975d3e36b0773420f2977a2bc1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b52b886df4da1aa864b07c34ef37a6c380668c2807119a274c71841e9f4a3779c12ec4d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aefdeb30258ed4d6bb73d144ae5039536c29c6a902f20d3d90c000a0c6def759a706d1bb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec4bc4a73accb552414122b1416ebfe55ddbb42da4a423f4c755235da7e68a316eec8d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18250dfa472cae9aa24b8deeeac47f1d7da9917a7dde290e4c6a1e433361d1ea0a43eb549;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7e23b57096a64e867404a6d20aea8fb0cd8b0139d975027fdb2bdb003086b6d0dc6bf6b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3e56f25fadae80f1fcde5a457f7b2095703aa0cb954f6f9b6f6a449a12c6afd13241b82;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d064c6fd79b8dbe766c24edeb709012e191ed4107c44e26b406492eb29139033a71b269;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22f77cc6afc0d463e0ed98731ac7fb40b8a053d60de11c01a9ad8d6f0a986205b03c0d82;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cb5995725f4903db63fa11ec244b79fbb165d8fd246d1d56b2a35ff3e1af4c042392fb76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h189296d7cfb5f888d7477171039c267f893e4985214267681b55e7af42deaf4a1f952f30b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1423fad983e93aa7f5918f0df6afc8dd3118f20a451a7ff413efa1b28f68ddca1719f6bb1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fcd2b4b8e5d6f66ef19922b15ede56d19e82d9523045edfc954fc57b16ba9cf60a6744c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha8e6dc9eac09a848512972db39f7a0b594ed51d2cfc022674017d1915f3fdd74af57e149;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h75ca307f947742302545d719ac42ab24212caf33c5603ca37fd1b521001d2b24043d4c83;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc3aa98f8d7b2d95c47a9f829d976d1cc1706cdc56e4ec9f3713b997fa7686917db524b0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3c10ac043df8848a14daf375ee707c4fb478ec68fc9e50bf6b46c6e6c6635115f3a197e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19914544d4c161b7c5bbcbf5a163b2b234a6225181aaefd2980c6bf94c69d830d4768f187;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h729a12fe5364caa37fd4a992a582542f9b6c9e14ed2941e2c640b4c0875fe02fee30f836;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3978c6fbaf1be39081933bcb00d83c2129b5af95f91323b099851ee3063c51f5a1c5e43f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h170172bcfde9f7ffd4bbbd7b520b911f830d468dee456716bca646120313e82619f5c9f03;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7091cf0fee89c0956ae7637fb1c5acea71babd668e8fbce893278badca481629fb616932;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38e28c821a34762d4c5982b75d68a482d3ea58d652498fe86cbc490dd91970575eb2420e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19753f3e8347551b39fc3953c00b1934f823b0c393fa5dfb4ea7fa05db1d3c0e1236f16e7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he489932290a2f72397260ea7f34406dd12b58430d2798df69467fe745a1137cd180adc76;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0b8edc8cc01da277632c859139780ffb2f9324437c1b561330aa36f7e467df0f282ac31;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha075cdadacbc36e0a71d23bd58ddd4d0a15f2627fe1223e43b5698eb047c30fa0c8f92d5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h91dab9a30564e7f1764e2bfa7ec5c601c1cdb4f7f5379ebd6dd1a8fff82673be4338961a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c14fd751e5ddf6c589f97114366192ff83f6afb12ffa79e7e86909ab5e607db36cd1ef4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8c29c514d5e9c549c8c25ca9558c684ebe7835c80c282d65b21dbe4ffe28496d040705f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h164af67de5d73efa7412e9d151ed06e362c459697e1f182a8aefc86ef009f82188377ac1f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc100e2f27e0ecaa97266531cd14798c566a9703edc82f2f531cad2e7d49d0401d1fee43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1970f9141a792112446e0431f67bd05428401676324d742ee81a64726517112f7e6e670c8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd9898ed9d53c49df8bb63b362dd84ffeb04b33d69c484ebca889e22aa18d33d051db3cb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183f763be65c5d64c060204ab86a8bbdce3ff33518da7add92fcd287e494138643f064183;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h964f11a8d768a9a950e9e9f1ac0deddc01c0fd6fa17ffc712d70e250d05e232f89fb04d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eac5ed2362cf22a2a31f160797d6162dc7ace259162db90857a90c5929e18fc1923b5468;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1891f2889c1d18ade7d0d76910f2497250dc4e4bf5f6e914be7655bd117acb3a068222fe9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd6b945a88fa72dbc8c14eee9aed01310e3c75034f758348878b9faa9e595539120438e2d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f920ca0bdeb68cd3ecd311f67a82736f8520e8b9cb861d5310fea4d58f3eedf471dad78;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c5acdb17ab483e8ae11c83e0979ec52051b4ff4ad41f11ee53624057e3045044f9cedb4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h176d5b61c258dde212977712b7bc13f2a75697176e54dba0721334985b556794d37f25078;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1796912ba84fa5bd8fe97d171b09a0814c831161fee7f36dce742b239dafda8121386c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ffa64cfea798c9002f76a0aa59e69f5b6cff2b456a576f6d8b306e26339794f87ed8dd6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e9c6965a023b88e9257a47fc1e9ebd6253502f1e03603aac5502259cbb477b42a43314a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa214c791851aeb46b595bc8beb81d3a7ba3638259cbaa367bef8f1ed6d11e01e3ac8ba2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18685eaf867ccac5e5b6c447eeb8c6e8cd31793c15e9cc417f51f8790ce8176d70edb775e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e704880a2ad0c5d79bf5f6c87ba700efb9a6046491b9ee9a42832d33d5855d965ee4ea0d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h58077d981218c412f7bcc5e1fb4843fa05f3454e32a8e0b124918bd4cc3a12b4839f2ea6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h39035f7035907bb56ece6ebef35a6b8130072146469357af7f010d1957e8b5872dcafd18;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe8dd2b7e7ab77cbabade278de5c8b5dd3e21e2eed65918ce6f3aa9b330cdfff5a6b44fd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64083134c821a6d896cb7e8adab9c83f001faa2ab3697167936936905b56c81ff0fb82d2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90f4784372d3ba732c0a5cfb68ad8863cc86ea3291d01e43e357701216ef290cb43b6685;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9f9c93ed15c5809793cbd9816d22a4cd22a17ba22354c1def13a5096b70edb39fe740adb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11a425afb7ca129175b64d14befdfd78d957daa21f6b8bd0ddd0eb6f5494be0717d146803;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf9dda24a9c00fc65d8aabb6a437623e0b70e94e0f260f3ff67a42c7eccc3ac2dfe071b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf84f2edb0dbcdbf788840a016468a44935c4751c651f54d8fabac5295f5399211a0423d7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1108f7ab4f6852915ccb8cd4764249e0cf47c002edbff53bb840b81fe19f218bc58298f83;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cbc5892ddc9b808be6ecab3b91833ffc63fa9063d7015fd6fc04feeb22afe02c739635d3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h680f6acf300c66cae06d603bbd7d4a76f25190b0a657453ebe31b4e41b6ef179f973ffbc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94dce6b464134023357aff9afffe9e3ecc39aefe8b69510bc8a51a3840c6d96c5dabb8df;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1457483a613f2a09b55c83e07e53092ae67356ac114bb346ab4b382e7a1de9de001995d2f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1734f711fc11bfab1360edb5a3a518302a77bbce8d1c7932840ffbdf8d90ace4f4edf73a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6a67e07bd3727b8321de9bab673c34607db3db8c67c0d75682f535d33d31069c6d0a038;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b0968d36306e9c100644e37291b79f0e891b18a60d8ee5d8e9319f8c343022e9c59f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f2b5f33d5f5002e672a2050edf76dfc56800e6c0b3ad1d6386b83cc6079b1843d858846;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182c1f0246fd20c00087fac378347b728620f99c03be19d75d75208bda709eb64b80069f7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h690a73986b155e49ee966f89342258bd5f9634f986bdd17bd4ed38d759e3e572e36a38a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18a56a466c6a81d3f337757a45a0295cfc2e1d20b25f9bf0082d7fa3b2230b5aaeeea2de7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f5269bb996adb3baee30f0901b184ef0d318f157439d67b4c7eb1d9c672ba11178f79d8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12df0c7bda5ddfb980dbc162eb60876f3cd2a73cd028cfdcef79d8e4f75dd34fbf0da5a6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15147e8dfead0970e435764a4d241989af8c6d8908ad78fa194103b035298187ebd004325;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14fd88673ecf0f374898329b9271f32af18768d4dbd5df64ecfc5f123ae998aa725d52e09;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fe9767076acda51c05afc5ccc7353f5bbd13ced992ae4c62b068b817d06cd559db2f2428;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1394428a97bd478e104801a887f4211fa0b3cf890eabdeb08ca5664e16313055f08c56dde;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef7a634bba37462b7b40ddd37b90e94b1dcf351b333b28b607142be5352aa8e44af522f3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b3cda23d258872a7da9dae7d62c3f8d973307196666a4945846e6cf9c05dbe158189041;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c649fbe952325fe8e8e75c9305497195466922f0af83153b34a418818c1246dfa11594e0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1130b6aa022bf9678d320ca8fd897a858372f217ba738675ca7957b6769fb7ccc546653f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1118023a1bb6460bc99bb52651c6ec844d4eb5e94d0f3a60b6439242156fc236e9d028f8f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cf231aa416f3a4459a776acd129f3c28548ffcee5e3fd640b22cddb747d1c894a8b5aea0;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd1446a7044abe669d8cb937ccc62e221add5c195f792d705a2540b6ad4b995a44fa791e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15489658b167b459d5c5ecb139f1d3597c28da029b0b90b4ea3f8b7eaace1180cf885af74;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f6de28ef9bf108e034edaf308e7c7b0d9a8a3b78ed2db3dd9c8410c9ec5dc578796e5e5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8d770615d4044a5f22bef0b788bc0f59d883fe8a90aef4e6c7059248f156bbad3f714ced;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72682e80bae21f74c145ba7f669189b5642fb9e6fb98639b8107383f5cebfd1dee11184b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b80c93fe3b2691046bdb54f237e03f9d03081f91d81f647ea2fe4d651f48adb09b9c789f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1feaa058d5f247ec4f609e913ab7247df1f853f637b74d2cece2cf8695ed13719db0451af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h50f97077ac6d5b3c1ed2d4de86c4c0824df754e7a18f1485cc8081adf9dba3e18ee347b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1619c38128a2c05e3583d61ac9741c8ca1c3ba3d890eb2a61fbfd4d53a6723b88a0b02704;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ea87d1a435d0376f6285ca5ed2728b1a6dccd977f9d811ecfcccffed4f915ccc75d5812;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf0447120dfb4e49afe99b3bc85ed8612881edf6ba258561251e7b6af8c5f599f46ea815;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1607da0035b2165849865290aace93ff53db38af048c54b0e841625e460641da99f85d4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135b4c3b27dc6da560a6a9e38dd85a399dc1ed5c7b20c2868ebd61d28e330d1767c886c21;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0fe1db2bc3e5fed51381489d295f8ff97920988273300f14fb0fa989c7a4754b50cfb1a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h232486454820220108c5a7dfe251acbd777a42c98007b8e3eb1c02181dbb8745de3a48f8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7bc0a651c9353a29d701fcbe56b34ca0010c374ffd23ab629cbb6b8031bc2bdae5d2b885;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h165149b7cb641f1db3b8b08c80428bc60667e8a0fd961d58483eae601e4bacf0daf2a9e2e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111a6c054a29ff546de40c4cb6ccfe0888b63e26bb95ea920b1e3b3149ddeac193e0a0747;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a88ee2f52ecdd6ebeae8e6e881b828c5028b723264de5bcfb75e972f417f5afb245643a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37aa812570ab37b34025e18556ebe08b3cb9ff6e3253b5ada0b4a719d31796f5f83d0483;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa7d12080e3e8f6f32f49b9a6db274dcaab6dab67ac4729686c1299b8be73ef069b077b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b14a6b5092e5370f210fcc0a10a8037b69aadd487cd3f3007510abb762d8dca27340b63c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h205c6fa25189955b69adde7a81a7a14e692abe25c0335fbe70a1b8b9110d0a9b1abbe90e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1101857b22d03ab68f449bd21a5a4526d5d34229412e78dd97e0a2e0fa06a3c44470d2f89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h382f52ff8d6c75980ceb4cb8a6c9c0c8e34437a958b4b44ba721d40990a492f50b02fdfb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc9cd8fdc8be09b7954e0811e1ed0c10792b2d87c16a41f71a601ba656bf0399f9a9e042;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12da40285d2d9dbedafc521f6bb33362cb0bb479e207885390fe7cde011a2b6f25bd76d67;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4fc463236337be4ab246a5a5ac83ae9d95c84b402c8bdfeb56322edb29747e760cfad4f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f8f78981299f5b8d709468b060fba91c2f2b405489674cd7e758ed5cf922f53ed216891;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1063871083d1ea0c4f0cfc42cce0d4ffa112bdfe81d92206ecc2ec55e3a8921512949c78d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd199c907aeef9ee2f298e194f0d56ba137a40d1b8bb895cd24301f3021b86672ab42829;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h20306307e4a3b1405d7a52d5f98fdaa4c827fc36917a66c00cc666e19bf8b6062c673965;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c994dfe18c6824f57a27b37ca2c6732f2a8deb721f436fec5474d3907f84ea76fbcc6e1;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e7813c007a46d870f23cbbf9ca031ed4a5c69595b0e91fe4d89698e9c8493e5838773a8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d6358e92e72008d28ad15e8271e8a5eda2196b0644303a67606811e78024cfbf1eb4c6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72902d92541f7211f1567574e0bb2055360e395c9e2fe152ee2d0ddce43ed2089f9fd9c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h157e198288b0b71a326b2fa64db712ed725a0cbfde8832859a308fc0fe5541ee02dcae66b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a1dc9276d928fccf9267b797a16d68de644d8c72dd02675e19c5c22d9a4a6d5d6aa0fde;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19090a7a70a99a45c905b6c0f08787d2d235725d91ac94800dfd0a8a215f2a4f9ef0b8694;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5c3a76d15cc8eee8186774335c2995bb2f61c379c83d54118d0bd7be58f606b184490a9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cbd3048ed687ebbbf754e0b8f5ca3b225d929e07c1ee5ca383f896d1855f74154998a21d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9349fd9d449096faa3837afc6a7bc3a4aff21de4e708a918a42cbf8205b552bff21d633c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h41167c233b68a43e502e73b8e75bdb7dfec9cfcbd0370abc72bd326190186ed623d6fe0d;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c391c48898840e4c749c9210bdde7837e994241c294a64ec7960094f6595b391b7e3a02;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1579acf73e2df77f2a6bfc86680f7775db776a60a1960716e2fec28ad351fe2e21833bb3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f7237aa2fb085779e09cccc549c0c768fc3dcadec43d9208f26767157011adebe31e81a7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf19a37f7c2ef5235cbc26d41f259fa8a09100cfdf6bf6545bbb1f4fa403e1669384a5a82;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107fd3ca49ed395ceb87f4348b5510c5e7381e26eebaa2aeed7c48e0f6676f846ddff6bf9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16cbbf3f1679c52b1f12e314341433c3ef0aa2895ba843dcacced5a727072e43137a7ea43;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c57c8c9387ffb7d546efb1ea2725229591769ec9aeb9c81e9e18f459dc08267041c85b1b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd94c0f27d858ec90a424d027054e2ccd97e91e4a942ca2fe414c4ae8945f11af3ca7ebd;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc80a7d307f6ff96bb3528b0b26b33dc5c20be3c1d73f51ed3eebed7ca23aa11e172819c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72af85e1c38cd733fb446efe0a9c7aef11b9de92a8f5960c9058025a72a851cf6b2ee4b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha407a1d88913555d76b9ee1ffd2ca32dd56ebd5a4ba898a006a7866197b55cf10ec70578;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1970625ecb2c7644563040dae5d70bab92236a72b046d8f76c79cb22fbfc3c67849f8ebd9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h193ea07d1eac694add1b3d3112670c5fe29b0a1f3631cd5892e7c0693ada3a40c0394c061;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hacb09eff4fdd02e2de59f70f65a8dff8ed42172c8fb5b2e5b436a47ba8d74963dcc1423e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6746c69c07ec7f6349691519a5d32926c9900d10be6c7fd8841a92bb6b0c85e6d418617;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115390371cad52d69bf2046813bf9deb1befbb88b23eb4372599ca11721587a1eb0083af;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h560302887ca56929717cce9553028a36c30db829631ad090a0614de17eb0bd46c6e8c3d6;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f414a6e8f62feccc8b9b21899aea2bfb5679343304227455cd4f5f32694d859309015de;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he3b7ed6aff987b134ab3cd5ccee70d6ef62cc5b151f986a68f3478ce30f4c6bfd07a85d9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15eae7e0df24f5cceacdf42a24b20171402ca39196862bb4a9fff9a094645eeb3ed662b40;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd29fb50e52c937303a5c9f9c394fedbd4d8ba71693dd0da35d895c6e75bf4d19ba6e539b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d1aa2094964028c043f7f5b279aa028d8a3c2dd1af8af5e02fc563f7f751136ea68c676;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14d867c5c740330383baf9b592490fbbfc671f51b0a95da2e8978a549d33820e1725e36b5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ebe977e0de0c03b439d674d0affe0e36b42891491f0d4187fc1aab9203d60a7320f47b9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5791a7d43e3a6adc9f3103f6ea05912453e482ea772d8df26426df47bf6cc407bced557;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c985076d35a49c98373452be50e92bc4fedfc28c192dff581d7dffa4f0ccc555b93267;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a36f1302810ad9e45dac8c3faea99b744c7ea7819485643f9295ea8b8510587d89d9ba03;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h101990f37f8e1460eb1c9b7ef1bc2c7abb69c50c1a2e28b250d008c51810f152dc2f2545;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14539aeb186763779f93e459fc8647be16dbc2048e01f9f22878b32d8f9c150356fa7a9b3;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1425ea12634777781c74e4457a9899196027c61ab4fdeec251c7cec0d6fcce0bc78df2d2c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7189af6c44b7c4e0b45009cf0e59b73f51bd857ef7f7bb3779bda5fcb1f8c7f43303f12a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c9883dd82480bf8abcfed6800189b84ce2ed4c2d0a1fb41959ef61de443b36b0e86a40f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed7488e9c6b1287356ed8b52d9e4b0630ae25338a013b882852a2a5e0abcddef277afc9;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182f3948e02bce0c8bc4540419c174086d3ad382e722c3e2cff9266af1ead6c73e1fa4528;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hacbdec012db29e668922cabca3abe13031213018b8c0fcfef39d192e59219ae1ed1f00ea;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cc37dc9eb76d1c1bfadcfdca6fa57cdaee1a494b5944069be29f54fa4f9d3f4a78d0f69;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4bd2857a6cc4cbf3254f2ba7eb182f284a9635eae278dda07ba227e5bdd669ef591491a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38e9b21bbd289941f2ea23a102b2de4e3e8799d27be527db4290acef857783098e177fd2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h171a395825a7e6bee8a0d9021ed21cb86dfb581d433064af943040f187fc63d958e72d02e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e7cda2bf2bfc0ba700f482c9461174e5595fee9fb241ce24d1504c6cdb433de3c2b11bc5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h816fd2412fa4c760037c3d4c851529cb8e96eaa960d43d7e43aa37d01713c4debc04a855;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ba3f31ac61f84427a16a074abf2afa4b58ba6fee090d781865afe10355ed9a5bc3c11c2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15401c9a35c763fbe45fd1feb65312cfcf476995bc0a56e4c48abbe41c9cc967282ac5660;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5cec7dbc66caf83825963baf74dd57cad28d694d4dc55c436f870d09fa15fa3b7176476;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11cc48797cfe704470a81b64627915b091ebde4567162793bc798f264bf4eb448605ef119;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2ca5b0388804f89da026c78f6c3719748ca6de1703a544452ab4410b9c91ef867c07237c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19636db2dbd748c22e7c541021046455796af06e0e2351b7f642b83f3e7804c705ce06791;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff955dad1a448857a82c54858ca17302adbb1cc904646a699929cacad4f885bb884c73fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d9853f932a603ee735ac46f677a9e0aabbf20586830b06816d3d0590b1f4bfe24f7576e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17083717051eadceba3863fba8a88ebab9dae9aadac33e9d383d9da61133c7972d64cc8ab;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d07a11396b38c881a5fb6fa65b6f20b041da6b05fbcf4401ab2561b04f8ce6e0352bb3dc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hedf63ddbed231996d40317860ed71886b5416a37743a5bcadb9f60d8cd654a7968874667;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13abf53835ddbb9ff895a3bfe7221afb8d61cc1962fb4584ae8fe76029f9a5e4f90122bdc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd069a3aad5f9308c35177a87a0a8bef1beb20dcbdab3eea1198d9e2bf56ff6c87dc8967;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c78584ce31f906c98c5e0877202ec35a29678a0aaba10f543d693158200e1bf66db47213;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17762bafc073621746a533f6f991e111ba48771ab9896785bac5f7d961443dd0ad379f946;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3fd840e57293d42b312c425e73412465749f04f059e17a51b82c24e03fe3127114b127f;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64d0f6160d8d333e633b26e00ed9f15e82887559aa6dea96179756f89d15295121006b39;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1a47cef1e280345067f2d19af7011468e7a0efbb13852aa6186b2fb3e82ebc46f4147fc;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc49b45e37f981e6c5a1b1c081e2f2a884a1fb40f0f0ef339141559bf03fb5d3f66ba81b8;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0693101ea1809726c4826e40c8ad7e255e7213313c7bf6207e80e51166e2bf08483842e;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h118c47ee12d6bd30fca09e05a8fa4f0a4a580234221d46773ba0a2dedda9f90bf41ee01fe;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a794df632f067cf6333d50a89aae85aa82063e316882b1191780a1e515840f00b7d910;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2569570650dfd7dba85c10abc0ee2999794117de5c1fda2fb44dd35e892c2e92bd92f014;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h148a4a70af980131ed0d98529d9472e8a56b3b173a32a031bb5cc0fe83d91ac4e2ac23ec;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183843e93cc98215b57944d66f6d23fb7a6fddb9fb2a52a595f45a245f85112afa8a86fdb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd84597f5e28fc746024c2455a152432774cb8c8669331fed30fed67c920572e806767f94;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h163a4a3db37d7fac43336b96faca1c9fa2e5773522deaaa6e7c198c6bde0c966774868a47;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h270effb45b324333a674b388e230f0f41f61647be8d89c200181664fdfc511a48af8def7;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114abb59fd1f68e33f3ee1cd391510d9515c3f8b213a6344b9a0f9b32d95e4dc4b1eddc89;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h79818875c80430e634951bae39f48c4517eb9e64cbd8ecd77e795cb65a02b3fd8908e33b;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a9736bff2326a42af41d2355aac99a8d35f0992c52143c019c142743884deb4efd087eaa;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9781926dd846c97b36f371c1ddd94fb5d4b4564b7ddda1e425e6eedfaa63b08196fcbf2;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62c52140d439f282dfe419fee5e3269ff4f9698e4be3fd70264edbdfa419e31cf606db1c;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1825b13d02770bfe98fe61ea8acb763f7450352ffab5219af407d6bf5c8ab2467adf8746a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd3457a1baa9178c1ac0b152279ed4426e2dc9ed0ba7a14b77c73904eb0ba4514dcb37bf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16edb4190160273a4150eda8767cda748c731cddb923ac878e13d66b24325a08fdd12b222;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h741c0649c8726618da5d60dc61181d27a7038ee7c03764f763f072468d963160eb085e25;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4bc51a88f9fb9b310b00f444c620d21e2c530d3f3616dec35c0f74e3173ed6bb3f38fbeb;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h139900496420d0808f4326d284989576d8132c3d40a7d2154aa560438fc746c1b5f70ae00;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h191bd587a9d49a8976da441a55c5ee21a940a03e3569551772b64fc5cb6656b23d5223388;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h72da98ec3c36903e74331ea0dc473a90aa3edb5639fa2ec47d4d5bc96bca5873e841ed0a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1679e18b4cfa865eee889194ba39f7864d9319442a803ca37820f9d629a08fff20b803ff4;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2cc4bf16614814c64b3f2c43e498191107d0d840a6fc175588bf953ac7846e933f1279f5;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e96c9be2730cf2d94b6fda2d4a105abacfc82f6bf1fe2ecb59aec4fdd472e551262e4f4a;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1715f2170d2704a3f8ff8b712d51d7aae683dd7e0b5dfc137dedd7c8fa2a384d772bba287;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b64173d46e4b95bc8193cf94951bda4d790882f078203ded62990efe3b5274686159a9cf;
        #1
        {src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b1417d4329ac394dc1239d1af176a434445bc4608584d0ec5674029c06182c4a2d2d5f5;
        #1
        $finish();
    end
endmodule
