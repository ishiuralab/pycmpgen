// probclass: mul
// size:      15
// stage:     12
// cost:      28
// elapsed:   7204.863266468048
module compressor (
      input wire [0:0] src0,
      input wire [1:0] src1,
      input wire [2:0] src2,
      input wire [3:0] src3,
      input wire [4:0] src4,
      input wire [5:0] src5,
      input wire [6:0] src6,
      input wire [7:0] src7,
      input wire [8:0] src8,
      input wire [9:0] src9,
      input wire [10:0] src10,
      input wire [11:0] src11,
      input wire [12:0] src12,
      input wire [13:0] src13,
      input wire [14:0] src14,
      input wire [13:0] src15,
      input wire [12:0] src16,
      input wire [11:0] src17,
      input wire [10:0] src18,
      input wire [9:0] src19,
      input wire [8:0] src20,
      input wire [7:0] src21,
      input wire [6:0] src22,
      input wire [5:0] src23,
      input wire [4:0] src24,
      input wire [3:0] src25,
      input wire [2:0] src26,
      input wire [1:0] src27,
      input wire [0:0] src28,
      output wire [0:0] dst0,
      output wire [0:0] dst1,
      output wire [0:0] dst2,
      output wire [0:0] dst3,
      output wire [0:0] dst4,
      output wire [0:0] dst5,
      output wire [0:0] dst6,
      output wire [0:0] dst7,
      output wire [0:0] dst8,
      output wire [0:0] dst9,
      output wire [0:0] dst10,
      output wire [0:0] dst11,
      output wire [0:0] dst12,
      output wire [0:0] dst13,
      output wire [0:0] dst14,
      output wire [0:0] dst15,
      output wire [0:0] dst16,
      output wire [0:0] dst17,
      output wire [0:0] dst18,
      output wire [0:0] dst19,
      output wire [0:0] dst20,
      output wire [0:0] dst21,
      output wire [0:0] dst22,
      output wire [0:0] dst23,
      output wire [0:0] dst24,
      output wire [0:0] dst25,
      output wire [0:0] dst26,
      output wire [0:0] dst27,
      output wire [0:0] dst28,
      output wire [0:0] dst29);

   wire [0:0] stage0_0;
   wire [1:0] stage0_1;
   wire [2:0] stage0_2;
   wire [3:0] stage0_3;
   wire [4:0] stage0_4;
   wire [5:0] stage0_5;
   wire [6:0] stage0_6;
   wire [7:0] stage0_7;
   wire [8:0] stage0_8;
   wire [9:0] stage0_9;
   wire [10:0] stage0_10;
   wire [11:0] stage0_11;
   wire [12:0] stage0_12;
   wire [13:0] stage0_13;
   wire [14:0] stage0_14;
   wire [13:0] stage0_15;
   wire [12:0] stage0_16;
   wire [11:0] stage0_17;
   wire [10:0] stage0_18;
   wire [9:0] stage0_19;
   wire [8:0] stage0_20;
   wire [7:0] stage0_21;
   wire [6:0] stage0_22;
   wire [5:0] stage0_23;
   wire [4:0] stage0_24;
   wire [3:0] stage0_25;
   wire [2:0] stage0_26;
   wire [1:0] stage0_27;
   wire [0:0] stage0_28;
   wire [0:0] stage1_0;
   wire [0:0] stage1_1;
   wire [0:0] stage1_2;
   wire [0:0] stage1_3;
   wire [5:0] stage1_4;
   wire [6:0] stage1_5;
   wire [6:0] stage1_6;
   wire [7:0] stage1_7;
   wire [8:0] stage1_8;
   wire [3:0] stage1_9;
   wire [11:0] stage1_10;
   wire [6:0] stage1_11;
   wire [13:0] stage1_12;
   wire [14:0] stage1_13;
   wire [14:0] stage1_14;
   wire [13:0] stage1_15;
   wire [12:0] stage1_16;
   wire [11:0] stage1_17;
   wire [10:0] stage1_18;
   wire [3:0] stage1_19;
   wire [3:0] stage1_20;
   wire [3:0] stage1_21;
   wire [2:0] stage1_22;
   wire [7:0] stage1_23;
   wire [5:0] stage1_24;
   wire [3:0] stage1_25;
   wire [2:0] stage1_26;
   wire [1:0] stage1_27;
   wire [0:0] stage1_28;
   wire [0:0] stage2_0;
   wire [0:0] stage2_1;
   wire [0:0] stage2_2;
   wire [0:0] stage2_3;
   wire [5:0] stage2_4;
   wire [0:0] stage2_5;
   wire [1:0] stage2_6;
   wire [3:0] stage2_7;
   wire [6:0] stage2_8;
   wire [4:0] stage2_9;
   wire [6:0] stage2_10;
   wire [4:0] stage2_11;
   wire [5:0] stage2_12;
   wire [8:0] stage2_13;
   wire [4:0] stage2_14;
   wire [5:0] stage2_15;
   wire [4:0] stage2_16;
   wire [9:0] stage2_17;
   wire [13:0] stage2_18;
   wire [4:0] stage2_19;
   wire [3:0] stage2_20;
   wire [3:0] stage2_21;
   wire [2:0] stage2_22;
   wire [7:0] stage2_23;
   wire [5:0] stage2_24;
   wire [3:0] stage2_25;
   wire [2:0] stage2_26;
   wire [1:0] stage2_27;
   wire [0:0] stage2_28;
   wire [0:0] stage3_0;
   wire [0:0] stage3_1;
   wire [0:0] stage3_2;
   wire [0:0] stage3_3;
   wire [0:0] stage3_4;
   wire [0:0] stage3_5;
   wire [0:0] stage3_6;
   wire [3:0] stage3_7;
   wire [1:0] stage3_8;
   wire [5:0] stage3_9;
   wire [1:0] stage3_10;
   wire [1:0] stage3_11;
   wire [6:0] stage3_12;
   wire [3:0] stage3_13;
   wire [5:0] stage3_14;
   wire [1:0] stage3_15;
   wire [5:0] stage3_16;
   wire [4:0] stage3_17;
   wire [14:0] stage3_18;
   wire [5:0] stage3_19;
   wire [3:0] stage3_20;
   wire [3:0] stage3_21;
   wire [2:0] stage3_22;
   wire [7:0] stage3_23;
   wire [5:0] stage3_24;
   wire [3:0] stage3_25;
   wire [2:0] stage3_26;
   wire [1:0] stage3_27;
   wire [0:0] stage3_28;
   wire [0:0] stage4_0;
   wire [0:0] stage4_1;
   wire [0:0] stage4_2;
   wire [0:0] stage4_3;
   wire [0:0] stage4_4;
   wire [0:0] stage4_5;
   wire [0:0] stage4_6;
   wire [0:0] stage4_7;
   wire [0:0] stage4_8;
   wire [2:0] stage4_9;
   wire [2:0] stage4_10;
   wire [2:0] stage4_11;
   wire [0:0] stage4_12;
   wire [4:0] stage4_13;
   wire [0:0] stage4_14;
   wire [2:0] stage4_15;
   wire [6:0] stage4_16;
   wire [4:0] stage4_17;
   wire [14:0] stage4_18;
   wire [5:0] stage4_19;
   wire [3:0] stage4_20;
   wire [3:0] stage4_21;
   wire [2:0] stage4_22;
   wire [7:0] stage4_23;
   wire [5:0] stage4_24;
   wire [3:0] stage4_25;
   wire [2:0] stage4_26;
   wire [1:0] stage4_27;
   wire [0:0] stage4_28;
   wire [0:0] stage5_0;
   wire [0:0] stage5_1;
   wire [0:0] stage5_2;
   wire [0:0] stage5_3;
   wire [0:0] stage5_4;
   wire [0:0] stage5_5;
   wire [0:0] stage5_6;
   wire [0:0] stage5_7;
   wire [0:0] stage5_8;
   wire [0:0] stage5_9;
   wire [0:0] stage5_10;
   wire [0:0] stage5_11;
   wire [0:0] stage5_12;
   wire [5:0] stage5_13;
   wire [0:0] stage5_14;
   wire [2:0] stage5_15;
   wire [0:0] stage5_16;
   wire [1:0] stage5_17;
   wire [9:0] stage5_18;
   wire [1:0] stage5_19;
   wire [5:0] stage5_20;
   wire [4:0] stage5_21;
   wire [2:0] stage5_22;
   wire [7:0] stage5_23;
   wire [5:0] stage5_24;
   wire [3:0] stage5_25;
   wire [2:0] stage5_26;
   wire [1:0] stage5_27;
   wire [0:0] stage5_28;
   wire [0:0] stage6_0;
   wire [0:0] stage6_1;
   wire [0:0] stage6_2;
   wire [0:0] stage6_3;
   wire [0:0] stage6_4;
   wire [0:0] stage6_5;
   wire [0:0] stage6_6;
   wire [0:0] stage6_7;
   wire [0:0] stage6_8;
   wire [0:0] stage6_9;
   wire [0:0] stage6_10;
   wire [0:0] stage6_11;
   wire [0:0] stage6_12;
   wire [0:0] stage6_13;
   wire [0:0] stage6_14;
   wire [0:0] stage6_15;
   wire [0:0] stage6_16;
   wire [2:0] stage6_17;
   wire [3:0] stage6_18;
   wire [2:0] stage6_19;
   wire [0:0] stage6_20;
   wire [5:0] stage6_21;
   wire [3:0] stage6_22;
   wire [7:0] stage6_23;
   wire [5:0] stage6_24;
   wire [3:0] stage6_25;
   wire [2:0] stage6_26;
   wire [1:0] stage6_27;
   wire [0:0] stage6_28;
   wire [0:0] stage7_0;
   wire [0:0] stage7_1;
   wire [0:0] stage7_2;
   wire [0:0] stage7_3;
   wire [0:0] stage7_4;
   wire [0:0] stage7_5;
   wire [0:0] stage7_6;
   wire [0:0] stage7_7;
   wire [0:0] stage7_8;
   wire [0:0] stage7_9;
   wire [0:0] stage7_10;
   wire [0:0] stage7_11;
   wire [0:0] stage7_12;
   wire [0:0] stage7_13;
   wire [0:0] stage7_14;
   wire [0:0] stage7_15;
   wire [0:0] stage7_16;
   wire [0:0] stage7_17;
   wire [0:0] stage7_18;
   wire [0:0] stage7_19;
   wire [0:0] stage7_20;
   wire [6:0] stage7_21;
   wire [3:0] stage7_22;
   wire [7:0] stage7_23;
   wire [5:0] stage7_24;
   wire [3:0] stage7_25;
   wire [2:0] stage7_26;
   wire [1:0] stage7_27;
   wire [0:0] stage7_28;
   wire [0:0] stage8_0;
   wire [0:0] stage8_1;
   wire [0:0] stage8_2;
   wire [0:0] stage8_3;
   wire [0:0] stage8_4;
   wire [0:0] stage8_5;
   wire [0:0] stage8_6;
   wire [0:0] stage8_7;
   wire [0:0] stage8_8;
   wire [0:0] stage8_9;
   wire [0:0] stage8_10;
   wire [0:0] stage8_11;
   wire [0:0] stage8_12;
   wire [0:0] stage8_13;
   wire [0:0] stage8_14;
   wire [0:0] stage8_15;
   wire [0:0] stage8_16;
   wire [0:0] stage8_17;
   wire [0:0] stage8_18;
   wire [0:0] stage8_19;
   wire [0:0] stage8_20;
   wire [6:0] stage8_21;
   wire [3:0] stage8_22;
   wire [7:0] stage8_23;
   wire [5:0] stage8_24;
   wire [3:0] stage8_25;
   wire [2:0] stage8_26;
   wire [1:0] stage8_27;
   wire [0:0] stage8_28;
   wire [0:0] stage9_0;
   wire [0:0] stage9_1;
   wire [0:0] stage9_2;
   wire [0:0] stage9_3;
   wire [0:0] stage9_4;
   wire [0:0] stage9_5;
   wire [0:0] stage9_6;
   wire [0:0] stage9_7;
   wire [0:0] stage9_8;
   wire [0:0] stage9_9;
   wire [0:0] stage9_10;
   wire [0:0] stage9_11;
   wire [0:0] stage9_12;
   wire [0:0] stage9_13;
   wire [0:0] stage9_14;
   wire [0:0] stage9_15;
   wire [0:0] stage9_16;
   wire [0:0] stage9_17;
   wire [0:0] stage9_18;
   wire [0:0] stage9_19;
   wire [0:0] stage9_20;
   wire [0:0] stage9_21;
   wire [4:0] stage9_22;
   wire [2:0] stage9_23;
   wire [6:0] stage9_24;
   wire [4:0] stage9_25;
   wire [2:0] stage9_26;
   wire [1:0] stage9_27;
   wire [0:0] stage9_28;
   wire [0:0] stage10_0;
   wire [0:0] stage10_1;
   wire [0:0] stage10_2;
   wire [0:0] stage10_3;
   wire [0:0] stage10_4;
   wire [0:0] stage10_5;
   wire [0:0] stage10_6;
   wire [0:0] stage10_7;
   wire [0:0] stage10_8;
   wire [0:0] stage10_9;
   wire [0:0] stage10_10;
   wire [0:0] stage10_11;
   wire [0:0] stage10_12;
   wire [0:0] stage10_13;
   wire [0:0] stage10_14;
   wire [0:0] stage10_15;
   wire [0:0] stage10_16;
   wire [0:0] stage10_17;
   wire [0:0] stage10_18;
   wire [0:0] stage10_19;
   wire [0:0] stage10_20;
   wire [0:0] stage10_21;
   wire [0:0] stage10_22;
   wire [2:0] stage10_23;
   wire [1:0] stage10_24;
   wire [5:0] stage10_25;
   wire [3:0] stage10_26;
   wire [1:0] stage10_27;
   wire [0:0] stage10_28;
   wire [0:0] stage11_0;
   wire [0:0] stage11_1;
   wire [0:0] stage11_2;
   wire [0:0] stage11_3;
   wire [0:0] stage11_4;
   wire [0:0] stage11_5;
   wire [0:0] stage11_6;
   wire [0:0] stage11_7;
   wire [0:0] stage11_8;
   wire [0:0] stage11_9;
   wire [0:0] stage11_10;
   wire [0:0] stage11_11;
   wire [0:0] stage11_12;
   wire [0:0] stage11_13;
   wire [0:0] stage11_14;
   wire [0:0] stage11_15;
   wire [0:0] stage11_16;
   wire [0:0] stage11_17;
   wire [0:0] stage11_18;
   wire [0:0] stage11_19;
   wire [0:0] stage11_20;
   wire [0:0] stage11_21;
   wire [0:0] stage11_22;
   wire [0:0] stage11_23;
   wire [0:0] stage11_24;
   wire [0:0] stage11_25;
   wire [4:0] stage11_26;
   wire [2:0] stage11_27;
   wire [0:0] stage11_28;
   wire [0:0] stage12_0;
   wire [0:0] stage12_1;
   wire [0:0] stage12_2;
   wire [0:0] stage12_3;
   wire [0:0] stage12_4;
   wire [0:0] stage12_5;
   wire [0:0] stage12_6;
   wire [0:0] stage12_7;
   wire [0:0] stage12_8;
   wire [0:0] stage12_9;
   wire [0:0] stage12_10;
   wire [0:0] stage12_11;
   wire [0:0] stage12_12;
   wire [0:0] stage12_13;
   wire [0:0] stage12_14;
   wire [0:0] stage12_15;
   wire [0:0] stage12_16;
   wire [0:0] stage12_17;
   wire [0:0] stage12_18;
   wire [0:0] stage12_19;
   wire [0:0] stage12_20;
   wire [0:0] stage12_21;
   wire [0:0] stage12_22;
   wire [0:0] stage12_23;
   wire [0:0] stage12_24;
   wire [0:0] stage12_25;
   wire [0:0] stage12_26;
   wire [0:0] stage12_27;
   wire [0:0] stage12_28;
   wire [0:0] stage12_29;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign dst0 = stage12_0;
   assign dst1 = stage12_1;
   assign dst2 = stage12_2;
   assign dst3 = stage12_3;
   assign dst4 = stage12_4;
   assign dst5 = stage12_5;
   assign dst6 = stage12_6;
   assign dst7 = stage12_7;
   assign dst8 = stage12_8;
   assign dst9 = stage12_9;
   assign dst10 = stage12_10;
   assign dst11 = stage12_11;
   assign dst12 = stage12_12;
   assign dst13 = stage12_13;
   assign dst14 = stage12_14;
   assign dst15 = stage12_15;
   assign dst16 = stage12_16;
   assign dst17 = stage12_17;
   assign dst18 = stage12_18;
   assign dst19 = stage12_19;
   assign dst20 = stage12_20;
   assign dst21 = stage12_21;
   assign dst22 = stage12_22;
   assign dst23 = stage12_23;
   assign dst24 = stage12_24;
   assign dst25 = stage12_25;
   assign dst26 = stage12_26;
   assign dst27 = stage12_27;
   assign dst28 = stage12_28;
   assign dst29 = stage12_29;

   gpc433_5 gpc0 (
      {stage0_1[0], stage0_1[1], 1'b0},
      {stage0_2[0], stage0_2[1], stage0_2[2]},
      {stage0_3[0], stage0_3[1], stage0_3[2], stage0_3[3]},
      {stage1_5[0],stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0]}
   );
   gpc607_5 gpc1 (
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5], stage0_9[6]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[0],stage1_11[0],stage1_10[0],stage1_9[0]}
   );
   gpc607_5 gpc2 (
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5], stage0_19[6]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[0],stage1_21[0],stage1_20[0],stage1_19[0]}
   );
   gpc607_5 gpc3 (
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5], stage0_20[6]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[1],stage1_22[1],stage1_21[1],stage1_20[1]}
   );
   gpc1_1 gpc4 (
      {stage0_0[0]},
      {stage1_0[0]}
   );
   gpc1_1 gpc5 (
      {stage0_4[0]},
      {stage1_4[1]}
   );
   gpc1_1 gpc6 (
      {stage0_4[1]},
      {stage1_4[2]}
   );
   gpc1_1 gpc7 (
      {stage0_4[2]},
      {stage1_4[3]}
   );
   gpc1_1 gpc8 (
      {stage0_4[3]},
      {stage1_4[4]}
   );
   gpc1_1 gpc9 (
      {stage0_4[4]},
      {stage1_4[5]}
   );
   gpc1_1 gpc10 (
      {stage0_5[0]},
      {stage1_5[1]}
   );
   gpc1_1 gpc11 (
      {stage0_5[1]},
      {stage1_5[2]}
   );
   gpc1_1 gpc12 (
      {stage0_5[2]},
      {stage1_5[3]}
   );
   gpc1_1 gpc13 (
      {stage0_5[3]},
      {stage1_5[4]}
   );
   gpc1_1 gpc14 (
      {stage0_5[4]},
      {stage1_5[5]}
   );
   gpc1_1 gpc15 (
      {stage0_5[5]},
      {stage1_5[6]}
   );
   gpc1_1 gpc16 (
      {stage0_6[0]},
      {stage1_6[0]}
   );
   gpc1_1 gpc17 (
      {stage0_6[1]},
      {stage1_6[1]}
   );
   gpc1_1 gpc18 (
      {stage0_6[2]},
      {stage1_6[2]}
   );
   gpc1_1 gpc19 (
      {stage0_6[3]},
      {stage1_6[3]}
   );
   gpc1_1 gpc20 (
      {stage0_6[4]},
      {stage1_6[4]}
   );
   gpc1_1 gpc21 (
      {stage0_6[5]},
      {stage1_6[5]}
   );
   gpc1_1 gpc22 (
      {stage0_6[6]},
      {stage1_6[6]}
   );
   gpc1_1 gpc23 (
      {stage0_7[0]},
      {stage1_7[0]}
   );
   gpc1_1 gpc24 (
      {stage0_7[1]},
      {stage1_7[1]}
   );
   gpc1_1 gpc25 (
      {stage0_7[2]},
      {stage1_7[2]}
   );
   gpc1_1 gpc26 (
      {stage0_7[3]},
      {stage1_7[3]}
   );
   gpc1_1 gpc27 (
      {stage0_7[4]},
      {stage1_7[4]}
   );
   gpc1_1 gpc28 (
      {stage0_7[5]},
      {stage1_7[5]}
   );
   gpc1_1 gpc29 (
      {stage0_7[6]},
      {stage1_7[6]}
   );
   gpc1_1 gpc30 (
      {stage0_7[7]},
      {stage1_7[7]}
   );
   gpc1_1 gpc31 (
      {stage0_8[0]},
      {stage1_8[0]}
   );
   gpc1_1 gpc32 (
      {stage0_8[1]},
      {stage1_8[1]}
   );
   gpc1_1 gpc33 (
      {stage0_8[2]},
      {stage1_8[2]}
   );
   gpc1_1 gpc34 (
      {stage0_8[3]},
      {stage1_8[3]}
   );
   gpc1_1 gpc35 (
      {stage0_8[4]},
      {stage1_8[4]}
   );
   gpc1_1 gpc36 (
      {stage0_8[5]},
      {stage1_8[5]}
   );
   gpc1_1 gpc37 (
      {stage0_8[6]},
      {stage1_8[6]}
   );
   gpc1_1 gpc38 (
      {stage0_8[7]},
      {stage1_8[7]}
   );
   gpc1_1 gpc39 (
      {stage0_8[8]},
      {stage1_8[8]}
   );
   gpc1_1 gpc40 (
      {stage0_9[7]},
      {stage1_9[1]}
   );
   gpc1_1 gpc41 (
      {stage0_9[8]},
      {stage1_9[2]}
   );
   gpc1_1 gpc42 (
      {stage0_9[9]},
      {stage1_9[3]}
   );
   gpc1_1 gpc43 (
      {stage0_10[0]},
      {stage1_10[1]}
   );
   gpc1_1 gpc44 (
      {stage0_10[1]},
      {stage1_10[2]}
   );
   gpc1_1 gpc45 (
      {stage0_10[2]},
      {stage1_10[3]}
   );
   gpc1_1 gpc46 (
      {stage0_10[3]},
      {stage1_10[4]}
   );
   gpc1_1 gpc47 (
      {stage0_10[4]},
      {stage1_10[5]}
   );
   gpc1_1 gpc48 (
      {stage0_10[5]},
      {stage1_10[6]}
   );
   gpc1_1 gpc49 (
      {stage0_10[6]},
      {stage1_10[7]}
   );
   gpc1_1 gpc50 (
      {stage0_10[7]},
      {stage1_10[8]}
   );
   gpc1_1 gpc51 (
      {stage0_10[8]},
      {stage1_10[9]}
   );
   gpc1_1 gpc52 (
      {stage0_10[9]},
      {stage1_10[10]}
   );
   gpc1_1 gpc53 (
      {stage0_10[10]},
      {stage1_10[11]}
   );
   gpc1_1 gpc54 (
      {stage0_11[6]},
      {stage1_11[1]}
   );
   gpc1_1 gpc55 (
      {stage0_11[7]},
      {stage1_11[2]}
   );
   gpc1_1 gpc56 (
      {stage0_11[8]},
      {stage1_11[3]}
   );
   gpc1_1 gpc57 (
      {stage0_11[9]},
      {stage1_11[4]}
   );
   gpc1_1 gpc58 (
      {stage0_11[10]},
      {stage1_11[5]}
   );
   gpc1_1 gpc59 (
      {stage0_11[11]},
      {stage1_11[6]}
   );
   gpc1_1 gpc60 (
      {stage0_12[0]},
      {stage1_12[1]}
   );
   gpc1_1 gpc61 (
      {stage0_12[1]},
      {stage1_12[2]}
   );
   gpc1_1 gpc62 (
      {stage0_12[2]},
      {stage1_12[3]}
   );
   gpc1_1 gpc63 (
      {stage0_12[3]},
      {stage1_12[4]}
   );
   gpc1_1 gpc64 (
      {stage0_12[4]},
      {stage1_12[5]}
   );
   gpc1_1 gpc65 (
      {stage0_12[5]},
      {stage1_12[6]}
   );
   gpc1_1 gpc66 (
      {stage0_12[6]},
      {stage1_12[7]}
   );
   gpc1_1 gpc67 (
      {stage0_12[7]},
      {stage1_12[8]}
   );
   gpc1_1 gpc68 (
      {stage0_12[8]},
      {stage1_12[9]}
   );
   gpc1_1 gpc69 (
      {stage0_12[9]},
      {stage1_12[10]}
   );
   gpc1_1 gpc70 (
      {stage0_12[10]},
      {stage1_12[11]}
   );
   gpc1_1 gpc71 (
      {stage0_12[11]},
      {stage1_12[12]}
   );
   gpc1_1 gpc72 (
      {stage0_12[12]},
      {stage1_12[13]}
   );
   gpc1_1 gpc73 (
      {stage0_13[0]},
      {stage1_13[1]}
   );
   gpc1_1 gpc74 (
      {stage0_13[1]},
      {stage1_13[2]}
   );
   gpc1_1 gpc75 (
      {stage0_13[2]},
      {stage1_13[3]}
   );
   gpc1_1 gpc76 (
      {stage0_13[3]},
      {stage1_13[4]}
   );
   gpc1_1 gpc77 (
      {stage0_13[4]},
      {stage1_13[5]}
   );
   gpc1_1 gpc78 (
      {stage0_13[5]},
      {stage1_13[6]}
   );
   gpc1_1 gpc79 (
      {stage0_13[6]},
      {stage1_13[7]}
   );
   gpc1_1 gpc80 (
      {stage0_13[7]},
      {stage1_13[8]}
   );
   gpc1_1 gpc81 (
      {stage0_13[8]},
      {stage1_13[9]}
   );
   gpc1_1 gpc82 (
      {stage0_13[9]},
      {stage1_13[10]}
   );
   gpc1_1 gpc83 (
      {stage0_13[10]},
      {stage1_13[11]}
   );
   gpc1_1 gpc84 (
      {stage0_13[11]},
      {stage1_13[12]}
   );
   gpc1_1 gpc85 (
      {stage0_13[12]},
      {stage1_13[13]}
   );
   gpc1_1 gpc86 (
      {stage0_13[13]},
      {stage1_13[14]}
   );
   gpc1_1 gpc87 (
      {stage0_14[0]},
      {stage1_14[0]}
   );
   gpc1_1 gpc88 (
      {stage0_14[1]},
      {stage1_14[1]}
   );
   gpc1_1 gpc89 (
      {stage0_14[2]},
      {stage1_14[2]}
   );
   gpc1_1 gpc90 (
      {stage0_14[3]},
      {stage1_14[3]}
   );
   gpc1_1 gpc91 (
      {stage0_14[4]},
      {stage1_14[4]}
   );
   gpc1_1 gpc92 (
      {stage0_14[5]},
      {stage1_14[5]}
   );
   gpc1_1 gpc93 (
      {stage0_14[6]},
      {stage1_14[6]}
   );
   gpc1_1 gpc94 (
      {stage0_14[7]},
      {stage1_14[7]}
   );
   gpc1_1 gpc95 (
      {stage0_14[8]},
      {stage1_14[8]}
   );
   gpc1_1 gpc96 (
      {stage0_14[9]},
      {stage1_14[9]}
   );
   gpc1_1 gpc97 (
      {stage0_14[10]},
      {stage1_14[10]}
   );
   gpc1_1 gpc98 (
      {stage0_14[11]},
      {stage1_14[11]}
   );
   gpc1_1 gpc99 (
      {stage0_14[12]},
      {stage1_14[12]}
   );
   gpc1_1 gpc100 (
      {stage0_14[13]},
      {stage1_14[13]}
   );
   gpc1_1 gpc101 (
      {stage0_14[14]},
      {stage1_14[14]}
   );
   gpc1_1 gpc102 (
      {stage0_15[0]},
      {stage1_15[0]}
   );
   gpc1_1 gpc103 (
      {stage0_15[1]},
      {stage1_15[1]}
   );
   gpc1_1 gpc104 (
      {stage0_15[2]},
      {stage1_15[2]}
   );
   gpc1_1 gpc105 (
      {stage0_15[3]},
      {stage1_15[3]}
   );
   gpc1_1 gpc106 (
      {stage0_15[4]},
      {stage1_15[4]}
   );
   gpc1_1 gpc107 (
      {stage0_15[5]},
      {stage1_15[5]}
   );
   gpc1_1 gpc108 (
      {stage0_15[6]},
      {stage1_15[6]}
   );
   gpc1_1 gpc109 (
      {stage0_15[7]},
      {stage1_15[7]}
   );
   gpc1_1 gpc110 (
      {stage0_15[8]},
      {stage1_15[8]}
   );
   gpc1_1 gpc111 (
      {stage0_15[9]},
      {stage1_15[9]}
   );
   gpc1_1 gpc112 (
      {stage0_15[10]},
      {stage1_15[10]}
   );
   gpc1_1 gpc113 (
      {stage0_15[11]},
      {stage1_15[11]}
   );
   gpc1_1 gpc114 (
      {stage0_15[12]},
      {stage1_15[12]}
   );
   gpc1_1 gpc115 (
      {stage0_15[13]},
      {stage1_15[13]}
   );
   gpc1_1 gpc116 (
      {stage0_16[0]},
      {stage1_16[0]}
   );
   gpc1_1 gpc117 (
      {stage0_16[1]},
      {stage1_16[1]}
   );
   gpc1_1 gpc118 (
      {stage0_16[2]},
      {stage1_16[2]}
   );
   gpc1_1 gpc119 (
      {stage0_16[3]},
      {stage1_16[3]}
   );
   gpc1_1 gpc120 (
      {stage0_16[4]},
      {stage1_16[4]}
   );
   gpc1_1 gpc121 (
      {stage0_16[5]},
      {stage1_16[5]}
   );
   gpc1_1 gpc122 (
      {stage0_16[6]},
      {stage1_16[6]}
   );
   gpc1_1 gpc123 (
      {stage0_16[7]},
      {stage1_16[7]}
   );
   gpc1_1 gpc124 (
      {stage0_16[8]},
      {stage1_16[8]}
   );
   gpc1_1 gpc125 (
      {stage0_16[9]},
      {stage1_16[9]}
   );
   gpc1_1 gpc126 (
      {stage0_16[10]},
      {stage1_16[10]}
   );
   gpc1_1 gpc127 (
      {stage0_16[11]},
      {stage1_16[11]}
   );
   gpc1_1 gpc128 (
      {stage0_16[12]},
      {stage1_16[12]}
   );
   gpc1_1 gpc129 (
      {stage0_17[0]},
      {stage1_17[0]}
   );
   gpc1_1 gpc130 (
      {stage0_17[1]},
      {stage1_17[1]}
   );
   gpc1_1 gpc131 (
      {stage0_17[2]},
      {stage1_17[2]}
   );
   gpc1_1 gpc132 (
      {stage0_17[3]},
      {stage1_17[3]}
   );
   gpc1_1 gpc133 (
      {stage0_17[4]},
      {stage1_17[4]}
   );
   gpc1_1 gpc134 (
      {stage0_17[5]},
      {stage1_17[5]}
   );
   gpc1_1 gpc135 (
      {stage0_17[6]},
      {stage1_17[6]}
   );
   gpc1_1 gpc136 (
      {stage0_17[7]},
      {stage1_17[7]}
   );
   gpc1_1 gpc137 (
      {stage0_17[8]},
      {stage1_17[8]}
   );
   gpc1_1 gpc138 (
      {stage0_17[9]},
      {stage1_17[9]}
   );
   gpc1_1 gpc139 (
      {stage0_17[10]},
      {stage1_17[10]}
   );
   gpc1_1 gpc140 (
      {stage0_17[11]},
      {stage1_17[11]}
   );
   gpc1_1 gpc141 (
      {stage0_18[0]},
      {stage1_18[0]}
   );
   gpc1_1 gpc142 (
      {stage0_18[1]},
      {stage1_18[1]}
   );
   gpc1_1 gpc143 (
      {stage0_18[2]},
      {stage1_18[2]}
   );
   gpc1_1 gpc144 (
      {stage0_18[3]},
      {stage1_18[3]}
   );
   gpc1_1 gpc145 (
      {stage0_18[4]},
      {stage1_18[4]}
   );
   gpc1_1 gpc146 (
      {stage0_18[5]},
      {stage1_18[5]}
   );
   gpc1_1 gpc147 (
      {stage0_18[6]},
      {stage1_18[6]}
   );
   gpc1_1 gpc148 (
      {stage0_18[7]},
      {stage1_18[7]}
   );
   gpc1_1 gpc149 (
      {stage0_18[8]},
      {stage1_18[8]}
   );
   gpc1_1 gpc150 (
      {stage0_18[9]},
      {stage1_18[9]}
   );
   gpc1_1 gpc151 (
      {stage0_18[10]},
      {stage1_18[10]}
   );
   gpc1_1 gpc152 (
      {stage0_19[7]},
      {stage1_19[1]}
   );
   gpc1_1 gpc153 (
      {stage0_19[8]},
      {stage1_19[2]}
   );
   gpc1_1 gpc154 (
      {stage0_19[9]},
      {stage1_19[3]}
   );
   gpc1_1 gpc155 (
      {stage0_20[7]},
      {stage1_20[2]}
   );
   gpc1_1 gpc156 (
      {stage0_20[8]},
      {stage1_20[3]}
   );
   gpc1_1 gpc157 (
      {stage0_21[6]},
      {stage1_21[2]}
   );
   gpc1_1 gpc158 (
      {stage0_21[7]},
      {stage1_21[3]}
   );
   gpc1_1 gpc159 (
      {stage0_22[6]},
      {stage1_22[2]}
   );
   gpc1_1 gpc160 (
      {stage0_23[0]},
      {stage1_23[2]}
   );
   gpc1_1 gpc161 (
      {stage0_23[1]},
      {stage1_23[3]}
   );
   gpc1_1 gpc162 (
      {stage0_23[2]},
      {stage1_23[4]}
   );
   gpc1_1 gpc163 (
      {stage0_23[3]},
      {stage1_23[5]}
   );
   gpc1_1 gpc164 (
      {stage0_23[4]},
      {stage1_23[6]}
   );
   gpc1_1 gpc165 (
      {stage0_23[5]},
      {stage1_23[7]}
   );
   gpc1_1 gpc166 (
      {stage0_24[0]},
      {stage1_24[1]}
   );
   gpc1_1 gpc167 (
      {stage0_24[1]},
      {stage1_24[2]}
   );
   gpc1_1 gpc168 (
      {stage0_24[2]},
      {stage1_24[3]}
   );
   gpc1_1 gpc169 (
      {stage0_24[3]},
      {stage1_24[4]}
   );
   gpc1_1 gpc170 (
      {stage0_24[4]},
      {stage1_24[5]}
   );
   gpc1_1 gpc171 (
      {stage0_25[0]},
      {stage1_25[0]}
   );
   gpc1_1 gpc172 (
      {stage0_25[1]},
      {stage1_25[1]}
   );
   gpc1_1 gpc173 (
      {stage0_25[2]},
      {stage1_25[2]}
   );
   gpc1_1 gpc174 (
      {stage0_25[3]},
      {stage1_25[3]}
   );
   gpc1_1 gpc175 (
      {stage0_26[0]},
      {stage1_26[0]}
   );
   gpc1_1 gpc176 (
      {stage0_26[1]},
      {stage1_26[1]}
   );
   gpc1_1 gpc177 (
      {stage0_26[2]},
      {stage1_26[2]}
   );
   gpc1_1 gpc178 (
      {stage0_27[0]},
      {stage1_27[0]}
   );
   gpc1_1 gpc179 (
      {stage0_27[1]},
      {stage1_27[1]}
   );
   gpc1_1 gpc180 (
      {stage0_28[0]},
      {stage1_28[0]}
   );
   gpc607_5 gpc181 (
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5], stage1_5[6]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[0],stage2_7[0],stage2_6[0],stage2_5[0]}
   );
   gpc1407_5 gpc182 (
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3]},
      {stage1_9[0]},
      {stage2_10[0],stage2_9[1],stage2_8[1],stage2_7[1],stage2_6[1]}
   );
   gpc607_5 gpc183 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5], stage1_10[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[0],stage2_11[0],stage2_10[1]}
   );
   gpc1244_5 gpc184 (
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9]},
      {stage1_13[0], stage1_13[1]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[1],stage2_12[1],stage2_11[1]}
   );
   gpc607_5 gpc185 (
      {stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7], stage1_13[8]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[1],stage2_14[2],stage2_13[2]}
   );
   gpc607_5 gpc186 (
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[1],stage2_16[1],stage2_15[2],stage2_14[3]}
   );
   gpc607_5 gpc187 (
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12], stage1_14[13], stage1_14[14]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[2],stage2_16[2],stage2_15[3],stage2_14[4]}
   );
   gpc607_5 gpc188 (
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11], stage1_15[12]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[2],stage2_17[3],stage2_16[3],stage2_15[4]}
   );
   gpc1_1 gpc189 (
      {stage1_0[0]},
      {stage2_0[0]}
   );
   gpc1_1 gpc190 (
      {stage1_1[0]},
      {stage2_1[0]}
   );
   gpc1_1 gpc191 (
      {stage1_2[0]},
      {stage2_2[0]}
   );
   gpc1_1 gpc192 (
      {stage1_3[0]},
      {stage2_3[0]}
   );
   gpc1_1 gpc193 (
      {stage1_4[0]},
      {stage2_4[0]}
   );
   gpc1_1 gpc194 (
      {stage1_4[1]},
      {stage2_4[1]}
   );
   gpc1_1 gpc195 (
      {stage1_4[2]},
      {stage2_4[2]}
   );
   gpc1_1 gpc196 (
      {stage1_4[3]},
      {stage2_4[3]}
   );
   gpc1_1 gpc197 (
      {stage1_4[4]},
      {stage2_4[4]}
   );
   gpc1_1 gpc198 (
      {stage1_4[5]},
      {stage2_4[5]}
   );
   gpc1_1 gpc199 (
      {stage1_7[6]},
      {stage2_7[2]}
   );
   gpc1_1 gpc200 (
      {stage1_7[7]},
      {stage2_7[3]}
   );
   gpc1_1 gpc201 (
      {stage1_8[4]},
      {stage2_8[2]}
   );
   gpc1_1 gpc202 (
      {stage1_8[5]},
      {stage2_8[3]}
   );
   gpc1_1 gpc203 (
      {stage1_8[6]},
      {stage2_8[4]}
   );
   gpc1_1 gpc204 (
      {stage1_8[7]},
      {stage2_8[5]}
   );
   gpc1_1 gpc205 (
      {stage1_8[8]},
      {stage2_8[6]}
   );
   gpc1_1 gpc206 (
      {stage1_9[1]},
      {stage2_9[2]}
   );
   gpc1_1 gpc207 (
      {stage1_9[2]},
      {stage2_9[3]}
   );
   gpc1_1 gpc208 (
      {stage1_9[3]},
      {stage2_9[4]}
   );
   gpc1_1 gpc209 (
      {stage1_10[7]},
      {stage2_10[2]}
   );
   gpc1_1 gpc210 (
      {stage1_10[8]},
      {stage2_10[3]}
   );
   gpc1_1 gpc211 (
      {stage1_10[9]},
      {stage2_10[4]}
   );
   gpc1_1 gpc212 (
      {stage1_10[10]},
      {stage2_10[5]}
   );
   gpc1_1 gpc213 (
      {stage1_10[11]},
      {stage2_10[6]}
   );
   gpc1_1 gpc214 (
      {stage1_11[4]},
      {stage2_11[2]}
   );
   gpc1_1 gpc215 (
      {stage1_11[5]},
      {stage2_11[3]}
   );
   gpc1_1 gpc216 (
      {stage1_11[6]},
      {stage2_11[4]}
   );
   gpc1_1 gpc217 (
      {stage1_12[10]},
      {stage2_12[2]}
   );
   gpc1_1 gpc218 (
      {stage1_12[11]},
      {stage2_12[3]}
   );
   gpc1_1 gpc219 (
      {stage1_12[12]},
      {stage2_12[4]}
   );
   gpc1_1 gpc220 (
      {stage1_12[13]},
      {stage2_12[5]}
   );
   gpc1_1 gpc221 (
      {stage1_13[9]},
      {stage2_13[3]}
   );
   gpc1_1 gpc222 (
      {stage1_13[10]},
      {stage2_13[4]}
   );
   gpc1_1 gpc223 (
      {stage1_13[11]},
      {stage2_13[5]}
   );
   gpc1_1 gpc224 (
      {stage1_13[12]},
      {stage2_13[6]}
   );
   gpc1_1 gpc225 (
      {stage1_13[13]},
      {stage2_13[7]}
   );
   gpc1_1 gpc226 (
      {stage1_13[14]},
      {stage2_13[8]}
   );
   gpc1_1 gpc227 (
      {stage1_15[13]},
      {stage2_15[5]}
   );
   gpc1_1 gpc228 (
      {stage1_16[12]},
      {stage2_16[4]}
   );
   gpc1_1 gpc229 (
      {stage1_17[6]},
      {stage2_17[4]}
   );
   gpc1_1 gpc230 (
      {stage1_17[7]},
      {stage2_17[5]}
   );
   gpc1_1 gpc231 (
      {stage1_17[8]},
      {stage2_17[6]}
   );
   gpc1_1 gpc232 (
      {stage1_17[9]},
      {stage2_17[7]}
   );
   gpc1_1 gpc233 (
      {stage1_17[10]},
      {stage2_17[8]}
   );
   gpc1_1 gpc234 (
      {stage1_17[11]},
      {stage2_17[9]}
   );
   gpc1_1 gpc235 (
      {stage1_18[0]},
      {stage2_18[3]}
   );
   gpc1_1 gpc236 (
      {stage1_18[1]},
      {stage2_18[4]}
   );
   gpc1_1 gpc237 (
      {stage1_18[2]},
      {stage2_18[5]}
   );
   gpc1_1 gpc238 (
      {stage1_18[3]},
      {stage2_18[6]}
   );
   gpc1_1 gpc239 (
      {stage1_18[4]},
      {stage2_18[7]}
   );
   gpc1_1 gpc240 (
      {stage1_18[5]},
      {stage2_18[8]}
   );
   gpc1_1 gpc241 (
      {stage1_18[6]},
      {stage2_18[9]}
   );
   gpc1_1 gpc242 (
      {stage1_18[7]},
      {stage2_18[10]}
   );
   gpc1_1 gpc243 (
      {stage1_18[8]},
      {stage2_18[11]}
   );
   gpc1_1 gpc244 (
      {stage1_18[9]},
      {stage2_18[12]}
   );
   gpc1_1 gpc245 (
      {stage1_18[10]},
      {stage2_18[13]}
   );
   gpc1_1 gpc246 (
      {stage1_19[0]},
      {stage2_19[1]}
   );
   gpc1_1 gpc247 (
      {stage1_19[1]},
      {stage2_19[2]}
   );
   gpc1_1 gpc248 (
      {stage1_19[2]},
      {stage2_19[3]}
   );
   gpc1_1 gpc249 (
      {stage1_19[3]},
      {stage2_19[4]}
   );
   gpc1_1 gpc250 (
      {stage1_20[0]},
      {stage2_20[0]}
   );
   gpc1_1 gpc251 (
      {stage1_20[1]},
      {stage2_20[1]}
   );
   gpc1_1 gpc252 (
      {stage1_20[2]},
      {stage2_20[2]}
   );
   gpc1_1 gpc253 (
      {stage1_20[3]},
      {stage2_20[3]}
   );
   gpc1_1 gpc254 (
      {stage1_21[0]},
      {stage2_21[0]}
   );
   gpc1_1 gpc255 (
      {stage1_21[1]},
      {stage2_21[1]}
   );
   gpc1_1 gpc256 (
      {stage1_21[2]},
      {stage2_21[2]}
   );
   gpc1_1 gpc257 (
      {stage1_21[3]},
      {stage2_21[3]}
   );
   gpc1_1 gpc258 (
      {stage1_22[0]},
      {stage2_22[0]}
   );
   gpc1_1 gpc259 (
      {stage1_22[1]},
      {stage2_22[1]}
   );
   gpc1_1 gpc260 (
      {stage1_22[2]},
      {stage2_22[2]}
   );
   gpc1_1 gpc261 (
      {stage1_23[0]},
      {stage2_23[0]}
   );
   gpc1_1 gpc262 (
      {stage1_23[1]},
      {stage2_23[1]}
   );
   gpc1_1 gpc263 (
      {stage1_23[2]},
      {stage2_23[2]}
   );
   gpc1_1 gpc264 (
      {stage1_23[3]},
      {stage2_23[3]}
   );
   gpc1_1 gpc265 (
      {stage1_23[4]},
      {stage2_23[4]}
   );
   gpc1_1 gpc266 (
      {stage1_23[5]},
      {stage2_23[5]}
   );
   gpc1_1 gpc267 (
      {stage1_23[6]},
      {stage2_23[6]}
   );
   gpc1_1 gpc268 (
      {stage1_23[7]},
      {stage2_23[7]}
   );
   gpc1_1 gpc269 (
      {stage1_24[0]},
      {stage2_24[0]}
   );
   gpc1_1 gpc270 (
      {stage1_24[1]},
      {stage2_24[1]}
   );
   gpc1_1 gpc271 (
      {stage1_24[2]},
      {stage2_24[2]}
   );
   gpc1_1 gpc272 (
      {stage1_24[3]},
      {stage2_24[3]}
   );
   gpc1_1 gpc273 (
      {stage1_24[4]},
      {stage2_24[4]}
   );
   gpc1_1 gpc274 (
      {stage1_24[5]},
      {stage2_24[5]}
   );
   gpc1_1 gpc275 (
      {stage1_25[0]},
      {stage2_25[0]}
   );
   gpc1_1 gpc276 (
      {stage1_25[1]},
      {stage2_25[1]}
   );
   gpc1_1 gpc277 (
      {stage1_25[2]},
      {stage2_25[2]}
   );
   gpc1_1 gpc278 (
      {stage1_25[3]},
      {stage2_25[3]}
   );
   gpc1_1 gpc279 (
      {stage1_26[0]},
      {stage2_26[0]}
   );
   gpc1_1 gpc280 (
      {stage1_26[1]},
      {stage2_26[1]}
   );
   gpc1_1 gpc281 (
      {stage1_26[2]},
      {stage2_26[2]}
   );
   gpc1_1 gpc282 (
      {stage1_27[0]},
      {stage2_27[0]}
   );
   gpc1_1 gpc283 (
      {stage1_27[1]},
      {stage2_27[1]}
   );
   gpc1_1 gpc284 (
      {stage1_28[0]},
      {stage2_28[0]}
   );
   gpc1316_5 gpc285 (
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage2_5[0]},
      {stage2_6[0], stage2_6[1], 1'b0},
      {stage2_7[0]},
      {stage3_8[0],stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[0]}
   );
   gpc607_5 gpc286 (
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[0],stage3_8[1]}
   );
   gpc615_5 gpc287 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[0]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[1],stage3_11[1]}
   );
   gpc607_5 gpc288 (
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], 1'b0},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[0],stage3_17[0],stage3_16[0],stage3_15[1]}
   );
   gpc1_1 gpc289 (
      {stage2_0[0]},
      {stage3_0[0]}
   );
   gpc1_1 gpc290 (
      {stage2_1[0]},
      {stage3_1[0]}
   );
   gpc1_1 gpc291 (
      {stage2_2[0]},
      {stage3_2[0]}
   );
   gpc1_1 gpc292 (
      {stage2_3[0]},
      {stage3_3[0]}
   );
   gpc1_1 gpc293 (
      {stage2_7[1]},
      {stage3_7[1]}
   );
   gpc1_1 gpc294 (
      {stage2_7[2]},
      {stage3_7[2]}
   );
   gpc1_1 gpc295 (
      {stage2_7[3]},
      {stage3_7[3]}
   );
   gpc1_1 gpc296 (
      {stage2_9[0]},
      {stage3_9[1]}
   );
   gpc1_1 gpc297 (
      {stage2_9[1]},
      {stage3_9[2]}
   );
   gpc1_1 gpc298 (
      {stage2_9[2]},
      {stage3_9[3]}
   );
   gpc1_1 gpc299 (
      {stage2_9[3]},
      {stage3_9[4]}
   );
   gpc1_1 gpc300 (
      {stage2_9[4]},
      {stage3_9[5]}
   );
   gpc1_1 gpc301 (
      {stage2_10[6]},
      {stage3_10[1]}
   );
   gpc1_1 gpc302 (
      {stage2_12[1]},
      {stage3_12[2]}
   );
   gpc1_1 gpc303 (
      {stage2_12[2]},
      {stage3_12[3]}
   );
   gpc1_1 gpc304 (
      {stage2_12[3]},
      {stage3_12[4]}
   );
   gpc1_1 gpc305 (
      {stage2_12[4]},
      {stage3_12[5]}
   );
   gpc1_1 gpc306 (
      {stage2_12[5]},
      {stage3_12[6]}
   );
   gpc1_1 gpc307 (
      {stage2_13[6]},
      {stage3_13[1]}
   );
   gpc1_1 gpc308 (
      {stage2_13[7]},
      {stage3_13[2]}
   );
   gpc1_1 gpc309 (
      {stage2_13[8]},
      {stage3_13[3]}
   );
   gpc1_1 gpc310 (
      {stage2_14[0]},
      {stage3_14[1]}
   );
   gpc1_1 gpc311 (
      {stage2_14[1]},
      {stage3_14[2]}
   );
   gpc1_1 gpc312 (
      {stage2_14[2]},
      {stage3_14[3]}
   );
   gpc1_1 gpc313 (
      {stage2_14[3]},
      {stage3_14[4]}
   );
   gpc1_1 gpc314 (
      {stage2_14[4]},
      {stage3_14[5]}
   );
   gpc1_1 gpc315 (
      {stage2_16[0]},
      {stage3_16[1]}
   );
   gpc1_1 gpc316 (
      {stage2_16[1]},
      {stage3_16[2]}
   );
   gpc1_1 gpc317 (
      {stage2_16[2]},
      {stage3_16[3]}
   );
   gpc1_1 gpc318 (
      {stage2_16[3]},
      {stage3_16[4]}
   );
   gpc1_1 gpc319 (
      {stage2_16[4]},
      {stage3_16[5]}
   );
   gpc1_1 gpc320 (
      {stage2_17[6]},
      {stage3_17[1]}
   );
   gpc1_1 gpc321 (
      {stage2_17[7]},
      {stage3_17[2]}
   );
   gpc1_1 gpc322 (
      {stage2_17[8]},
      {stage3_17[3]}
   );
   gpc1_1 gpc323 (
      {stage2_17[9]},
      {stage3_17[4]}
   );
   gpc1_1 gpc324 (
      {stage2_18[0]},
      {stage3_18[1]}
   );
   gpc1_1 gpc325 (
      {stage2_18[1]},
      {stage3_18[2]}
   );
   gpc1_1 gpc326 (
      {stage2_18[2]},
      {stage3_18[3]}
   );
   gpc1_1 gpc327 (
      {stage2_18[3]},
      {stage3_18[4]}
   );
   gpc1_1 gpc328 (
      {stage2_18[4]},
      {stage3_18[5]}
   );
   gpc1_1 gpc329 (
      {stage2_18[5]},
      {stage3_18[6]}
   );
   gpc1_1 gpc330 (
      {stage2_18[6]},
      {stage3_18[7]}
   );
   gpc1_1 gpc331 (
      {stage2_18[7]},
      {stage3_18[8]}
   );
   gpc1_1 gpc332 (
      {stage2_18[8]},
      {stage3_18[9]}
   );
   gpc1_1 gpc333 (
      {stage2_18[9]},
      {stage3_18[10]}
   );
   gpc1_1 gpc334 (
      {stage2_18[10]},
      {stage3_18[11]}
   );
   gpc1_1 gpc335 (
      {stage2_18[11]},
      {stage3_18[12]}
   );
   gpc1_1 gpc336 (
      {stage2_18[12]},
      {stage3_18[13]}
   );
   gpc1_1 gpc337 (
      {stage2_18[13]},
      {stage3_18[14]}
   );
   gpc1_1 gpc338 (
      {stage2_19[0]},
      {stage3_19[1]}
   );
   gpc1_1 gpc339 (
      {stage2_19[1]},
      {stage3_19[2]}
   );
   gpc1_1 gpc340 (
      {stage2_19[2]},
      {stage3_19[3]}
   );
   gpc1_1 gpc341 (
      {stage2_19[3]},
      {stage3_19[4]}
   );
   gpc1_1 gpc342 (
      {stage2_19[4]},
      {stage3_19[5]}
   );
   gpc1_1 gpc343 (
      {stage2_20[0]},
      {stage3_20[0]}
   );
   gpc1_1 gpc344 (
      {stage2_20[1]},
      {stage3_20[1]}
   );
   gpc1_1 gpc345 (
      {stage2_20[2]},
      {stage3_20[2]}
   );
   gpc1_1 gpc346 (
      {stage2_20[3]},
      {stage3_20[3]}
   );
   gpc1_1 gpc347 (
      {stage2_21[0]},
      {stage3_21[0]}
   );
   gpc1_1 gpc348 (
      {stage2_21[1]},
      {stage3_21[1]}
   );
   gpc1_1 gpc349 (
      {stage2_21[2]},
      {stage3_21[2]}
   );
   gpc1_1 gpc350 (
      {stage2_21[3]},
      {stage3_21[3]}
   );
   gpc1_1 gpc351 (
      {stage2_22[0]},
      {stage3_22[0]}
   );
   gpc1_1 gpc352 (
      {stage2_22[1]},
      {stage3_22[1]}
   );
   gpc1_1 gpc353 (
      {stage2_22[2]},
      {stage3_22[2]}
   );
   gpc1_1 gpc354 (
      {stage2_23[0]},
      {stage3_23[0]}
   );
   gpc1_1 gpc355 (
      {stage2_23[1]},
      {stage3_23[1]}
   );
   gpc1_1 gpc356 (
      {stage2_23[2]},
      {stage3_23[2]}
   );
   gpc1_1 gpc357 (
      {stage2_23[3]},
      {stage3_23[3]}
   );
   gpc1_1 gpc358 (
      {stage2_23[4]},
      {stage3_23[4]}
   );
   gpc1_1 gpc359 (
      {stage2_23[5]},
      {stage3_23[5]}
   );
   gpc1_1 gpc360 (
      {stage2_23[6]},
      {stage3_23[6]}
   );
   gpc1_1 gpc361 (
      {stage2_23[7]},
      {stage3_23[7]}
   );
   gpc1_1 gpc362 (
      {stage2_24[0]},
      {stage3_24[0]}
   );
   gpc1_1 gpc363 (
      {stage2_24[1]},
      {stage3_24[1]}
   );
   gpc1_1 gpc364 (
      {stage2_24[2]},
      {stage3_24[2]}
   );
   gpc1_1 gpc365 (
      {stage2_24[3]},
      {stage3_24[3]}
   );
   gpc1_1 gpc366 (
      {stage2_24[4]},
      {stage3_24[4]}
   );
   gpc1_1 gpc367 (
      {stage2_24[5]},
      {stage3_24[5]}
   );
   gpc1_1 gpc368 (
      {stage2_25[0]},
      {stage3_25[0]}
   );
   gpc1_1 gpc369 (
      {stage2_25[1]},
      {stage3_25[1]}
   );
   gpc1_1 gpc370 (
      {stage2_25[2]},
      {stage3_25[2]}
   );
   gpc1_1 gpc371 (
      {stage2_25[3]},
      {stage3_25[3]}
   );
   gpc1_1 gpc372 (
      {stage2_26[0]},
      {stage3_26[0]}
   );
   gpc1_1 gpc373 (
      {stage2_26[1]},
      {stage3_26[1]}
   );
   gpc1_1 gpc374 (
      {stage2_26[2]},
      {stage3_26[2]}
   );
   gpc1_1 gpc375 (
      {stage2_27[0]},
      {stage3_27[0]}
   );
   gpc1_1 gpc376 (
      {stage2_27[1]},
      {stage3_27[1]}
   );
   gpc1_1 gpc377 (
      {stage2_28[0]},
      {stage3_28[0]}
   );
   gpc425_5 gpc378 (
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], 1'b0},
      {stage3_8[0], stage3_8[1]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3]},
      {stage4_11[0],stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[0]}
   );
   gpc607_5 gpc379 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[0],stage4_12[0]}
   );
   gpc1_1 gpc380 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc381 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc382 (
      {stage3_2[0]},
      {stage4_2[0]}
   );
   gpc1_1 gpc383 (
      {stage3_3[0]},
      {stage4_3[0]}
   );
   gpc1_1 gpc384 (
      {stage3_4[0]},
      {stage4_4[0]}
   );
   gpc1_1 gpc385 (
      {stage3_5[0]},
      {stage4_5[0]}
   );
   gpc1_1 gpc386 (
      {stage3_6[0]},
      {stage4_6[0]}
   );
   gpc1_1 gpc387 (
      {stage3_9[4]},
      {stage4_9[1]}
   );
   gpc1_1 gpc388 (
      {stage3_9[5]},
      {stage4_9[2]}
   );
   gpc1_1 gpc389 (
      {stage3_10[0]},
      {stage4_10[1]}
   );
   gpc1_1 gpc390 (
      {stage3_10[1]},
      {stage4_10[2]}
   );
   gpc1_1 gpc391 (
      {stage3_11[0]},
      {stage4_11[1]}
   );
   gpc1_1 gpc392 (
      {stage3_11[1]},
      {stage4_11[2]}
   );
   gpc1_1 gpc393 (
      {stage3_13[0]},
      {stage4_13[1]}
   );
   gpc1_1 gpc394 (
      {stage3_13[1]},
      {stage4_13[2]}
   );
   gpc1_1 gpc395 (
      {stage3_13[2]},
      {stage4_13[3]}
   );
   gpc1_1 gpc396 (
      {stage3_13[3]},
      {stage4_13[4]}
   );
   gpc1_1 gpc397 (
      {stage3_15[0]},
      {stage4_15[1]}
   );
   gpc1_1 gpc398 (
      {stage3_15[1]},
      {stage4_15[2]}
   );
   gpc1_1 gpc399 (
      {stage3_16[0]},
      {stage4_16[1]}
   );
   gpc1_1 gpc400 (
      {stage3_16[1]},
      {stage4_16[2]}
   );
   gpc1_1 gpc401 (
      {stage3_16[2]},
      {stage4_16[3]}
   );
   gpc1_1 gpc402 (
      {stage3_16[3]},
      {stage4_16[4]}
   );
   gpc1_1 gpc403 (
      {stage3_16[4]},
      {stage4_16[5]}
   );
   gpc1_1 gpc404 (
      {stage3_16[5]},
      {stage4_16[6]}
   );
   gpc1_1 gpc405 (
      {stage3_17[0]},
      {stage4_17[0]}
   );
   gpc1_1 gpc406 (
      {stage3_17[1]},
      {stage4_17[1]}
   );
   gpc1_1 gpc407 (
      {stage3_17[2]},
      {stage4_17[2]}
   );
   gpc1_1 gpc408 (
      {stage3_17[3]},
      {stage4_17[3]}
   );
   gpc1_1 gpc409 (
      {stage3_17[4]},
      {stage4_17[4]}
   );
   gpc1_1 gpc410 (
      {stage3_18[0]},
      {stage4_18[0]}
   );
   gpc1_1 gpc411 (
      {stage3_18[1]},
      {stage4_18[1]}
   );
   gpc1_1 gpc412 (
      {stage3_18[2]},
      {stage4_18[2]}
   );
   gpc1_1 gpc413 (
      {stage3_18[3]},
      {stage4_18[3]}
   );
   gpc1_1 gpc414 (
      {stage3_18[4]},
      {stage4_18[4]}
   );
   gpc1_1 gpc415 (
      {stage3_18[5]},
      {stage4_18[5]}
   );
   gpc1_1 gpc416 (
      {stage3_18[6]},
      {stage4_18[6]}
   );
   gpc1_1 gpc417 (
      {stage3_18[7]},
      {stage4_18[7]}
   );
   gpc1_1 gpc418 (
      {stage3_18[8]},
      {stage4_18[8]}
   );
   gpc1_1 gpc419 (
      {stage3_18[9]},
      {stage4_18[9]}
   );
   gpc1_1 gpc420 (
      {stage3_18[10]},
      {stage4_18[10]}
   );
   gpc1_1 gpc421 (
      {stage3_18[11]},
      {stage4_18[11]}
   );
   gpc1_1 gpc422 (
      {stage3_18[12]},
      {stage4_18[12]}
   );
   gpc1_1 gpc423 (
      {stage3_18[13]},
      {stage4_18[13]}
   );
   gpc1_1 gpc424 (
      {stage3_18[14]},
      {stage4_18[14]}
   );
   gpc1_1 gpc425 (
      {stage3_19[0]},
      {stage4_19[0]}
   );
   gpc1_1 gpc426 (
      {stage3_19[1]},
      {stage4_19[1]}
   );
   gpc1_1 gpc427 (
      {stage3_19[2]},
      {stage4_19[2]}
   );
   gpc1_1 gpc428 (
      {stage3_19[3]},
      {stage4_19[3]}
   );
   gpc1_1 gpc429 (
      {stage3_19[4]},
      {stage4_19[4]}
   );
   gpc1_1 gpc430 (
      {stage3_19[5]},
      {stage4_19[5]}
   );
   gpc1_1 gpc431 (
      {stage3_20[0]},
      {stage4_20[0]}
   );
   gpc1_1 gpc432 (
      {stage3_20[1]},
      {stage4_20[1]}
   );
   gpc1_1 gpc433 (
      {stage3_20[2]},
      {stage4_20[2]}
   );
   gpc1_1 gpc434 (
      {stage3_20[3]},
      {stage4_20[3]}
   );
   gpc1_1 gpc435 (
      {stage3_21[0]},
      {stage4_21[0]}
   );
   gpc1_1 gpc436 (
      {stage3_21[1]},
      {stage4_21[1]}
   );
   gpc1_1 gpc437 (
      {stage3_21[2]},
      {stage4_21[2]}
   );
   gpc1_1 gpc438 (
      {stage3_21[3]},
      {stage4_21[3]}
   );
   gpc1_1 gpc439 (
      {stage3_22[0]},
      {stage4_22[0]}
   );
   gpc1_1 gpc440 (
      {stage3_22[1]},
      {stage4_22[1]}
   );
   gpc1_1 gpc441 (
      {stage3_22[2]},
      {stage4_22[2]}
   );
   gpc1_1 gpc442 (
      {stage3_23[0]},
      {stage4_23[0]}
   );
   gpc1_1 gpc443 (
      {stage3_23[1]},
      {stage4_23[1]}
   );
   gpc1_1 gpc444 (
      {stage3_23[2]},
      {stage4_23[2]}
   );
   gpc1_1 gpc445 (
      {stage3_23[3]},
      {stage4_23[3]}
   );
   gpc1_1 gpc446 (
      {stage3_23[4]},
      {stage4_23[4]}
   );
   gpc1_1 gpc447 (
      {stage3_23[5]},
      {stage4_23[5]}
   );
   gpc1_1 gpc448 (
      {stage3_23[6]},
      {stage4_23[6]}
   );
   gpc1_1 gpc449 (
      {stage3_23[7]},
      {stage4_23[7]}
   );
   gpc1_1 gpc450 (
      {stage3_24[0]},
      {stage4_24[0]}
   );
   gpc1_1 gpc451 (
      {stage3_24[1]},
      {stage4_24[1]}
   );
   gpc1_1 gpc452 (
      {stage3_24[2]},
      {stage4_24[2]}
   );
   gpc1_1 gpc453 (
      {stage3_24[3]},
      {stage4_24[3]}
   );
   gpc1_1 gpc454 (
      {stage3_24[4]},
      {stage4_24[4]}
   );
   gpc1_1 gpc455 (
      {stage3_24[5]},
      {stage4_24[5]}
   );
   gpc1_1 gpc456 (
      {stage3_25[0]},
      {stage4_25[0]}
   );
   gpc1_1 gpc457 (
      {stage3_25[1]},
      {stage4_25[1]}
   );
   gpc1_1 gpc458 (
      {stage3_25[2]},
      {stage4_25[2]}
   );
   gpc1_1 gpc459 (
      {stage3_25[3]},
      {stage4_25[3]}
   );
   gpc1_1 gpc460 (
      {stage3_26[0]},
      {stage4_26[0]}
   );
   gpc1_1 gpc461 (
      {stage3_26[1]},
      {stage4_26[1]}
   );
   gpc1_1 gpc462 (
      {stage3_26[2]},
      {stage4_26[2]}
   );
   gpc1_1 gpc463 (
      {stage3_27[0]},
      {stage4_27[0]}
   );
   gpc1_1 gpc464 (
      {stage3_27[1]},
      {stage4_27[1]}
   );
   gpc1_1 gpc465 (
      {stage3_28[0]},
      {stage4_28[0]}
   );
   gpc1343_5 gpc466 (
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0], stage4_10[1], stage4_10[2], 1'b0},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[0]}
   );
   gpc607_5 gpc467 (
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[0],stage5_18[0],stage5_17[0],stage5_16[0]}
   );
   gpc615_5 gpc468 (
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4]},
      {stage4_18[6]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[1],stage5_18[1],stage5_17[1]}
   );
   gpc1_1 gpc469 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc470 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc471 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc472 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc473 (
      {stage4_4[0]},
      {stage5_4[0]}
   );
   gpc1_1 gpc474 (
      {stage4_5[0]},
      {stage5_5[0]}
   );
   gpc1_1 gpc475 (
      {stage4_6[0]},
      {stage5_6[0]}
   );
   gpc1_1 gpc476 (
      {stage4_7[0]},
      {stage5_7[0]}
   );
   gpc1_1 gpc477 (
      {stage4_8[0]},
      {stage5_8[0]}
   );
   gpc1_1 gpc478 (
      {stage4_13[0]},
      {stage5_13[1]}
   );
   gpc1_1 gpc479 (
      {stage4_13[1]},
      {stage5_13[2]}
   );
   gpc1_1 gpc480 (
      {stage4_13[2]},
      {stage5_13[3]}
   );
   gpc1_1 gpc481 (
      {stage4_13[3]},
      {stage5_13[4]}
   );
   gpc1_1 gpc482 (
      {stage4_13[4]},
      {stage5_13[5]}
   );
   gpc1_1 gpc483 (
      {stage4_14[0]},
      {stage5_14[0]}
   );
   gpc1_1 gpc484 (
      {stage4_15[0]},
      {stage5_15[0]}
   );
   gpc1_1 gpc485 (
      {stage4_15[1]},
      {stage5_15[1]}
   );
   gpc1_1 gpc486 (
      {stage4_15[2]},
      {stage5_15[2]}
   );
   gpc1_1 gpc487 (
      {stage4_18[7]},
      {stage5_18[2]}
   );
   gpc1_1 gpc488 (
      {stage4_18[8]},
      {stage5_18[3]}
   );
   gpc1_1 gpc489 (
      {stage4_18[9]},
      {stage5_18[4]}
   );
   gpc1_1 gpc490 (
      {stage4_18[10]},
      {stage5_18[5]}
   );
   gpc1_1 gpc491 (
      {stage4_18[11]},
      {stage5_18[6]}
   );
   gpc1_1 gpc492 (
      {stage4_18[12]},
      {stage5_18[7]}
   );
   gpc1_1 gpc493 (
      {stage4_18[13]},
      {stage5_18[8]}
   );
   gpc1_1 gpc494 (
      {stage4_18[14]},
      {stage5_18[9]}
   );
   gpc1_1 gpc495 (
      {stage4_20[0]},
      {stage5_20[2]}
   );
   gpc1_1 gpc496 (
      {stage4_20[1]},
      {stage5_20[3]}
   );
   gpc1_1 gpc497 (
      {stage4_20[2]},
      {stage5_20[4]}
   );
   gpc1_1 gpc498 (
      {stage4_20[3]},
      {stage5_20[5]}
   );
   gpc1_1 gpc499 (
      {stage4_21[0]},
      {stage5_21[1]}
   );
   gpc1_1 gpc500 (
      {stage4_21[1]},
      {stage5_21[2]}
   );
   gpc1_1 gpc501 (
      {stage4_21[2]},
      {stage5_21[3]}
   );
   gpc1_1 gpc502 (
      {stage4_21[3]},
      {stage5_21[4]}
   );
   gpc1_1 gpc503 (
      {stage4_22[0]},
      {stage5_22[0]}
   );
   gpc1_1 gpc504 (
      {stage4_22[1]},
      {stage5_22[1]}
   );
   gpc1_1 gpc505 (
      {stage4_22[2]},
      {stage5_22[2]}
   );
   gpc1_1 gpc506 (
      {stage4_23[0]},
      {stage5_23[0]}
   );
   gpc1_1 gpc507 (
      {stage4_23[1]},
      {stage5_23[1]}
   );
   gpc1_1 gpc508 (
      {stage4_23[2]},
      {stage5_23[2]}
   );
   gpc1_1 gpc509 (
      {stage4_23[3]},
      {stage5_23[3]}
   );
   gpc1_1 gpc510 (
      {stage4_23[4]},
      {stage5_23[4]}
   );
   gpc1_1 gpc511 (
      {stage4_23[5]},
      {stage5_23[5]}
   );
   gpc1_1 gpc512 (
      {stage4_23[6]},
      {stage5_23[6]}
   );
   gpc1_1 gpc513 (
      {stage4_23[7]},
      {stage5_23[7]}
   );
   gpc1_1 gpc514 (
      {stage4_24[0]},
      {stage5_24[0]}
   );
   gpc1_1 gpc515 (
      {stage4_24[1]},
      {stage5_24[1]}
   );
   gpc1_1 gpc516 (
      {stage4_24[2]},
      {stage5_24[2]}
   );
   gpc1_1 gpc517 (
      {stage4_24[3]},
      {stage5_24[3]}
   );
   gpc1_1 gpc518 (
      {stage4_24[4]},
      {stage5_24[4]}
   );
   gpc1_1 gpc519 (
      {stage4_24[5]},
      {stage5_24[5]}
   );
   gpc1_1 gpc520 (
      {stage4_25[0]},
      {stage5_25[0]}
   );
   gpc1_1 gpc521 (
      {stage4_25[1]},
      {stage5_25[1]}
   );
   gpc1_1 gpc522 (
      {stage4_25[2]},
      {stage5_25[2]}
   );
   gpc1_1 gpc523 (
      {stage4_25[3]},
      {stage5_25[3]}
   );
   gpc1_1 gpc524 (
      {stage4_26[0]},
      {stage5_26[0]}
   );
   gpc1_1 gpc525 (
      {stage4_26[1]},
      {stage5_26[1]}
   );
   gpc1_1 gpc526 (
      {stage4_26[2]},
      {stage5_26[2]}
   );
   gpc1_1 gpc527 (
      {stage4_27[0]},
      {stage5_27[0]}
   );
   gpc1_1 gpc528 (
      {stage4_27[1]},
      {stage5_27[1]}
   );
   gpc1_1 gpc529 (
      {stage4_28[0]},
      {stage5_28[0]}
   );
   gpc1316_5 gpc530 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[0]},
      {stage5_15[0], stage5_15[1], stage5_15[2]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[0],stage6_13[0]}
   );
   gpc607_5 gpc531 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5], stage5_18[6]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage6_22[0],stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[0]}
   );
   gpc1_1 gpc532 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc533 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc534 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc535 (
      {stage5_3[0]},
      {stage6_3[0]}
   );
   gpc1_1 gpc536 (
      {stage5_4[0]},
      {stage6_4[0]}
   );
   gpc1_1 gpc537 (
      {stage5_5[0]},
      {stage6_5[0]}
   );
   gpc1_1 gpc538 (
      {stage5_6[0]},
      {stage6_6[0]}
   );
   gpc1_1 gpc539 (
      {stage5_7[0]},
      {stage6_7[0]}
   );
   gpc1_1 gpc540 (
      {stage5_8[0]},
      {stage6_8[0]}
   );
   gpc1_1 gpc541 (
      {stage5_9[0]},
      {stage6_9[0]}
   );
   gpc1_1 gpc542 (
      {stage5_10[0]},
      {stage6_10[0]}
   );
   gpc1_1 gpc543 (
      {stage5_11[0]},
      {stage6_11[0]}
   );
   gpc1_1 gpc544 (
      {stage5_12[0]},
      {stage6_12[0]}
   );
   gpc1_1 gpc545 (
      {stage5_17[0]},
      {stage6_17[1]}
   );
   gpc1_1 gpc546 (
      {stage5_17[1]},
      {stage6_17[2]}
   );
   gpc1_1 gpc547 (
      {stage5_18[7]},
      {stage6_18[1]}
   );
   gpc1_1 gpc548 (
      {stage5_18[8]},
      {stage6_18[2]}
   );
   gpc1_1 gpc549 (
      {stage5_18[9]},
      {stage6_18[3]}
   );
   gpc1_1 gpc550 (
      {stage5_19[0]},
      {stage6_19[1]}
   );
   gpc1_1 gpc551 (
      {stage5_19[1]},
      {stage6_19[2]}
   );
   gpc1_1 gpc552 (
      {stage5_21[0]},
      {stage6_21[1]}
   );
   gpc1_1 gpc553 (
      {stage5_21[1]},
      {stage6_21[2]}
   );
   gpc1_1 gpc554 (
      {stage5_21[2]},
      {stage6_21[3]}
   );
   gpc1_1 gpc555 (
      {stage5_21[3]},
      {stage6_21[4]}
   );
   gpc1_1 gpc556 (
      {stage5_21[4]},
      {stage6_21[5]}
   );
   gpc1_1 gpc557 (
      {stage5_22[0]},
      {stage6_22[1]}
   );
   gpc1_1 gpc558 (
      {stage5_22[1]},
      {stage6_22[2]}
   );
   gpc1_1 gpc559 (
      {stage5_22[2]},
      {stage6_22[3]}
   );
   gpc1_1 gpc560 (
      {stage5_23[0]},
      {stage6_23[0]}
   );
   gpc1_1 gpc561 (
      {stage5_23[1]},
      {stage6_23[1]}
   );
   gpc1_1 gpc562 (
      {stage5_23[2]},
      {stage6_23[2]}
   );
   gpc1_1 gpc563 (
      {stage5_23[3]},
      {stage6_23[3]}
   );
   gpc1_1 gpc564 (
      {stage5_23[4]},
      {stage6_23[4]}
   );
   gpc1_1 gpc565 (
      {stage5_23[5]},
      {stage6_23[5]}
   );
   gpc1_1 gpc566 (
      {stage5_23[6]},
      {stage6_23[6]}
   );
   gpc1_1 gpc567 (
      {stage5_23[7]},
      {stage6_23[7]}
   );
   gpc1_1 gpc568 (
      {stage5_24[0]},
      {stage6_24[0]}
   );
   gpc1_1 gpc569 (
      {stage5_24[1]},
      {stage6_24[1]}
   );
   gpc1_1 gpc570 (
      {stage5_24[2]},
      {stage6_24[2]}
   );
   gpc1_1 gpc571 (
      {stage5_24[3]},
      {stage6_24[3]}
   );
   gpc1_1 gpc572 (
      {stage5_24[4]},
      {stage6_24[4]}
   );
   gpc1_1 gpc573 (
      {stage5_24[5]},
      {stage6_24[5]}
   );
   gpc1_1 gpc574 (
      {stage5_25[0]},
      {stage6_25[0]}
   );
   gpc1_1 gpc575 (
      {stage5_25[1]},
      {stage6_25[1]}
   );
   gpc1_1 gpc576 (
      {stage5_25[2]},
      {stage6_25[2]}
   );
   gpc1_1 gpc577 (
      {stage5_25[3]},
      {stage6_25[3]}
   );
   gpc1_1 gpc578 (
      {stage5_26[0]},
      {stage6_26[0]}
   );
   gpc1_1 gpc579 (
      {stage5_26[1]},
      {stage6_26[1]}
   );
   gpc1_1 gpc580 (
      {stage5_26[2]},
      {stage6_26[2]}
   );
   gpc1_1 gpc581 (
      {stage5_27[0]},
      {stage6_27[0]}
   );
   gpc1_1 gpc582 (
      {stage5_27[1]},
      {stage6_27[1]}
   );
   gpc1_1 gpc583 (
      {stage5_28[0]},
      {stage6_28[0]}
   );
   gpc1343_5 gpc584 (
      {stage6_17[0], stage6_17[1], stage6_17[2]},
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3]},
      {stage6_19[0], stage6_19[1], stage6_19[2]},
      {stage6_20[0]},
      {stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[0],stage7_17[0]}
   );
   gpc1_1 gpc585 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc586 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc587 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc588 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc589 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc590 (
      {stage6_5[0]},
      {stage7_5[0]}
   );
   gpc1_1 gpc591 (
      {stage6_6[0]},
      {stage7_6[0]}
   );
   gpc1_1 gpc592 (
      {stage6_7[0]},
      {stage7_7[0]}
   );
   gpc1_1 gpc593 (
      {stage6_8[0]},
      {stage7_8[0]}
   );
   gpc1_1 gpc594 (
      {stage6_9[0]},
      {stage7_9[0]}
   );
   gpc1_1 gpc595 (
      {stage6_10[0]},
      {stage7_10[0]}
   );
   gpc1_1 gpc596 (
      {stage6_11[0]},
      {stage7_11[0]}
   );
   gpc1_1 gpc597 (
      {stage6_12[0]},
      {stage7_12[0]}
   );
   gpc1_1 gpc598 (
      {stage6_13[0]},
      {stage7_13[0]}
   );
   gpc1_1 gpc599 (
      {stage6_14[0]},
      {stage7_14[0]}
   );
   gpc1_1 gpc600 (
      {stage6_15[0]},
      {stage7_15[0]}
   );
   gpc1_1 gpc601 (
      {stage6_16[0]},
      {stage7_16[0]}
   );
   gpc1_1 gpc602 (
      {stage6_21[0]},
      {stage7_21[1]}
   );
   gpc1_1 gpc603 (
      {stage6_21[1]},
      {stage7_21[2]}
   );
   gpc1_1 gpc604 (
      {stage6_21[2]},
      {stage7_21[3]}
   );
   gpc1_1 gpc605 (
      {stage6_21[3]},
      {stage7_21[4]}
   );
   gpc1_1 gpc606 (
      {stage6_21[4]},
      {stage7_21[5]}
   );
   gpc1_1 gpc607 (
      {stage6_21[5]},
      {stage7_21[6]}
   );
   gpc1_1 gpc608 (
      {stage6_22[0]},
      {stage7_22[0]}
   );
   gpc1_1 gpc609 (
      {stage6_22[1]},
      {stage7_22[1]}
   );
   gpc1_1 gpc610 (
      {stage6_22[2]},
      {stage7_22[2]}
   );
   gpc1_1 gpc611 (
      {stage6_22[3]},
      {stage7_22[3]}
   );
   gpc1_1 gpc612 (
      {stage6_23[0]},
      {stage7_23[0]}
   );
   gpc1_1 gpc613 (
      {stage6_23[1]},
      {stage7_23[1]}
   );
   gpc1_1 gpc614 (
      {stage6_23[2]},
      {stage7_23[2]}
   );
   gpc1_1 gpc615 (
      {stage6_23[3]},
      {stage7_23[3]}
   );
   gpc1_1 gpc616 (
      {stage6_23[4]},
      {stage7_23[4]}
   );
   gpc1_1 gpc617 (
      {stage6_23[5]},
      {stage7_23[5]}
   );
   gpc1_1 gpc618 (
      {stage6_23[6]},
      {stage7_23[6]}
   );
   gpc1_1 gpc619 (
      {stage6_23[7]},
      {stage7_23[7]}
   );
   gpc1_1 gpc620 (
      {stage6_24[0]},
      {stage7_24[0]}
   );
   gpc1_1 gpc621 (
      {stage6_24[1]},
      {stage7_24[1]}
   );
   gpc1_1 gpc622 (
      {stage6_24[2]},
      {stage7_24[2]}
   );
   gpc1_1 gpc623 (
      {stage6_24[3]},
      {stage7_24[3]}
   );
   gpc1_1 gpc624 (
      {stage6_24[4]},
      {stage7_24[4]}
   );
   gpc1_1 gpc625 (
      {stage6_24[5]},
      {stage7_24[5]}
   );
   gpc1_1 gpc626 (
      {stage6_25[0]},
      {stage7_25[0]}
   );
   gpc1_1 gpc627 (
      {stage6_25[1]},
      {stage7_25[1]}
   );
   gpc1_1 gpc628 (
      {stage6_25[2]},
      {stage7_25[2]}
   );
   gpc1_1 gpc629 (
      {stage6_25[3]},
      {stage7_25[3]}
   );
   gpc1_1 gpc630 (
      {stage6_26[0]},
      {stage7_26[0]}
   );
   gpc1_1 gpc631 (
      {stage6_26[1]},
      {stage7_26[1]}
   );
   gpc1_1 gpc632 (
      {stage6_26[2]},
      {stage7_26[2]}
   );
   gpc1_1 gpc633 (
      {stage6_27[0]},
      {stage7_27[0]}
   );
   gpc1_1 gpc634 (
      {stage6_27[1]},
      {stage7_27[1]}
   );
   gpc1_1 gpc635 (
      {stage6_28[0]},
      {stage7_28[0]}
   );
   gpc1_1 gpc636 (
      {stage7_0[0]},
      {stage8_0[0]}
   );
   gpc1_1 gpc637 (
      {stage7_1[0]},
      {stage8_1[0]}
   );
   gpc1_1 gpc638 (
      {stage7_2[0]},
      {stage8_2[0]}
   );
   gpc1_1 gpc639 (
      {stage7_3[0]},
      {stage8_3[0]}
   );
   gpc1_1 gpc640 (
      {stage7_4[0]},
      {stage8_4[0]}
   );
   gpc1_1 gpc641 (
      {stage7_5[0]},
      {stage8_5[0]}
   );
   gpc1_1 gpc642 (
      {stage7_6[0]},
      {stage8_6[0]}
   );
   gpc1_1 gpc643 (
      {stage7_7[0]},
      {stage8_7[0]}
   );
   gpc1_1 gpc644 (
      {stage7_8[0]},
      {stage8_8[0]}
   );
   gpc1_1 gpc645 (
      {stage7_9[0]},
      {stage8_9[0]}
   );
   gpc1_1 gpc646 (
      {stage7_10[0]},
      {stage8_10[0]}
   );
   gpc1_1 gpc647 (
      {stage7_11[0]},
      {stage8_11[0]}
   );
   gpc1_1 gpc648 (
      {stage7_12[0]},
      {stage8_12[0]}
   );
   gpc1_1 gpc649 (
      {stage7_13[0]},
      {stage8_13[0]}
   );
   gpc1_1 gpc650 (
      {stage7_14[0]},
      {stage8_14[0]}
   );
   gpc1_1 gpc651 (
      {stage7_15[0]},
      {stage8_15[0]}
   );
   gpc1_1 gpc652 (
      {stage7_16[0]},
      {stage8_16[0]}
   );
   gpc1_1 gpc653 (
      {stage7_17[0]},
      {stage8_17[0]}
   );
   gpc1_1 gpc654 (
      {stage7_18[0]},
      {stage8_18[0]}
   );
   gpc1_1 gpc655 (
      {stage7_19[0]},
      {stage8_19[0]}
   );
   gpc1_1 gpc656 (
      {stage7_20[0]},
      {stage8_20[0]}
   );
   gpc1_1 gpc657 (
      {stage7_21[0]},
      {stage8_21[0]}
   );
   gpc1_1 gpc658 (
      {stage7_21[1]},
      {stage8_21[1]}
   );
   gpc1_1 gpc659 (
      {stage7_21[2]},
      {stage8_21[2]}
   );
   gpc1_1 gpc660 (
      {stage7_21[3]},
      {stage8_21[3]}
   );
   gpc1_1 gpc661 (
      {stage7_21[4]},
      {stage8_21[4]}
   );
   gpc1_1 gpc662 (
      {stage7_21[5]},
      {stage8_21[5]}
   );
   gpc1_1 gpc663 (
      {stage7_21[6]},
      {stage8_21[6]}
   );
   gpc1_1 gpc664 (
      {stage7_22[0]},
      {stage8_22[0]}
   );
   gpc1_1 gpc665 (
      {stage7_22[1]},
      {stage8_22[1]}
   );
   gpc1_1 gpc666 (
      {stage7_22[2]},
      {stage8_22[2]}
   );
   gpc1_1 gpc667 (
      {stage7_22[3]},
      {stage8_22[3]}
   );
   gpc1_1 gpc668 (
      {stage7_23[0]},
      {stage8_23[0]}
   );
   gpc1_1 gpc669 (
      {stage7_23[1]},
      {stage8_23[1]}
   );
   gpc1_1 gpc670 (
      {stage7_23[2]},
      {stage8_23[2]}
   );
   gpc1_1 gpc671 (
      {stage7_23[3]},
      {stage8_23[3]}
   );
   gpc1_1 gpc672 (
      {stage7_23[4]},
      {stage8_23[4]}
   );
   gpc1_1 gpc673 (
      {stage7_23[5]},
      {stage8_23[5]}
   );
   gpc1_1 gpc674 (
      {stage7_23[6]},
      {stage8_23[6]}
   );
   gpc1_1 gpc675 (
      {stage7_23[7]},
      {stage8_23[7]}
   );
   gpc1_1 gpc676 (
      {stage7_24[0]},
      {stage8_24[0]}
   );
   gpc1_1 gpc677 (
      {stage7_24[1]},
      {stage8_24[1]}
   );
   gpc1_1 gpc678 (
      {stage7_24[2]},
      {stage8_24[2]}
   );
   gpc1_1 gpc679 (
      {stage7_24[3]},
      {stage8_24[3]}
   );
   gpc1_1 gpc680 (
      {stage7_24[4]},
      {stage8_24[4]}
   );
   gpc1_1 gpc681 (
      {stage7_24[5]},
      {stage8_24[5]}
   );
   gpc1_1 gpc682 (
      {stage7_25[0]},
      {stage8_25[0]}
   );
   gpc1_1 gpc683 (
      {stage7_25[1]},
      {stage8_25[1]}
   );
   gpc1_1 gpc684 (
      {stage7_25[2]},
      {stage8_25[2]}
   );
   gpc1_1 gpc685 (
      {stage7_25[3]},
      {stage8_25[3]}
   );
   gpc1_1 gpc686 (
      {stage7_26[0]},
      {stage8_26[0]}
   );
   gpc1_1 gpc687 (
      {stage7_26[1]},
      {stage8_26[1]}
   );
   gpc1_1 gpc688 (
      {stage7_26[2]},
      {stage8_26[2]}
   );
   gpc1_1 gpc689 (
      {stage7_27[0]},
      {stage8_27[0]}
   );
   gpc1_1 gpc690 (
      {stage7_27[1]},
      {stage8_27[1]}
   );
   gpc1_1 gpc691 (
      {stage7_28[0]},
      {stage8_28[0]}
   );
   gpc607_5 gpc692 (
      {stage8_21[0], stage8_21[1], stage8_21[2], stage8_21[3], stage8_21[4], stage8_21[5], stage8_21[6]},
      {stage8_23[0], stage8_23[1], stage8_23[2], stage8_23[3], stage8_23[4], stage8_23[5]},
      {stage9_25[0],stage9_24[0],stage9_23[0],stage9_22[0],stage9_21[0]}
   );
   gpc1_1 gpc693 (
      {stage8_0[0]},
      {stage9_0[0]}
   );
   gpc1_1 gpc694 (
      {stage8_1[0]},
      {stage9_1[0]}
   );
   gpc1_1 gpc695 (
      {stage8_2[0]},
      {stage9_2[0]}
   );
   gpc1_1 gpc696 (
      {stage8_3[0]},
      {stage9_3[0]}
   );
   gpc1_1 gpc697 (
      {stage8_4[0]},
      {stage9_4[0]}
   );
   gpc1_1 gpc698 (
      {stage8_5[0]},
      {stage9_5[0]}
   );
   gpc1_1 gpc699 (
      {stage8_6[0]},
      {stage9_6[0]}
   );
   gpc1_1 gpc700 (
      {stage8_7[0]},
      {stage9_7[0]}
   );
   gpc1_1 gpc701 (
      {stage8_8[0]},
      {stage9_8[0]}
   );
   gpc1_1 gpc702 (
      {stage8_9[0]},
      {stage9_9[0]}
   );
   gpc1_1 gpc703 (
      {stage8_10[0]},
      {stage9_10[0]}
   );
   gpc1_1 gpc704 (
      {stage8_11[0]},
      {stage9_11[0]}
   );
   gpc1_1 gpc705 (
      {stage8_12[0]},
      {stage9_12[0]}
   );
   gpc1_1 gpc706 (
      {stage8_13[0]},
      {stage9_13[0]}
   );
   gpc1_1 gpc707 (
      {stage8_14[0]},
      {stage9_14[0]}
   );
   gpc1_1 gpc708 (
      {stage8_15[0]},
      {stage9_15[0]}
   );
   gpc1_1 gpc709 (
      {stage8_16[0]},
      {stage9_16[0]}
   );
   gpc1_1 gpc710 (
      {stage8_17[0]},
      {stage9_17[0]}
   );
   gpc1_1 gpc711 (
      {stage8_18[0]},
      {stage9_18[0]}
   );
   gpc1_1 gpc712 (
      {stage8_19[0]},
      {stage9_19[0]}
   );
   gpc1_1 gpc713 (
      {stage8_20[0]},
      {stage9_20[0]}
   );
   gpc1_1 gpc714 (
      {stage8_22[0]},
      {stage9_22[1]}
   );
   gpc1_1 gpc715 (
      {stage8_22[1]},
      {stage9_22[2]}
   );
   gpc1_1 gpc716 (
      {stage8_22[2]},
      {stage9_22[3]}
   );
   gpc1_1 gpc717 (
      {stage8_22[3]},
      {stage9_22[4]}
   );
   gpc1_1 gpc718 (
      {stage8_23[6]},
      {stage9_23[1]}
   );
   gpc1_1 gpc719 (
      {stage8_23[7]},
      {stage9_23[2]}
   );
   gpc1_1 gpc720 (
      {stage8_24[0]},
      {stage9_24[1]}
   );
   gpc1_1 gpc721 (
      {stage8_24[1]},
      {stage9_24[2]}
   );
   gpc1_1 gpc722 (
      {stage8_24[2]},
      {stage9_24[3]}
   );
   gpc1_1 gpc723 (
      {stage8_24[3]},
      {stage9_24[4]}
   );
   gpc1_1 gpc724 (
      {stage8_24[4]},
      {stage9_24[5]}
   );
   gpc1_1 gpc725 (
      {stage8_24[5]},
      {stage9_24[6]}
   );
   gpc1_1 gpc726 (
      {stage8_25[0]},
      {stage9_25[1]}
   );
   gpc1_1 gpc727 (
      {stage8_25[1]},
      {stage9_25[2]}
   );
   gpc1_1 gpc728 (
      {stage8_25[2]},
      {stage9_25[3]}
   );
   gpc1_1 gpc729 (
      {stage8_25[3]},
      {stage9_25[4]}
   );
   gpc1_1 gpc730 (
      {stage8_26[0]},
      {stage9_26[0]}
   );
   gpc1_1 gpc731 (
      {stage8_26[1]},
      {stage9_26[1]}
   );
   gpc1_1 gpc732 (
      {stage8_26[2]},
      {stage9_26[2]}
   );
   gpc1_1 gpc733 (
      {stage8_27[0]},
      {stage9_27[0]}
   );
   gpc1_1 gpc734 (
      {stage8_27[1]},
      {stage9_27[1]}
   );
   gpc1_1 gpc735 (
      {stage8_28[0]},
      {stage9_28[0]}
   );
   gpc615_5 gpc736 (
      {stage9_22[0], stage9_22[1], stage9_22[2], stage9_22[3], stage9_22[4]},
      {stage9_23[0]},
      {stage9_24[0], stage9_24[1], stage9_24[2], stage9_24[3], stage9_24[4], stage9_24[5]},
      {stage10_26[0],stage10_25[0],stage10_24[0],stage10_23[0],stage10_22[0]}
   );
   gpc1_1 gpc737 (
      {stage9_0[0]},
      {stage10_0[0]}
   );
   gpc1_1 gpc738 (
      {stage9_1[0]},
      {stage10_1[0]}
   );
   gpc1_1 gpc739 (
      {stage9_2[0]},
      {stage10_2[0]}
   );
   gpc1_1 gpc740 (
      {stage9_3[0]},
      {stage10_3[0]}
   );
   gpc1_1 gpc741 (
      {stage9_4[0]},
      {stage10_4[0]}
   );
   gpc1_1 gpc742 (
      {stage9_5[0]},
      {stage10_5[0]}
   );
   gpc1_1 gpc743 (
      {stage9_6[0]},
      {stage10_6[0]}
   );
   gpc1_1 gpc744 (
      {stage9_7[0]},
      {stage10_7[0]}
   );
   gpc1_1 gpc745 (
      {stage9_8[0]},
      {stage10_8[0]}
   );
   gpc1_1 gpc746 (
      {stage9_9[0]},
      {stage10_9[0]}
   );
   gpc1_1 gpc747 (
      {stage9_10[0]},
      {stage10_10[0]}
   );
   gpc1_1 gpc748 (
      {stage9_11[0]},
      {stage10_11[0]}
   );
   gpc1_1 gpc749 (
      {stage9_12[0]},
      {stage10_12[0]}
   );
   gpc1_1 gpc750 (
      {stage9_13[0]},
      {stage10_13[0]}
   );
   gpc1_1 gpc751 (
      {stage9_14[0]},
      {stage10_14[0]}
   );
   gpc1_1 gpc752 (
      {stage9_15[0]},
      {stage10_15[0]}
   );
   gpc1_1 gpc753 (
      {stage9_16[0]},
      {stage10_16[0]}
   );
   gpc1_1 gpc754 (
      {stage9_17[0]},
      {stage10_17[0]}
   );
   gpc1_1 gpc755 (
      {stage9_18[0]},
      {stage10_18[0]}
   );
   gpc1_1 gpc756 (
      {stage9_19[0]},
      {stage10_19[0]}
   );
   gpc1_1 gpc757 (
      {stage9_20[0]},
      {stage10_20[0]}
   );
   gpc1_1 gpc758 (
      {stage9_21[0]},
      {stage10_21[0]}
   );
   gpc1_1 gpc759 (
      {stage9_23[1]},
      {stage10_23[1]}
   );
   gpc1_1 gpc760 (
      {stage9_23[2]},
      {stage10_23[2]}
   );
   gpc1_1 gpc761 (
      {stage9_24[6]},
      {stage10_24[1]}
   );
   gpc1_1 gpc762 (
      {stage9_25[0]},
      {stage10_25[1]}
   );
   gpc1_1 gpc763 (
      {stage9_25[1]},
      {stage10_25[2]}
   );
   gpc1_1 gpc764 (
      {stage9_25[2]},
      {stage10_25[3]}
   );
   gpc1_1 gpc765 (
      {stage9_25[3]},
      {stage10_25[4]}
   );
   gpc1_1 gpc766 (
      {stage9_25[4]},
      {stage10_25[5]}
   );
   gpc1_1 gpc767 (
      {stage9_26[0]},
      {stage10_26[1]}
   );
   gpc1_1 gpc768 (
      {stage9_26[1]},
      {stage10_26[2]}
   );
   gpc1_1 gpc769 (
      {stage9_26[2]},
      {stage10_26[3]}
   );
   gpc1_1 gpc770 (
      {stage9_27[0]},
      {stage10_27[0]}
   );
   gpc1_1 gpc771 (
      {stage9_27[1]},
      {stage10_27[1]}
   );
   gpc1_1 gpc772 (
      {stage9_28[0]},
      {stage10_28[0]}
   );
   gpc623_5 gpc773 (
      {stage10_23[0], stage10_23[1], stage10_23[2]},
      {stage10_24[0], stage10_24[1]},
      {stage10_25[0], stage10_25[1], stage10_25[2], stage10_25[3], stage10_25[4], stage10_25[5]},
      {stage11_27[0],stage11_26[0],stage11_25[0],stage11_24[0],stage11_23[0]}
   );
   gpc1_1 gpc774 (
      {stage10_0[0]},
      {stage11_0[0]}
   );
   gpc1_1 gpc775 (
      {stage10_1[0]},
      {stage11_1[0]}
   );
   gpc1_1 gpc776 (
      {stage10_2[0]},
      {stage11_2[0]}
   );
   gpc1_1 gpc777 (
      {stage10_3[0]},
      {stage11_3[0]}
   );
   gpc1_1 gpc778 (
      {stage10_4[0]},
      {stage11_4[0]}
   );
   gpc1_1 gpc779 (
      {stage10_5[0]},
      {stage11_5[0]}
   );
   gpc1_1 gpc780 (
      {stage10_6[0]},
      {stage11_6[0]}
   );
   gpc1_1 gpc781 (
      {stage10_7[0]},
      {stage11_7[0]}
   );
   gpc1_1 gpc782 (
      {stage10_8[0]},
      {stage11_8[0]}
   );
   gpc1_1 gpc783 (
      {stage10_9[0]},
      {stage11_9[0]}
   );
   gpc1_1 gpc784 (
      {stage10_10[0]},
      {stage11_10[0]}
   );
   gpc1_1 gpc785 (
      {stage10_11[0]},
      {stage11_11[0]}
   );
   gpc1_1 gpc786 (
      {stage10_12[0]},
      {stage11_12[0]}
   );
   gpc1_1 gpc787 (
      {stage10_13[0]},
      {stage11_13[0]}
   );
   gpc1_1 gpc788 (
      {stage10_14[0]},
      {stage11_14[0]}
   );
   gpc1_1 gpc789 (
      {stage10_15[0]},
      {stage11_15[0]}
   );
   gpc1_1 gpc790 (
      {stage10_16[0]},
      {stage11_16[0]}
   );
   gpc1_1 gpc791 (
      {stage10_17[0]},
      {stage11_17[0]}
   );
   gpc1_1 gpc792 (
      {stage10_18[0]},
      {stage11_18[0]}
   );
   gpc1_1 gpc793 (
      {stage10_19[0]},
      {stage11_19[0]}
   );
   gpc1_1 gpc794 (
      {stage10_20[0]},
      {stage11_20[0]}
   );
   gpc1_1 gpc795 (
      {stage10_21[0]},
      {stage11_21[0]}
   );
   gpc1_1 gpc796 (
      {stage10_22[0]},
      {stage11_22[0]}
   );
   gpc1_1 gpc797 (
      {stage10_26[0]},
      {stage11_26[1]}
   );
   gpc1_1 gpc798 (
      {stage10_26[1]},
      {stage11_26[2]}
   );
   gpc1_1 gpc799 (
      {stage10_26[2]},
      {stage11_26[3]}
   );
   gpc1_1 gpc800 (
      {stage10_26[3]},
      {stage11_26[4]}
   );
   gpc1_1 gpc801 (
      {stage10_27[0]},
      {stage11_27[1]}
   );
   gpc1_1 gpc802 (
      {stage10_27[1]},
      {stage11_27[2]}
   );
   gpc1_1 gpc803 (
      {stage10_28[0]},
      {stage11_28[0]}
   );
   gpc2135_5 gpc804 (
      {stage11_26[0], stage11_26[1], stage11_26[2], stage11_26[3], stage11_26[4]},
      {stage11_27[0], stage11_27[1], stage11_27[2]},
      {stage11_28[0]},
      {1'b0, 1'b0},
      {stage12_29[0],stage12_28[0],stage12_27[0],stage12_26[0]}
   );
   gpc1_1 gpc805 (
      {stage11_0[0]},
      {stage12_0[0]}
   );
   gpc1_1 gpc806 (
      {stage11_1[0]},
      {stage12_1[0]}
   );
   gpc1_1 gpc807 (
      {stage11_2[0]},
      {stage12_2[0]}
   );
   gpc1_1 gpc808 (
      {stage11_3[0]},
      {stage12_3[0]}
   );
   gpc1_1 gpc809 (
      {stage11_4[0]},
      {stage12_4[0]}
   );
   gpc1_1 gpc810 (
      {stage11_5[0]},
      {stage12_5[0]}
   );
   gpc1_1 gpc811 (
      {stage11_6[0]},
      {stage12_6[0]}
   );
   gpc1_1 gpc812 (
      {stage11_7[0]},
      {stage12_7[0]}
   );
   gpc1_1 gpc813 (
      {stage11_8[0]},
      {stage12_8[0]}
   );
   gpc1_1 gpc814 (
      {stage11_9[0]},
      {stage12_9[0]}
   );
   gpc1_1 gpc815 (
      {stage11_10[0]},
      {stage12_10[0]}
   );
   gpc1_1 gpc816 (
      {stage11_11[0]},
      {stage12_11[0]}
   );
   gpc1_1 gpc817 (
      {stage11_12[0]},
      {stage12_12[0]}
   );
   gpc1_1 gpc818 (
      {stage11_13[0]},
      {stage12_13[0]}
   );
   gpc1_1 gpc819 (
      {stage11_14[0]},
      {stage12_14[0]}
   );
   gpc1_1 gpc820 (
      {stage11_15[0]},
      {stage12_15[0]}
   );
   gpc1_1 gpc821 (
      {stage11_16[0]},
      {stage12_16[0]}
   );
   gpc1_1 gpc822 (
      {stage11_17[0]},
      {stage12_17[0]}
   );
   gpc1_1 gpc823 (
      {stage11_18[0]},
      {stage12_18[0]}
   );
   gpc1_1 gpc824 (
      {stage11_19[0]},
      {stage12_19[0]}
   );
   gpc1_1 gpc825 (
      {stage11_20[0]},
      {stage12_20[0]}
   );
   gpc1_1 gpc826 (
      {stage11_21[0]},
      {stage12_21[0]}
   );
   gpc1_1 gpc827 (
      {stage11_22[0]},
      {stage12_22[0]}
   );
   gpc1_1 gpc828 (
      {stage11_23[0]},
      {stage12_23[0]}
   );
   gpc1_1 gpc829 (
      {stage11_24[0]},
      {stage12_24[0]}
   );
   gpc1_1 gpc830 (
      {stage11_25[0]},
      {stage12_25[0]}
   );
endmodule
