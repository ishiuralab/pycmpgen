module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [20:0] src22;
    reg [19:0] src23;
    reg [18:0] src24;
    reg [17:0] src25;
    reg [16:0] src26;
    reg [15:0] src27;
    reg [14:0] src28;
    reg [13:0] src29;
    reg [12:0] src30;
    reg [11:0] src31;
    reg [10:0] src32;
    reg [9:0] src33;
    reg [8:0] src34;
    reg [7:0] src35;
    reg [6:0] src36;
    reg [5:0] src37;
    reg [4:0] src38;
    reg [3:0] src39;
    reg [2:0] src40;
    reg [1:0] src41;
    reg [0:0] src42;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [43:0] srcsum;
    wire [43:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3])<<39) + ((src40[0] + src40[1] + src40[2])<<40) + ((src41[0] + src41[1])<<41) + ((src42[0])<<42);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9797185716de642772cb6a5f9f2b4ea9a48c82d85352adad44c3559a148709560f793a86cb3d1764b64faca959758be4542d6a963ffd08efd79ed2ef7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6edae7c7061bd79ab0b4fc06c1ebb5db0f3a466a13d8a019f1d54160daa8b26007709f862791ad90967ff8806593ce2c6fce4402a82952f66f56c3d3a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35c572a3f520204aa603b021713ef194e128d6d3907bf5df7bf4153b3288aa54eb49e622bc042d7dc95ebcbaef7686d370922847a4182770dfbc63140;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha091ea4b5061b548f515c819acdc8811611b07259c4fe84147ee13a14b4c81edc98a6ffe70ebe4c31cdae27e85e1cd612a17a43eb9c9085b82e19c063;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9052609c2148f7a81c6bb225e2795949e98d6fd3e9ecdbf1ab74195375c7c3e55404f3d02117e04632b2b086d8487cbe261900dc7d9499abf52fbd2fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1fcc84c2d01c364bcefc3f1f56366b2635c10b3e43017c1603b8db043c23966ba08fc31abfdb998c3313eb52ed3f8787f66b7c9e9a4d3cfa0d3c958bd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha64631015c725cb3d1505b289e157aa78f3434df91c9f7a8aff315db4d6c21bb95778eb1d638d5c92838dd1a82c0b7db07be27c6594ddce71fcf9fd6f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3652dec45fac0eba30f5e1ff2fcf2e45437ae1660ceedd142f2d60f5678f68d496d836c804b98f38f1877f013a8cd87810cf90499d72164744d0adc36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b7882941f12a300292fae62cdf64f0871a17802f281bc704af5de678c23fd02549d74d4596c5dc120aea8540259ec2591d4de50ba02fbdda4289309f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31afacce20c613b3a4464b69cf470f8642f7abc899f5d923e9c3d44357b4ff60220b27fed9146f2bb686e72b1af523ddf514469d58ce681b3edaa0bff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7254b9f1a26f506e2c9fd9d7c3e8cc205beda33a5cfcf1d51d46b0c6d3b161265c46229d403c3a0252b172d25fca20a88259a13be3aa84a9ca2f7e7e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h274104b32ac6bd03e24d32a05d142fac39d41c16b375705916c645000ce9a5367c82dff9bae6d764363f47a49ad8ca37aece0bacf6bd724be5e5ef635;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h274380640505ec82b17e25a65f4ad38c70997548d10f22de39e180b0ab5f09347259810439fb04889dc39b5c6bbf5c2d3965063198306ee7fd7f1c801;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4e5cd0c6ad4d4bd7a7b3820fcdbe1ff18373ce6a7f1aaeec6d9be1be40dd2cf74c9b495577f02daa1d3aa2b81eba39b3a7a641830ecc751f31cfcd37;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c2d00a0ac726b130475dfe7d5110f04a10148011fb7e56e4ddfa3e5e9a90cbf9f50e802550b284a044c5cae93b0e4d038043c4c133045f7f570ad152;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6393591fd1312a61b36e00336ccee59b1f3b3bb6605975832611c268d5f46bd9d865a4b1702a3ab4b32daa7a0c8688227062bc8197a502d010cd7ada;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h845a2c2af5d09c41891e3b79992699ab10c603e7f4146bb8824647832a5aa73a1e90592af0d9f161976cc40829965efb59e14b017410883cec0d79ae9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66fac6e16232f0ce8e7a7d5acdc17a3c5008ac4dc3530de2f5813dc622a7fe3b347f0fbeacba14b0a8e3c33660fbe3e99204aaec61378f8913336bbfc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8291ce4ec2dfad7480613bc3b614838c9af8bf5440723793efaba7fd3c7157af17cbb31b473d4ad034065982772fcc44dc1969049eda09e10899209ee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e5de174bea36c1ab1b7f26cd36e1486dd5644eb479542c25d4d61b7629b16d2d8fe46c7d73890ade082d370f28e12e136676f476876492adadf5180a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfeb4f4944296973e88e205b30e4290e5986338d58f4517a12e9e8da577961ec965969edd4a2e5569d229c4ba8d25e94042b36cc94e4c2f0d7ade0a0f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab5edca511b89ed902d87a02dd2e7ecde8cf2ba6d492d6ae8634172eb92b12a25d31426d6c95f160ad0a0a542a13295b31f835ea03ef8a2d9f506f60c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6e35a2b1f3ebec19718cfd4c7c517ee548e92d6faca20f4e8d69bc3e3e35dc0cf55d9eea71d4b8fae7c056bb892b17e9680eb9d5657e7572c69105b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h426e71ea825a25bc62e2bc2dcd087c1a3c011918008c3c560c1c869e49ff48dbfaaab73f0ad0fa2f0939d3fe0176d94f53ed9fe2473cd703e9b4b4ff7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h748dee77992b53fb4843553d399e057e2eeb5cbc0466caf86ccdb4740de0cf94761fa840563419cd91a9aea24e645e527eabb6a607305b817dfc04084;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d0a6b67449c8ca085295856db566dcefb7439b1885ebe2540f89e68096ed47517e91ad48f2ffc32ddf3381b5888dd34c6ef8c4019aa7d2ef52dd502a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9498ad24f86e79b1c8adebb242157a8f5f9c86ca257544a777617270cd51697c1915b4969b190440d1f5ad5c490377b2ba018b8fdaf5ddf7d8869fd3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h489dbe89e0201da1d971d069d9ba5630cf6a4fa9ac355a76e6a8b5601f4d71cc100b64907ce0c63cefc2f9bf35e147982429b8af0d14f1b0b47278017;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h118ca893f06abd52a5fe2e07b522f98814f058ee84a064da7946e94ca7c352cf4666f6edd84ed1866fc860389f87cede9ad3d6aebae30ad732c36e6e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47b1b503c361245765827d6a4cbd3face91e6ff33f7d3fe5b88e93d9ddba619b1911dfe7fa2d32195ca8c2e8515f53e76fb95abe7ec900d479e4559bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ab4cd9448288a5e4e676dfe0af2386de6e4520bb7a60291ea7a2827b4e9c7a921162fa1182f6d1618ea9eb70b69da57971bb2976c424271ea23c909e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9455ffc67201094d9dde79a810d29b9a8c9d6edf5bc854a1361f7d701facb227aa05a48c65f850174abd37676752d2be664734f74fd88adc5ee11e913;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he382043b9449a702e9256c1debd04156f158f2a1a1e98c78de001298bcfea974546b47c6f3ae20ce0047009fd34870e0aad8f5b1018a3fcad3385d168;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b15fee924d25fa9294640dfd264d8e15cb4c089bc036b674aa80011dd22a8da0c9fba9067319dd61cbef87b2254a1a0568e86b7f89785f38e2fe96bd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35d111d3c1f386a9f591a906327ecca8dc2cd232731559188eae1bd4ac9c9f7dac9098ad3ee7f8fc471ea35083c10e866ee5a82dd948b50525fa55b25;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d766518c7cd724c4f67f13feb43004f20e06986d491366441b6fa5a6edba2af8a0097023d8aa20e8c442ff212dd36b19b1b05f7fa4101ed1a3456e98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ed74439f48d036c945bc472af547ca877a57b9f7d7a37eb0c9348daf6d89d76a3178513cbe02ddd80a3fa081b30213fb4634f907cb5c2d71250d9819;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5535c208231dadcbcee91dd1451ffffd872da5c2fb7572058094843a1b4cea77050075031dc6f49d61e3f6e2fd3ad5a62b50f1f541fe4d7dc90c6bf16;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4529f6933b1d8e57a84f98801a88f8ee57d5c8350876e8c3b776b18bf4981fff92fbf0d2ad748b56190a0f6f7670a1c8dbf64e9d89ae4570bcf3a8bbb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b1bc9c010fec70cf7860412bf04862cf1b26243cbf2d43db673f389b703a233e6859a744f866da4ab76a6c2606656282105938fcf8a3797c62d0b3f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9aefb7145dac2b17f93c3da9073a6b33df86aaebe885328da7d958f6e6d0e6ab793a7dc231b4349d8fbf34fef24de36c9717dc36fc5fbb695938dbf02;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86e0a9765d218a56ba2fca95c37f8e9058c85de7c33a82a849908ce9d83df347333a6593aae199f3769d0ab8dd676e91f9f3164aeb152d7651647d24e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0a66490867dfaedd8c6cf7c559dead4d992756f99f4a1257343820457219e8910b81ac1f25ffd46b782db62bbc8fd980019791ea7b9bf5ca59b5058c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h581fc4a2903fdedd31fb5b4d45707581cec5e8509053b0273bb5214112433ed49d84928f75799bfb617e717751761cc299c5bc034796d8b4a1bf2bb7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8fde5a749cbe78db94f6a2f3dbe697e5f0fabef105b47acdfba45a8188785b3c2ae03174703d1b2bd3a59b7062d4c09faca4ccba359d76e8b9fa4ddc4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8700458fdcf5d4884e117d24f7044e3d990ad3bbd88454e06e9ae24d77a029540b00947b6808bb5f41608930cc383078f1ed5fa8c98182b81a6711ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h976aebd25af9864c2f1195b888a442ff0b80f8586946dc86e0b313ff7f2e37b49a0ca5ef48d0d8d4a9cda165cc4ad6548373fffbd084ccf61db6a6cf3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf62662ca514fc59455b3a401db0cda941e2a93975ef978552378ac40d5e640c514968472d0fff75a2c87c872e40f5f5d744ff070f2dd0739084684d76;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d0d99472c24fc7921a50793266bb43483b6d88b78c834d847689965b49dd99aface74bbccaa777a652d677f5323370c645f1a4fd0245669873d0a467;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hee2e0a822b41338bec9d8c82317f31a27c90d4494a784ea4e74ab9ecff7734abd3cf988f02c55d6cbb2e082ea867d14d0e77fa5b45a5350e73afe7a39;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he103efbcf49a0b343ce54560ca44c54c1335d641f3e235f4b6d3b1cd8496c2872fb3062b6308c12c2bc658d25a7c35cb144b05152eeb47d115637514f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72fb0b567abe6164b775ee70815296f3362f05fc7dbf341e0ceaded21127bb6721593298876ecace47681c8e6989baffab9b7a915b0452dd577c91f1b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc976d26dd0a37ad371140f2ae29661ce9754c53e8afa7cf85c9985a49e5e498896cda79c6bda922cf4b4f964cc16c1b57e287c56023602bf7470be3a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4915229a315d7eff8815a4370eec0b21489ddb89efbf782c2640d882518f12c5b34ce0f568025e0dc493c103cd59b3e1dbf6c400554a9e8514d521a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85d77d9eb3c711cbb6e30c03a0d2bf4c7a84d7a7eab5f91feae865764dcc0704a06eedee811735c197cdde4af7752cf18495d1ba04b32e3f216c563de;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18168bbe6e6515977414a66f098f45c70d00c5e4bb4a3886c4e9cbdee6b43804f4d8285fb836cffc2303b54301f338bc2ef91641e4154833acfeb4b56;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7915bf651bc0769174aeeceb2886e91745f32868153c42cac50fd25540fcb2b3519373a932737a1e682083f493f185079bd0c3bc5909a0962ce0eaf09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ba344b2b4ebc961ce54d2451a8a2ad36b18d56a0aa5508d772b94b4b6d00a289226aa70678d7ccc90b1104e32761641cfeeb70272d72ff7558dc38b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ae941d5a18e8958b202493d1618eb07a2d47c09360ad7f6a2240eeb66dfb39264155ca2f6eb8b8cc8d14cb10cb617867336879ac4eda3bf2e46280b3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h517e31b1989ee65d9fb0636e7a8e827bd5d4891686d7eb6600a84dbc638220544ddc9e29b7d2ff12d1530edd6358295724c3935ec92805200b21b1ad3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11e4e283a995ca6075b65f72366fa767aef68b45ac24d518d2016fffd886b551348692cad5088d80079d8aefe9ffd495b7ceb3d147db91ed192f2f787;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1deb0ae9a045de1a5e6a68d5b4c35703cd97417367aef03ce5ff1c2520277ec455b6531955fb6363e4e5c56e02690a0fd018ba600acbf1ca875e1ca4e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3dd8a9a8c95354df079130b55a908181c957571300feaaa3d65c0edf16975e8e781def33abd4f65d2e2aef995dc9e4e474ff4a75eadfd9c18dc1149c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2a92ca67c326cb27aa9fe74bc90b3249dbc69c987f95d87f54af8386cf494ee2a86580b9b8903420f9fb37ff98dff09b6d7f6e90a75972d6c3e61f30;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heee94f2c94ef54fe8a54b0d9f34172381eabe3789dd8f975e6421f039794c58a1d888f8ccda1585c5a9bda90787ad45c79eb1641a0c8c178681d2bbf9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f8d60aa405930abef7f4d51c421ef112b46923a9c04e2094d8f049d92aa9f4b2f34442f6cd1d1cdbdc0af622e8cfee19afe31b67c6b3576e3178bcb3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5888ea92ea7fbba5606f33a5af3d85f0b41630f280f7b9dfaf5ec9921877c97ca9dd362a8963bfccf631e2c3f95cb97663d6b35198de5f1ea854432de;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2e383d3c225e2f98f7e9ff8c499665ecf570a8ca2380d12c40033a19515a8f67188c02428355bc1681e5b5ec3beb32180d52f4511491fe55186a6893;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae36573239c813bec80acdff355b481cf951f457aaa98b5778355f5f71cfebaab07b175c9f67eedf9a5ba22cd50d63aecddef9f342f9f7d45b2a64395;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a8215e2ea09f187404dece3b2a11af6e50ba39409e04299c6117c376f3f36db57f209eda2b0ba93b230bfcb8203a0358921f3ccb43e3dafde5c44dcf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha765c1969085de12bb9cf01bbfc90d5235feab052175cf7b48c2d050a47ddbcfe580f17f74d72e245a9cd939aace3cad6756327fd1a2ed6999e92164f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffb0e34ebf66ea8276ee9620e1994ca909be6199085e73bd868c0e8b60102fb7d5b6f44b9a511bc7180e6dfc54475b9b1e16c8ad5065852cbb8c5cc8a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1953b36eca6e8157dfdb888562e4784b65dd3d8307be9a7678ffb819e016ea946c39ccb8352450b4393357a180487e88578473193682000a2a324b6f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h172233bb2d1166ccc6497a9dd26068599a9420a36bcae4402ae3db4688a6e35d565ba7c17dff6c3f5b2e4fc61bf76310d6296c7d29e76e45dd83521a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h356e809c2ff7571fba0d215b1fbde7c7f77d63a91df8cff60ca4c598adbd675e19d71a9c982f7530edb4468cb4c075ec8388624a9b2a2749b4a30fb48;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ae363cc9995b8ea8274e3089dd1f79686a38876d790686cb741c3146ff94d43394d88e4c4483128077f6978a315fe907cbceea32281bb67e47a39750;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b6b8533fa36e0ace04ea4d578692ed133e241882b605ad69d5123f65e8074dc0f3f2b710a549f29b77ad171430dc80638784edf12842eada8f331b8c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb45b4f55e2dc6d295e14f228ca48bf91957a8b259ba763d8eaae25a426915f75ada208a681230da58ddc7ef908167d11e7c131e5861b897e5fc69c04e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e62b6ca1878f456b0beddbaa4fabfe66be40224b4b0e7b638dd894a8dec7032acb06f1a9036207c11a1ffae5ea62040d0a14a7158d33d5121494d76;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28507e2a97eea18f50540dc2a4cf3d50ee8b7b7b2473775b7e812b574fde2a03614efab3c22118e83d53e549bdbea3779aee8c3bdf7e654be045e526f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h809a07c08f34e34dd8f6bbcd84a50b2b4698c39ce8a0eea00307920ef73d0b89449003d261382cc53d63576192605a604dec89e39ddb17d32ffa926b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa775f3d0ff5eaf0790f41cc1120d2a9ebf2f157d69ad1386e1a107fc5b259aa92d32392c1514b85c6f89ba90d6d0d3c1557fa8f8222d4f7d7fd74756;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ac27f2a9179987c880767fe55950eb3567778278d678d7695d6cdcdaf1f2e24ef08e5f115cd3e8bfe5b8b7c11f964e97cb86a3e8b184400e36354cc5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63261ffbfc576c26b86e635e39054fcbc7e575410c39bd6067d804a6005f5dc30602542e51baa3b8dea9d26bdc653872bbeffd0257206f00a3aa88c20;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46da9c0c763bd7f453655890aaddebea0f1c53e3c73342f1c0258895bcf73fb353a667055633bfcc74d962ae41464f9d9eb6335ec96e70c936be55f87;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha80d0b6a0b4fbb14c8f28d4953dce024176769e31e2c3d70f67db620cea9e4eef5b227adfd78a36036ad971fff45249959e34a96137b4b830e08374;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfea9520065d40785f2cc11d0d2304ae43b391c82e0a0a83ce5dda8c977fa1cf70bc6eda0995212276b80699e7df363e76c95064ebe2a607afba9c0629;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a69b55a89f9a5ae023e943f7b02129bd0e06c67610b971742dc511ba70f1e3c2bd35b3eeb39f8a96a1eaffc94f62f0d8f85f636d96120c4fd9035182;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a43ca0502d76ac12b8041905a8a108341507554f509cb7df8a08d7ac2e5ba34187a68879898f3a33adb2c14ea48a7fb942a3cbcc24ac3d52d5cfe535;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb328ae83824fee25f732d5dd879c94394c790455398b425cb881dec2f1ca1f694f8b8a6387099266d3eff572eeb5d113c46c710c3154d649963173a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54913b4f45d91f0595dfb11dbd680a9903b99895de190b3549b4c0d5da47eafb05cbcf2b9212121a4f1cc77582a480614055124ade351ad59bcf844eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5357d36ed9e950ad1b6c8a62722819dd44db44e818ff169150dec714818c47f72fdb6477b8ac9e2585be58698672a88bf69dd8e2c82343752411346c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25bb6887cb563fd8adc1db9e8ca22bef5a4ee82b93b344d7d82dabe0655c4beee1ca1ea142032af48196d177dc5a67684f62cca37c157162d5961ea74;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a01b8313887d1117eefe2c2ce86f435c80b1570cf52059c10591bab347c1ff057218c5fd6f659bd10e88d598c47d4ae58d2bc7809d41d22f834290ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27225f4a91830d6d526830a075d54bcac7c53101ff37a3f0942f3f1088b8ada5ca788648f93b33364bc82034b9772fb0facb0302188c9e21290ddf343;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b95d879e1946d7f2863352de635d22c66e3aedcbb7ea0f61cc088e578a9bb8c667534e3a1d7dcbd76ad793e827262d39d0e66d7bbab26956f7059bf7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb65a2c2246733dde78a18d2d5cb43ffb8ec2b677d735e9c78db1fc4aef1b4431ac44b8248c6615e14ca4c03be7daac526503e18e7e5beff20a6915e2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84a7198df4b01f4ed3e9c348a7ffb529b5579d9f8658f46ad545d374cf2dd9291f7a145b13ebccb61f61bd46794a8c282ecceecab5cf7c290a736091b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5c81f9acb88b72bbec53146022912dece1245ec84c8a761999b1bca356ec9c09d56d75a0cac6bbc27e362ef91c787b6c6c4fa5ae83041c0dd443783b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h730cde1024ae0a0350b073d19b700474791d53da49bc17b175750ba6f548afece1c894bb6243dff8366eb050eccc143253695554183b399a6126c43f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h140b3487ff094a9ad6f551dc923df0fa0139bf335911d03ce9f247491293b1f2fc4104a5c2ea3d84f8712b553e0368b379edcce68e2525b88faeae19f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h388074713344d34d3828af79bfba45c9582352a3e1ff3042650c613662c6475b02a7dbbfbef80ad8d7e2cea1d44ee5d72406362bd7f8846e6e9b17b78;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b00213d4bd161fb9399e574f3328ebd14801e9910f9746572c4b4a899e21f6388270e96a7bbf2298289f4249d5fe66e33c0526c675f4189a03c5cf21;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36f22b3795544c5d64f31483915ee607b79a35a147dce8f3dfe51fb5affc34fa66e9b289ca94d54c36df4afbafe502ed9f193fb5205aabc7283d86650;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cd6fbea641a34b99fc3ad12a971701bd2327e090d7e6994229e67d5e7fe8ea4b4ccb409d53e6d69ebc285a2de87f707b420ea6b7e77a2c3f40c6703c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha2e1dbb59e0789e76ad0edec79d3514999ae04704997f613d85bc0b8ceb9b4ea26408a99c9881e260781bf19a3988dce41d23eb62b0d3d3e3d2e46d7a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h658300b765fda3fae6ee3f7607e043b46b6fd80b425c8d3621c0ba86c325b9b469d8af7d16370d941eaa2929f021e2fcd481cbb552cd0df22be3570e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95cd040847f2159d637c3cc99394fcf8fb602820f8622b0d890590fb72f70e50e3223d48257379deeb6bfe097e1bb1ce7c1782c7e8fe8fc3ba5c7a5de;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haefc5cc943a0358190e2926ed3dbea2633567dc2f0452407ecf2b0c727166274d742e488ba2137c3891c17ea01b425b6e056342f41caf81bf54f5b760;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1eb631c8f7e88c4e685b25c72da2ea682f3332657af9edb92aa2f83ba68b75a5ec8ca2055b156c316accae09c1081a9cc28fbfb66e5b96049214435ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3bb53734aa8fc3fbaaffc04b39d5d3ab33c19233743929f9bb68c7527bc237e54e2552fb5d5acd81a24934b07f6d76f3c1eaa298f8e06e1cc6476624c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h518774dd21345368836427b38178a951b9b0d9ec9fb9734ce484ad9b5bd1362bf0d82640080a41b852461c6612c15d52057ca96c7390d1eca82affa2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65fd3a203c5aed7e006bb1ed291bea0fa2d0f4fedbf43bc09d56d8c52d25606fa4ee5f6e6deb4b22bb111a69d0d4f16d1f7b831f572900e91006c2c09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h865e4d9cf6a5430912fd3cdea45c53625f5ef515a98c09e3bb1017686a29f388e17a1dd43988d9b7d1af0fb405e54b859960e16f89ece3f90682146e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91009612c0fc350cabd86fdc8c132846fde9aa0cc46a3915a2d576fc6254431f87530c1865d2183a78f22cad6945cb21092db76938e0b02d37fd2a15e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd93d53633bd46411d1bf37392cbec33e68d53ac0bf428696a27bab9560865c48e1baa25dfd997dca4de0fca3a1a3999b2556303b1885c0a57bf15aa10;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbeca6d6c109a472dc5ef35aeb6ed702f90afaea673755d56bc46045703f1476a711836bc58b8e0dea08cdc8f2478aa38ae20b0ab8ddcce7df35ee533b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c808db9fc8ebbb29fe3be9ef4b9794a81afe7dde552538f7c9e4d0bbed53f280acda03a22af1e4e2b411a47ad065c00a9ef5e4764dde72ac7be3336;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd1afb0d5c287ef32068e1a5f316715e2c8f8dc4b436db0ea0b01b23b9885072d05c7efa20d7218f1ee2dfab74ee5d1ede10c9cb482696fe57387a119b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd54afe6a0c13c353179254fed3cf860516b874b212dacf5cec64e387bebc832e2c4a031c25f8073a7442b67add0e9c4c8429d989a3f0d587745a2c714;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e3ecb6228959c5d839b9506b816c1864ecdf6af2e7ed9836838b395872b66afa45798cd767d6d44776aea148a7052742c758e7c33580aa8f49486204;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99266435a93175418147681456c5920ac493c14e99ff6ef10a296f18c94b16c18b92f1b5c5227f1762bc0aa821803f794f31f7ea383025f009dc4df1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f0f0596ef19a344dcb4b669e78dab9aba206edb585396177c845b1d88e7e8558a9800ab4db7a44ae306ed49c03b3fce2c009ee1fb84c82e296feb819;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5f887ec44b79972c678f7545bc1a9db80b942c3f2c22c82a7daed353dce2b9e61f5ed1a9963a5b2aba65b4208e8017471f38a29fc4d39813725e4e876;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c63a46c4dc41c32fcddfff881af31b4a477fea9972ea1894d1cf7b63f0e5e2d73f0ff40df36aa656174880b8e67a409ec4c06aa652bd30a48f3834df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb79de2822af81e5750c59ce15177836f73cdea1665b68b3552859f684f8c3aa350fd1ffc9e3177459e3770b19987d53b25522af4e5f0ad71883397ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h274d093d6e169ad8fd84f6a3c8a93738ca581b8852805b2592867114a207f99cd962bc9af4e9289252cde24c79b272b64ec87ca1a1ad5bcc2ad65c9c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8aca4e6454fe4c8cf21c1e6a443bc2079de5fdd784ce1ed59d28416b2b826b6d7ce58b1978da489488f1a1fa537c5059262283989870c6b9a3d68f1f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h323cb190062254ac84a1bd3dc94a6b5f1319ce079e82e8b0f09a766e884909d887855e4b73ff669ae6554a6b69da6f5232a2214a0c9ffed2ec992bf1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78c0f19d515b5922bad3618f15908927c1724e404c1794e1413c83e67997d9755be41f36905165837d8d06ccf6eef82782b168a25a9ec6f7552dd9579;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42291129ed908f4d56a471cb9931cf60f871a9d71853bb9a971d54a35c238b7c061fc5a2c7c38527d5ee1254c961fc33db4b0c68c9f9903cd152cc61f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92cc594d4c8fd5453715fc18818a405acc1ea374e42ce28388ee7e24c543c8d28155acd693eac2c3889e09b9eb909be3fa8fb6b27ab04d14c95d8cd7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h871d98c33862a3539151712c7772ca2d14b65b8da23182c79b6c0d161a2ddcf5cee14110197f0d446db41f125ca902ff7487f60ef62d967e789d2c705;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54e4e8cb0d0dc5ec5b6a7a5a5f63c47c8b2891ae8128efbb38b8891d3df1e7bf7c4af28921c5da8c96d0c7283aa942c7efc6714b2fb512f12e21e05f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3230d7e5cd349209632f2a5d20f399568ffb6f99811887fc034b184925025888a14737a7d4802801883bc884587804ef2f3c5e1fee352e587be86829f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbea7f7bf990597d8349f6aac3f84038184964eb15e0ff41509ac052098ef822f9a18520e2bae18ab816147e106253a1c1e6ccc47a3cb506380cadf2a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he374af91ef96bdce814a14a6de5eef31197433c2c6c21362e579246a44f2d94331156e3198a09fde3ffd27889c4e90895cd3792086c8fbd8479ca8e26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5e92a60b7c9e46af58c00780a54a3b22708c5b1bde76f041cd91bda1894c62de63a656dd653b50d12b155f940c43797132603615afe9db32998de1b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d56c0338746b4886a65f37c3d6608a5375375c1a53a7ac4e76aff2db28764565589a1d2317b5fd5dee035fbe98404a745db6d662d13bc02bfd6ea97;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab5762c9ab1c84670c28b81f34d59295afafde38e54e8db28d8fad8902d84a0b40bf57fb8d37f0e4c1dc4503a6dc64bbdfe91f0b5dc54bc3d4a710131;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h346b3ecc15ffb3f9d572c403ada057782c7d51ecb5258703715484158703760eced32262eb8effc4ab1a9eb7373546408083bb998646837ebcfacfb3b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32a783e6f753ba6c264db63981d22ec82cc62a58d4acf67feb97a8b5a58906f725a7939a594a6a6eb20ecc98edfaf5ba630f7066f11aa3bae2e7889f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hde571869103583f6d660f19bf91d4f754018a5ecdf2ed5372520be994da5d90a80c5fdd86c2e9812d0ec22c96c2175f93276c4938b1d2f4429ed24d0f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9123d08779dc97daa8f9f3f08b88724295ef5c1fb610740c72b9449fb780687fc1693cfa3380785877251c7b6ac49e70b926063628aafa91991c4a7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha84d2705ff69fb51876bfb9a8be5e8188da527bb2fe753f531ecbe927619947c8fc220c58563a1cfc4b3c7d1c23925e083aa37463c31f0af72bdbdb5a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb68306ae89b73a0ffd52ba7ed55109275bd4f33d851bc297ea97f1d2d5b4d70b6f5b758ae3e7824dcf7dbae44d809d31b294bfd0d8f58ae38c0c8f1dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h85354618c55b96e71e0a93e4f53eed7c86b23b93ff1fad59e7c5935c33357a7ab40bca60195b2239d1650648ff6b944e35352c81b52730b8ee17575cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2d43a3a49d5ab5016360813ba58ceaea7566faaec6cb18c16d90135fc4c4ee8550a45833a83ce411a63a7e7485ee827d948310bc116ffc4572c9bf37;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h696f83b8eaa0d5f59715b48670a434da90665e5d3207e54fc779188d25f0f5882e38f2563bfa712c49e9e09ff786f3c0bc170e6d975d20b558300d9aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1abc10532e55f9e9a651c7017d5e7f667703a74750b08fcdb0800ac0844bc542119b617070c5577b4416edc30f1f03d349e97db329160de259c5bbeb9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he023c499afaadb5d77687989912d64ccbdcd57e499d6da05e3ae694c0604af9316d4a60c2d04009baf94cb9ce89b80ab461de3f2d34a86ff25481d3f8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67f028ae7b7c78bf9d8ddc97b251b42f2a741d48e81cac98aff38240eb3339d1a3b681258ab82edbf8b2f6790168310a4ad6780a6832e5fe3d549053c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h520037299f492b681a16c68288059207570ea79ce3781626cce29457c9fdf02a1054a391e6f15f598e8ac85d9a081b30f2abf976b82a65f664eda7ac3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0d92bce9037eee57e1b3e9f79a8913376399941fc467ef34626575d2ef9fb97811b5521fd3848fcf876a91ab9aa1d640c48983052fe9ff8befb2cb51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc77c3014f6732f043191c876fc815f5e5fafcc41ef1b7673d3f0b0ba4f18ca0799769f3c215120be5dce2f7d257cfb5131e1a510e46e91365790f99b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e04dc81d3bf6081640a7be778f11ab4d69de05daed90560b07c703ae3a07e1fa83fea472557bf3060740d3bc01749abf124190217a4ed3a940980796;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8f7bea87e79b76c4da06799c151a81e1bf3642fd266be4672e5046da4510b876175da6d92a9bb65cf5064a31440f58a81ba9f6c1a01f1cc9de147c272;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d4c6fce0d273780b842b441915e243dea60919d37320e40a3dfd1400f22a4951c57732735a5acc296bff773bdbe25df5d3dc60205a578512f5782ce9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h478abf8e03c8125452895bb47cab5510334d7020a70604d8f6e7e7d746a7fcf49670db92e779af85ce9211e5bdf889ec5a5a2a19420dca52a16c1fa30;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcea0e6480bb0ea38d9bdca07832bdfd3e533dacbd4be413dea66ddde5b145f09fd874f79657de3a8b222e3affdb3f375f54e2418556713ab303a72cc2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3278f509bafe757815f91c3b332eda02dd2ba1f16ab93218832437d017608d6220766805fb73cc601fe7efb75f5185aef54a401d60a3add599a24ee7f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbddddacf7f271ea2c074ee5a06a4767b0c8412f55cefcb3cc64e69d2b0858463257a76f31da89ea8c2f5a4bdef5c17a2c440f16656865e348a992ac55;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9335a0a2994f2f3bf6ffb81cbcd4b49ed0f6940ab76ae0fab369822809e05345cdef166a2a0581cb57f3024ef527e90ba7ef5fb7d0710bdc4f0876ab6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e20e38f1ac80f7d76b4eb89498abb0517cb7cf076d1a83babf433bc0d52160dd9eb99183fe6b980f2e31772d92093aa041dd005836580a50b26cc92b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha879782da08b7160b372262a059c7808a5bb37ae784842778de92416e03c6a2fb0451a97736e809e12f4a65da9cb26a54d475f2007bd473b4454387eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ca4deca13c24f7a5bb5b7c9df3a4202268705c2659b6833b50911741fc3e085ab840d3a3e18e01c7ed823494d136f77e50e65fa7dcb9ed80f46b6fb0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd1190eb6b6beef2c087aa47da772bdee6eeb05847dcaffb6d87aa916c42a4b9f6c6538e27b232e182952cab7d5c5e802b540cb0a18d2f797cf2c1b11;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef6b7cf695e93e13a9b77ffb560b78368ff56ee4259285bfa643eefca9d2d9515337385737ad5189f400c2014e7cb4194990efb91112215f53a53d3bf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d6dc377b3b1b194dffcb4875eeb15e0c42d6fa91329776515d10c1ba8ce0cf0f1be2b6c2553ff674b1c444609a4a6c50a54f3327e7654d5dbc4e5bd2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3401457e99da7b344da364e9865559b255e81aaad10efd590cc6239c7e649878f2e6b75fd90f7e4fe01c2a2f4b39043b052ac6e4409d394d93cec9e76;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5744e085a8f552039a8011bc146ba88393db22e98fd9a1f47e6a7f608b81776910a452dde800cfd13c86835a6736f8eda2c6a22baca839749bc17770e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h304446d7b399673fe55987410d048aa95765993fbd5b28e4df6ba055aee37c19bb70b0a89394c4e692fa2f1f277834c2c3fdb2d17e3fab5b49d22542a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8f498d7a2c58a774fa1a8d15569020c2566894d3ef66a932db8266b31341ba45c4fc6c1c2144e759b59957c9b322c004a857383b3e94825878bf9f3e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h388c32becb0cdae7441ef78ed12705e7b5089f0ddbb2be3873dff192effc86fc821685d417111816cc69019f88e009c660c98326b93178417cbe455e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h997961729f98b243a3982c1ddf13b66866e4c7647e626bf5323d21dc1eaeb198144c9addb4a8878c9af14fb262952b307c795655d0a19079abc9e907d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ef5a48efbe40e0257b71c55793e709658b99e5bb9f460f62fb1fedc3389486958d1896dcb1648f9c61bcb446fed72e18a5d85d98e9c1438247e4e7cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a11dc1351a480d3cd2684b210a8dabe2e48d7104ad1352479d44a3a1ce795cfd7d3caafad860ac6ef345d25e103974a2e7627af2520c83dfaf2f31a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ba28dd05184997d1796b010d95413869cb5c9d87f92f06bad074bba998f430565f75f3f4af45c771d84d92dbc8e2060a253d54cc823e0032dbc7c715;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0cb9284b72bf462d6dbacbc22605979a478715c3cb9d94c66ce7bfe308ccb84422a54d63a64799c3909e7a755520975509f3b8e268aa5d44ea6ab07a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ff7593b8e6ac876eeb74227776fc264b7227ec4cdc8c6949879e2d3c329cd38bed6a04bbd13e0bf05e08fa5760e979f3135d8b643c4af0b9fb20606e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65c7a5651ec76d07d1542363cfa5faf9e962383e4ba694b406b4c0398909dbb81a2d7ad8ba2173c1229e97da6d5c662e6ec31e4ffd77467538a210045;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3712ee0550c2b9f52f5da0ead738e8067cffeaa364d3d594d732bccebb7d634d458a2763cfcd27059c94b424d101c1b90479413bfb6cd0a51fbca4cd2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3445902aec29b9684401828143b072ee7d4b9a68aa9714b4d705f7f7ce78462581a7d6362372f61356ec2d9742e5cc19ca8953bdec4f7d4c9c2a5d027;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15b069123b55af6b278c690705d41a4b787a28bec23bb5de19f76f566500ee36bb472d33bdf22643900ee3a0aa351bdbfb9ea8a5965218a530cde6b0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ba197d3a074d50854605f7ae52013751058f09013a6955b136ed56069d32f35067626d6a31f763a531b61822e2a8141e2fbf51d0b3e1518854e1042;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2869d27bf9ef5e1fb78b5a54f87e014b1404c048cae6e59779d8c29e6ca7b48fa6f7eab218af04687c416275542f0d65c177c04ea76859df12e86b188;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a40f6f3675ebdb555da157a8491b03dbb9406c8982baac1a3d8a2b869f2482d36123194258b87deaee62ab8eb53406f57e29e26554d86ea2b34ee88f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e0093f5a5d6d293dbb83e7538a8833ef6fb22ed9a102eae97babb40f7dcdd09b07c855eed45c0326b69061c3d5d6c33d1e941710f85fa5179d129483;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd42738c0b3316297e574e76c36ae2d149c51fce5e71095da3df1211692c382190b4dd975b538be37b4e15a57604a619504ff0757ad0ebd67cbd649e24;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h375f2b583c5340b6765ccc4db451572fba31c1c2072fe877e499b438d2af43d971383efc251b62374d2e04d3cdb362020f5c2dcfb56827a769929419f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91638de5c0ef2e7792cd9c625bee806e7eb18cbda0111ba72b7aeea152d55f84e404d25f6008620bc78eb211679c9e24f31750a389a99ba81b7215f36;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d18be8456b60ba1ea0589ec37b5743b59a19652e4074397c903781809be8102c4198046e1e1714950e928cb3df23cfac048103551aac7abf455c5ced;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf43f5625fa6a405472377d7f1f235fd80e2ae004093fb6110aa0b8925a3cfd4b0949e3c581da4272c8ba6252a2dfed83fca668814603653c0744d65e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f2ca78ba3ae600d657b13c0e8d85eff47b397995ac8c29cd41473a6fb7b308c017660a9ccc6764deca5832dd21aafc53e892dca5770848b4254eae5a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he52686964f00232dc2b3c0a6507c4a1868f2aa153ed0139405a3dc36ab25692f58bdcc7c5a0d58e0e7d65f7d9a9a5bb5f53b95d08bbc5dd2ed5b13a7b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21800cebdc13f271080a20e59298ebf97057e36c5b59434640ece0c368535d38f789c1745c7778298a4fe92d4ab3eaaf322e335c2bc79f41a6bfc40d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f08051bbaea2be4335deeda64b11b47396abf759e589e497b1f7680dd96f538d37d77f3d0166d81da3ec1bdf4c0321b2d8fe9b15114d087add9ced5b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he54eacae0c3eedd95f2501a90b3a91103f2bc653b0fe50b55d44c56cbdf30adc20ac54b4c324d3bec30d9fb9d2e3cdbfa3d0dcd982feaea89d9998890;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd32153e4e807046ccdd1312ab9ae48bd7b6dd84b24adc6bd309d8c7db62fb5636ffd4db121a9c7071632bfbdce498d6b6d3b09234195aa22d86c6640a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdabedcd6e295b90519dc9b95ca78adb72cc4710954c50e25eebf48659c5a60b7df1fccb549117839e6494db8295e481545fe9489c8c9c25d70e04a967;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e9e3a538897669b3a38c79fa2296b1cd157c3d5efbf9e853638a8ef3be41e503de985cfaa3a64faf3ece60921a359df64ce3c0ae5538e7be8b5d1067;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1d0cc749aa633c1b88ae24d27974da83ea6527a6e97875db6c77f1d9b5e6a0326eaf818d5cd7e646f05a475ed55d2d82e3c1ac5df41e2ec7f9cf9801;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h322aff1f1ff5e3bd810df5084341b59e78abfde574afd84239dd324072f68af8c60615c7277de29d8bc890cec9abf44168ad989e2c039bfded008df51;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha373802efb27146a7dd1706d3948f4a1ab1de1f757313e85cc4e28b43efa90978464933e3934d13ed7644b1e4a6c00bdd19f400ed0fbbd469c8de168c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9edbfa14c7ba88b3a037c43528597e68fb8651833ff7b65c25a8dca6afe21f1e7fcd56c69ba40dd7520ffcd250f3c6b5a671c856872b76f11eb42f8b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53b83f25ca54017d14c07c54ca2f66b0651d2f0461874c0605fdf00dc05eaaef7c7f1162f6a2b5d2f51dab21be67568f674286e7b1ea8d185109cb0c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h191d780d77d82cc30a3574e4d87b2e73a76bb0dacda05e5713548a6aa3ca5498ad2ae9a215fd68c5cf4ca48aabeacb1f905327ecbd5393f8980d576e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20abff49c9c50047d05fdbae418a76be52e0938fdbc3baa89eac311078a339ea7b2ecaa5bbeb618287516b75a90a567525d75c161a28b264e9a2a7471;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h54612c2eeb3edf85f99b46b5f7bbb04adcff8eae936228cecf5a4c6e9cd289450d1a25233c8b7f93b74da77adedc8e51f7bd5fd1fe37137b26c1723a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha48768ffeaa82ecec62a39e05b2cfe410621ff7ec37b9e46a240be5fa041f0e471bce2f41c1e0798743c8a219160639ef53b630e7ae3bef8fcde79082;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b10f030952e4e0dc192d2c68ddc4e50bd84c05afbf7fc013355c113603007e4cf12fe8bfa6065e6a98cf9f06225bae78c88aab5216a86521cef37560;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h361856d56d61a90b295ade39dbf936803f93661245058736be5cd8f4df04323d72f496e8f89f9cfbec7a519b350f1318e020d46ddb93f95decf8c6e63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95e9287dc9b2ef5d5720ac11ca62922cd298c7faad2a0759618699b432567021e79bd8aebaf9a9dda07a98b9d2aee97b9e8fdafaf68b7b0d5632c413e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb96c6713517958ff111527b154032ca06df935faf5034653d8a72c626d4d1e5d0012265f689d9343925e000f8e0b4e256dba8797e0a005a9e84a7187b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfbf3db6a8e3b575b01c39c80ff7fa67e42948415f7074b47fa940a545d0868c4492d8f68be9b6f582bf6d52fe481b62e774ef1ab4c6b8abb1f3556b03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b9832f67cb330f7892581b4d23567f7640d6fef3c471a0ab64c66682439a6a23d88ae3559947ae5143d246f7c780721da3d9a542f4d5dcac5d6a335f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf87bd8ab446a8859116aa92189f27bd1f73f67e4df56d4e021ff2568a9ae6e7d749f7966d503e4b57ac8358ee0e4ad4b2e2f1361f35a84c0c920d7ef6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49a09250cf21e11f57c5cb4f2b50c4e8b4df4b68a6a34c7fa0b21243d179bd1bdad29cdedf4990871dcb3c21409f778ffa297bbe358651587e9411540;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5dde0c15f34e44f40006c40019995af992c0a9f22b214c56935e3b0580e52e61646c31353e170fc07cf9dcbdfd7a62b84dbbc70f825ca492425483363;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3abc9df4aae72787fb1e80843891088009d2759b1fc41d22d6c4acb7e7f06aa98db3fcced7727cd1c99bdb2fe754fd959858db88ba4a0290ff787bbe7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb9cd8664ff220455340ba67510e71a3ed61ee7579493c320c68d0d67f3c7ee18eda81dbc5e69cdab20d910809f835bf3aa0de2d7004f0d2b98f5109dd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4013b9b4258289849a93fe5307a3d7e00216d2571e070db7d9ec8c9309ffd60d71e1ea756acfab750795a7bb6c1d579d49ebb689ef143b368de9dd653;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa7bd45880df0c92945fe4000ff131291f9df2b89d70b292edecbe14e4887380ef38f4b2cea99fc8b637ade070b3b6c0a93fa42480add7099a9d54705;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc08f241282aa7ea2e390dc36e1e64574b5f886e0777b17997181a49f5f7342a80ebeaa294f516e3b93a3308c19a5a13934889d1476b7de48da4d64442;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc872e8ec9a3bb1272e2f0b344821bae1325e199c9df7d187e96074930e4fae7a32d1d472ef3716a847fdc94f319c3d699c25127bf803f3bdd9296645f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba861b26b59ffd8e5004f0cb1116d1c4ea4d432385bf93d7b97fcc3043df8f3c6c95e2e8baae0fff386823cad799f420e33f00dd905eeae073567a501;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb423d814150673d4a9dcd21dddaf727ddf0c7af196467baec06a2f64f5ee932623ec318f5cac43f3a597a018d52a72333d10a77fbec9ace244afb5da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha1ac882e2f806d095395b829f833195123042eaddd276b01764b28f4344a0f4c9226968a59ab2d073298887b18660752d014a9033f8eee51d8242a82f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26cb38429054108936d992e5fafdd7e3eb2734d6bd7c22e2851d27ea3ba7ff20ee8061ea6a515a703e4255b83153b3e34c31bb8fb2de46a55419e5bfe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h850c5ebbb26f21135069be4b21da1f5ff01cc482736147f7593867d29f7f2e236075aab0ad16d7c2634235d8ee35034041b4a8d3f98a78d97f4abd871;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58be42a2ba1075bdd2a6cbf960088be7af65721e0bfb4ce38e4e89b842205d598099356ccb2d84b525960fe5aed3c38372a98ea8208fcb85c54aa1c6e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25967c6b59a1a675cc0ba7f3f75262d07fec3e8734be979c708c7db2e8b5a60a7aadefa4dc6817805c5dbda5b55a160ac2c62786cae76334538820fcd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74d3a27c4be10f7c42fc9bdf8233b2caab29ff2f22927b1607c03213397990474e260292fbde78627d9a383e4aa383a1cb0ddc3dc78c18d2e992da010;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2aaaa4a270f449c089ecca793e982e5ca8bb50e7e6318e819bf7f8e9e8b82bbd0fd2c1e5a9246046b5ed8857e6bf79f7fe66837308758feb983cd019;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha60ac1adb812e5d115742f8504dab461035c34617be725f325e184c80a196f6d98dee240f0187711f7e218e14a1467b969c288c1a73dceae49da512cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89541382e1b2918771a83a0939aa74daff273d396c883a04d534559b24e786d9d9d0de5b72ede7c2e2e0e11626630a357154909ab78f3616ef17714d2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2d92d29280d2285c9fdc24c69587ed2f73e2c91b28c31d40b400ae84a2f4e3f053ac62022b1abe7f83d570e9393378ad38740760d71a01b90b98f71d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h617ea019aae93b37ea3bb5bee45ce2c6c6f62bb8e7b100fe3bb6acdb00253d3c83bdc2bc189c3bac8f2205ce2eb191ecf998ef28bd6cd8cdc5757a81c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d84b3e2876123e82455fd1bb708f58489fdf87e3e22e248fbf346c325f54307137ce7376a0e5d0fb84e3fb79d43189ea6dbdd9560f6e0980b2177f59;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha22a32994adb8d1ca22f8899333b5d83d37c0cfa57b86a96e91840eaba34d173fce5acffe7336e26ac2d894db73b24e67ba7a1d5d9f7b1ddbfbfa744e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0d20e99b4b2c62f00f36e74ada448817c1d8f718bbe61d65f12bf09a5ebffd9266fe2a19754af27f67d068dbe61f993aa59a1c43233b39c10fb74d0e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hecbe7f10dc663ad82eadc58538ea2ce6c61a0cfbf8c1bf04b817182943708e2691e1e1b80a3bc5a841f095768a65fb189b344e178d5600f6712ae1f3a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf000b09df661216934ab4676b8b12714953b858e925aa2a2f5847cc99f9b2192f6592481f1edee22bf5ca8c26e516a017d0e287c78bf24ee10d096da3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f48f4a5647d8991d0302ce9aed5be332f291fc47aeaf75c8b0f1f9029a5243f77dd3302fb389878b9674a5a803c0e12143adf226d7f8bd26ba7b41a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcea8f354946d33641b93790457c8b0e2edbb8976711799e050ff1d8f13ff1d74e5396cca2458475bf723e6c789e3019bdbd41571db82657df5ecc430e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e978ed85f339ab93d52ee10d9be8a2561148e274b14f3871ec719f1de610d255c8f1b8166a64453003e83bc2d238b12c4eb85b69667161b6173b482f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebb98eadc5d88a9f8f7110d7aa9a6fbe00f198bed2a77b41729165f2df682034da1a2a507d48683152ac6b8398fc125e5a792be84e953ff5234bd8638;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4c7b57166364300b6779f8d9984530a68153b30ab6660bf83551b7ea32b435d2d48c96ac0040692ea1e6459e4ee10408adbde62ed9a6fb75549045fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49bc8a4bee3206c4036114842d4fac37bdb9f2442052b9cc02cfbc8b2ad622999f231e18a66c2045b896250f0078da5ca4e9fc1d07405f0485a7f755d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6ae9e35c61c49a6346fdd1f9f7b616f1918ce4dd219ddd652034c06c827d0a3254acd1aeca3e51d391f469f47250663db3f019e208fdae2197a0db06;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90eec32e8a9a00feb180d2a9c67a474ce9767cde41511d031eb13e28af878231155f2218d9d45f41be316ebf7786bbc1157c772c9b2ca57de67f67c16;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa19f42d4cbc31e20aeb71d05298a72ffef617e9371dc3d88a014fe3abb56dde5beca0ec04523dd4634bcbf995d5fd158e9ac5809421d74b6d11e1a09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h200a6b1b1798750a16bb968dd1514962dd8f50463c141c7b5434263e9f85e761542e334b70c2aa87f12716a5aa4cd129bf9e944a2d7aa2b06d03f1215;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b543f85f39e717a47fbabf91ca13103f34024b1fa871a211db912aab8f18a7edc30b0fdc1c8a1bc4b1cbbd3545c2faa56e6997dfed5b51d6560238d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h753ae24fa27e65f10e5421fcfeb75a108c922ce3af6e11d483f716a962c81b8375949a295fa7a1d70a6c78da562bf42f05ecbe6aa006937c56dc3f21c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d5f1e4254e3049b80633bcedd2cda7f37e88b753cd1562327aa7a107320efbedf0154a47b7e9f895cb1ff170d7194ba8194d4c6d07548d8a2774817a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd9979e350b2465f4dcb1868de40bf2e3e297342a340129fa6488a8ad512897dab254a90b7db5c701df8da699b955a278a01e1ec239fa77f57a59f6f46;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd14793e2effea21313a8e01ce1d7024d47a4a1685d7e5fc3329b747213b4f89d5809de71050adfc38e983b7538347e73ee7428a28645a0aec36e071f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5e08f53c0e9735822df22e2537cafe1c93ebf508002292df27e8f361ffc92d38baf0948a42e7ffa254cd006fe91beb4c2f9e12234836ae3019cdcbf2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h46707fea601b6a0f8cd1d7d2304ef3654d7e6dd9831196bfed107aff29d3d42efa81eb51dbe149dbf6862e379854397db4eeacfe7d8a4a02467c38391;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d9145659177503d7d945c0018b70913163e0ee9847a2259b8064dee7cad826a57da3959f47cf8caf22c6b03f67ed5fcb130c7e9ad00ffd9fd7ee68dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56072ba4b31eafb62e2a193da33d39e57a5ca7fe71af40224b8ebdb8bc24ef227f044439c0c4e6b5064b7e07302f68c14be746f64fc861b1cd3f7890b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc22d7fc7f7bb94a73cc057edb2a16f634551d4def04963b0134a84c74313199d6cd9526065b627556d3bddee780d4fce0171ebac81712ccd3c8a32c80;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84047ce9c0be86980976b8bfca0b32efdd849e156ab0d2a5a9342bf9b56344970ca50134926c56584366682b240e9721fd572a0d20262ce9ed755255c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h90cfd68095b31bc169e92bd48ff2feca5ce60a7c608d05aa8adc20708e561189e8506e0b415f3b1de1e0854d7549447de3e6758ca364b55113df519be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h50c7c9ae4bd08defa31d1c7905ab216e63d892d66214666c5eb8da918407db3e28feeb915ad90da8d32ac1304e795618314021a5889732f721869c5b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6bb8778587ab4f3b313ba10db6b869b1fa924834e09b6aa95b39cc214d3f03d049d477aaf43640558be43f33d5d072b1e1d428aff06d18e5dc1626a43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e97aa891daff64c8ec52f1faff559b8ad33572325d3616654e2af34ce685c9e43d06fc1f26c50d0bf72d5b4e1414b79d3f07bdfe2798aeb1d6fbd8c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he701c21f03f4b02eb85d03030a960b6e141693a087f9e4c14b1ab85128639af4e94e25559169c8cbff40a7967bd84d808b04d8d45e4023f52b4b7e293;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67f153d95c845961d372defda9b94fcc3c66d0d6604a2392700b9e8f7c2415555861441752c2c4380d0cce704bb6c68fdbde119dfcf37b1dcaefde1db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6867b0ba8b5902ffbe639c4f99f059ebb5dffda47e3c46452d2235d3318004826af22fb39535ba4e1002f1b27f33f8c089e966d1ff60a3dbf895fedfb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0fce0cbf8f3ce425104edb14de1d0032d7bb7dd46247496b6d68f17ea6bb0c9502aec654314ac2ac51ebc0e094ce4d834aaf6553b9abe1237ca973ca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0b2dd699db938bede128eae6f4dc17184b5eecf05262d719f86cf85e0e29406b2801f52f8e55d37323fb779f0bb07b30d4b371568356ec2a6acb1010;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h10d92189fbe22bcf2702455bdf90560e505e3a01896e0707f115deba4505be448d667278ff928a4bf61e913e4366556ecd538c249655010722a493008;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h717dc2384b6933cc0f0402dfcff7aea2c54fdbfeba46d2ee7a226fc681e97f35bef35fcdebbeabceb44584e9e9151d7fb0e05d30de073d321f47691be;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h902dfb0f8c48c1fa0edd92d531139dbd6d82e4241a83acce39646e07a51190615db6053e5402ac756f9da55dc61940c7a6be3a14a29ed58ad5cb3ce3c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he82d0411f52e777c11ffdb3e20ebb66e815d6bc74da8b1f3e49edd98c0f24a978e1f252615ffa0745d49d473a0b2dec9ba337e0fd9d201135d3a7be37;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88b4629da0a57b4bf2d690e1bd1bd5756213aaf8085192449de30d5e7d233255383289429fe1e80359bbc3153d85290c8b2d8ed034d85c7e33302ebee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfeb509bd71a892b5275d230ce78a38cf201e6060aa43c6f3528fc31b33be66007b34a5b6bbb7f5eaa7e797610b526bfb7f344a2e72918dd2fb637f38e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he011ab4607fe96e3c37bf4a3b68cc8753420b11da6d88fac3935f64868c8fd61fc2ef60db1689d37900d44f9d9c2556870c5482ae75e8f7d1b88d7cc9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heef9dc31d8abe2ee675c9dd2040681f12a36b86f24815a87b5755ed23310f446a438f3a5a8233e49772e5ff7499f199d94dcb183f841a32150d941a9e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc20557d2875747cefcbc7b66d1fd58b7411ceb71e52857d77095b7882c889beb4c784944afd1f39915c0a93d375a55edbbfb2132bd01bb20e20280765;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e3663eff15b5d6036fffeac9c4a96640879e512cbc968f175852f4590766227c08d6c3008fc3d7f6aaf403446ca7d933122a59967ca332658ee819b4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa788941f5df578393d7d8f2273310de7e4533bf2fdaa6f77813a12aa65cc149ed8c8fcae510a02f3ed0e6443fb08b2d1780d7569a065fc0ee1644db6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29308258f35658a265253e31cb32be9c71881e940fadf6d434b11d737450e38319304ba419581c5a1a3d74ed0c11494aa957558e8fc48b6740e1ce4b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6b5ba95338f81eb0a806297e9ba90df53cd21960efe6ded843a33fe73e32cac70eeaec5ea435291c20de7c9e9f5a79aee96091ce7f014a313bf60a69;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19cd4d1828ea13db5e239f754fa32076838a54cae5913491a8ab75a6a3192c089347c4efaece4f53f652db0ff98154bcd5538291bb0046f94fde455a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h679dc18bc4309fc15a60d10308c9b06ea903a52820792c1d8589db51c27cbdd2d3076706f7465a282f3959ddea35950d7e7fab46a512e97ed6b166a42;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79fea7b0d851456196272044a07fc4fe90cadbb84ed2d6504405537a1f3890426e9974f1a9c7d0e999c5c10b19e384423c5716bafadc4d67476400127;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he805b6f30dab25dec5bea163b737df3ce735eacd4ccfec747dd5b6233c3bacab0ce8e12b10f412ecaf83e825381e1626913bd808e1cd43337651566e4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h397c0adc92203b314a15864f377430aec625eecca7b8064619f7cc9a66371005c7ca4c1375fdf33de2aeb239f08dc6ba1a42560abd679caf4c8aed421;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8cd63921e8561a3f92db2ab60ac67a80f5e83f3fb3ea2d5c7faa740c081adf2fe14f6b46ec70c8376dd31764142fbb418401043012ce1d9639fd3fbb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2f6b22716a3e95d1c29c8e0a41570fd01c720925736ad5662b3b91e0c315e9ed955db9478da32f32b5c6f8c3001154ba35175318f0a59bae01b7d91b7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3536c664f4f9b57150dc09d7d1a273b86449fcff36e4ae43578abb43a95fc6486db41cb37358d86ecf6a73a505836c1bc50b7a6d6411c34c79826de89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd2b683fa1cfe1d91bf37e9270c55b8deab80782713c46b12113c1513c987fadc281f7505bcdb77dcb227ad106df845e71cc4d1ab2dc648e47b91629e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ac4d2af30d0f53b2d20e4a2ff78ca153d2941504346379950ea1d8134fc9556b94000c34e3ef7c231827048ab852d3437c012a957fc74cd87cbb39f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf14d163d8a3849894cebab11171987b98e7dcbed8d20d2da7788f8fa69e2f8f7178c0f6a27b1430e58b84c4fbf1e22a5e5c1feadedcce9bbcee4f379c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab164ff9095de6082e00296200aabf11b66ae2a96786a23835a2a16fc4682ce20406a0845c80c7d105bf62915c9d62e2fa6811fe72a3eb5e9da1157bd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17b6d0298ab86eefd05f2910533f44d9038633e3c658bf885db953d5169399ae4fe5789b5baa3c5df0a4378803766ebdd135b3125806f455cd1183554;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d7258e62c50d668f9a29260b6cae593827783349d3a6d077e888d245954f982ff7ca50fea541ba5dc7746c47580c8663041fe1a04b3943a340a5d628;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0e9436b01d5e9b4b6e42c428db3fd08a4a6cd8294a983c7a86da165eb652ed34a2cb25232f74784e0d2a5969b0265ca997be384baf1961853147ae99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha14016e0e31a86f08b86043b57bb60defe368edd0d8c4682b87c0f1a19f1da85ec818f5b495834ce76633b27eec81d9a749fec5c66e372036f618a5ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a1f7e26ce55343d336af5539d7429d62fe28814bf927f69c5a78803fcec11f1384491734ceb98f08e44d87554194ad09206e2fdca0af62c35ecc9c8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d8eb970eec4d780e76301709885a5a07809d3dc71e14329b77eb6fd163c349d4d0a802d2e835da3340fefa93482444befcb5fc3e75a99e84b6386b43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ce714a73357a0472e131b27c6ad91c7312ee9b4c944848c08a942f4f8e6b80da74fb203c788eecb211eb751d21f2bc2e2fcc7b7c42abbd5029d804e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9dd02e62f5e6bba3176f6249685e584efdb2546cf0a8ec3977b3de960136c9cb4b38cfff20ee71bffe6696cf79e715ea51473dd59420fb84914e0f42c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6ddc58f342a82bbaaed6217a3527b94471bb5cc7661cf930e31c131ec180651027195bb6b9a95798a7405f2bf0da4d89fb71573c9ee1a693afed2fbc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h34170357f080f218086098e6f2933aee1535608c19fc0d5f71e9590e26495573ce9abae15a2c9a4eb8197802aef93341facc74d6c35c313e9f24a2e67;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h293a0501901ae2a97ac0880c6ce85f8bab2d670830398d9bf3febe7b231cd5ccf64f64c5074a060c8488f6e29829ca4afeb915f9625e78692e6267001;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b09987fe33db70f83dfe2f22d3131f536343b11d46fc1af0ac49625b4af6c5d3672e5b36688a951ad936093e7cd958685780f962c7d98aac38d91dda;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11182a3e43762ebc1bb586acbdf59c12e55f70f57e56827e33c95cdcd0637ada18206499a13473768d89754ae488b84199b78f76defddbee7f165e38f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h427e73ea8c227d5747ebb2d98eb2e4e188208ad75ca307545fccaad293183c7f1597c3ccbd92e4ee8bcac3a4017e72ad5d9b5fd17c2c53fc52aa81d8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62bbba6144ea5abf0a9277ec6c5b00ce3aa581dbef17b36be82be3712fcd93d997c951cdfa2e9cd8933ba1ba9321e8941c0b844cce24b99f61df5fdb0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45a5b4476b8091a7a1f04bee286f8f83ee030ab50c2837ad08889cf3fe6fb8856fc323d6f5e24c799a3e261aa5a06a4a58f15eb5dbbd6f07e006bd433;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h941c7f8825093f137b7d4cd1723369d8ecdac07dbe60415351106230c21e32d7b6456db713205a683e2511c6903d4f3209a8f7682c0c0c33d9ecc8941;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55a0b59a41f72a273bbf94cc3f8870424c1f8394a0eb7279c5ce5b16572eb97f9be2a53e7cdada99c2fafdd15195c3818a9cffe9564414504a32eca73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h408a28b76ba5181b22c201ceec11bf5d608844e422082c2e2510029203858a95f3a367281886e52fdecacf800396b148f78555b7cd37b003f257cfbbf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h455209d4139b0541a55500442e3a17a001b3b7a629edd5627cece828c3db02014b38b3967ce0e95b60a442f471d2e4799b9a6eada2456684f299138d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5134cb96406e139d6029c4d777e58b4aea7d556c6ce78a1f765682a0e07dcdc38333c71ac85e006007e6df64cbb12de99607ac32c2ceecb6dfbac4d13;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h728e56e6098654e6d9c23ba3d43d028208373d118d1498cf835d09d6a54f9c2b1d87dfeb8a04c97846dfbc5b5db4f981ab2ab7a8df41f8844b8b4aa30;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc5776095f85f4e69ebf31340f1a24aedf0256bb2c08be4353fdface19d94625a0d498c7429932d2d152bb1ba7d3e87ffa1511b38b7a47e3c27de7b15;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h574d37ccb97f6da54624419b4bc9b8d647542501e3264fb5eb799aed3687ba14664302ccd1f958d22512645b770af75f134e2ce26b520d03236a5049f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75e02b62814e88e7aa9da84031951aec7fc237868000c3f214fb406a1724b558f89a71ae4bcbccae45c47cb19c3a32b25cbb937dfa8d348f89658af61;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f51e9f1608789b85b4eb113c01efad157c6a7709d63b3230cbd303e134745ebe962431b2fa112436938d38b147ade224db259d3ff9aa5bfa29d20f2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61e4ba44e39f5c8b68a64ac43299643b66b73d415503574df1abb49f2ec8dc9d994af13bf07522c8c9743b2a9358ee5ac13c906616d5010a1e1603155;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77b1c5ed9e710dc55f9e9e3f165aa0c104e66ca29bee9347068f2a88c75a5886f4237f9e6211d8bb743766603cee6f62f4a476af4f803dc37c222d3f0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbfdc30b4affc94e7193ebd893dac0b14409b0c61e52f5b800d2790b3b086452cdb5f530933fab6f7028de1f12e0dc2119c6dba0e69f3ac0aee349edf1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13e54c651918eae4275a4196bdf38927448aaf38b51a9d21f92f15a2979f75b483baae4a89c0dd50595435fa78e87475926c40c2e3f53ff46dd5e226;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h58bf08b050cad139c472ca28dcdb06a9ea48e2396541423b8f0d962a233960448a47951db56b739dd460491d37fcb2d37be5bbd95559e2f7bb0ffb61;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf3a6b1b05a6e5b2cd651f5e7e092877d89ad36ecb16263cd5d644f52d3a1139fd53747389a133049fe6178d32b4500b494afe82ebb77576a0c21bd05e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h136c26b6285a7fe60d7569932b794eb0212cf260ee66416670702fa9f394fec73a37c647719eb7b23e55545d63515f117bc5606bb225f93968fbd3792;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h975540537998866af6216606d260f55d36be39acf0749395512628586488d0e5e10f3fc7d3700a2038566e62729a24b945b46e5458b0ab689026a3af5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4c6937b841c33a9735c48aeb0de5f0f4158f1220f02107d826062f6b6d3a98d3d88d693c073451c38341bf98739570ffadb56bcaf7c0222b562b35aec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd511b26dbbc8df7e63c243986f7ed1cd6aaab2a73d78e1e947a68b01d5745ea4ea50e68db604234d343a927ba8de00029ffbb796fc049507f24edda09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49fade0d87e354a8fcff5197c31810794048d887e28c00b70f9e3329314b583c6f43984d48c8d5ecb6514922d996e8351d84fde56bb98aeb46929905e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f72fc3a9b4bf7b8c1928f52d758d7e7bd3638ba3c6c75c0426fdcdc54bd186f450c18c3e5569dc78880225c12747aaf5d6ce151a1993674770887567;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcb9f614dbc81666a30e14162c55e95276a267a7a9dfbed0322ca062a369f9bde640a081cd5ddff426ac5744e536f333005f3958ed8ec69c967d0ab08b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcfea4881e789a6d0388c1d532c4b56dcf0cc98809c0871eefd16b739824dfaee748405465036097faf3736253279eea89a5661f1d9791e88823fd66fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0c474ee9ce0aa0ae5072a92c7f02cc36cd87368093c0daa1cb04ec76ff40614dd7174b1e3492b8c1c6693f244d038804ebab8d91a1319d440c93810f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3726a07414c17c6cc7139d2794f4982e06a907e9fb20e1c59a238d1ff9f5dd7edaa08a6b0c0cf11057a3966642793b35703aeb22957402fda4230572;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ae1e20d0efa1703b179ea8e153774fd9bc86f82d855f1054c5a80f1b78d73c8e7669fe1e1aa34df93cb31f1a278e9b9f3e3e6b3c195c184791c0b4c6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66796a7803cd589801bab84a793ce29aecd0d30ff163ecdf5fc23325772bbb338685a460947d6bae7fe2845ec0eca2f2511d3f44dff08b20e3f6df708;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he94fd8fbbd6ba95fec679f1216f13723250d1ffd1ea7a6892e75f09f24addc659eeeb078b7ad15b14537d2acbe9b1c07a4021aa553ff4fc12bbcf2c63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49a6f284e5a5006efc5c17d7f178c9afdc9975a2a76681fa8016771accc466a2be66b27563ee049babe6659e3e7708c1810bbac5be2dd0c42ba09fdc2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h91981882efeebabf75334d0eb11f4467288c6b7afc1ebc6f7ea1bdd314deffa3fccd7d118b76f21c54c2d6926b2466e5127975435ea320865deebe068;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59a2b5c5029df564b482a55f3bdadb8e091ae1b989a8002a6549a549ffc5afe425021c8ee8f6087175447f85fdaf614b401440ff703fb8cd87d5aec15;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8e1ba73cd127977a52eebd2953889573277740035690c73bae6a26e00538b670fa9ff7f085a69544c5bb98fc76d03c39e5b35cbbf547ce462c086e58;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36e5a60601636766fbb6a3935355b9583387d89c4df4a23728b4a3823f3e60b28eb13b80c154b0ae2ec7367a025d52e3fd5e048a04031ed71cf4e1235;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99c90c093719e5199b88bc24f16aed79143622f2499f770d334e0b822004af19e215864a049ec5ce542ccefcb630dadea26db3dff940b1f37c1bd3ff7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5002980908b638ae9d7794a9a929f07bf8ba8c8fe724f5e1b9ea4b917d162dcde70aefb578d37bb2e935296bf1831674e6ae02a60b4f793c2b72887d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d512ae6faaf0ce884ddbd2654df71cfa89efd304a44733565cc910accae8bad00f6194aee4f0a8b7d92f807958ee50d38493ce66622a5986747b6bbc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd491bfad74d6077dfe802881ed15bc5fe5140c7489c959a7531dd366232d0aa9cd0e6913a5a80a754576934ea6021586396c89644327c9e71ac571c99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ba1685ee4efe77f609cff2c26088c644958afd4de57cfca9a7f0e3925597e97c7bb3cf9b76f9178f355d7006268c3438be6e8e3a3353800d12e9098c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h787e8f4128407dad74784e6480dc01a87c9468f86b6962da7b0a4e4807206e72823e0d926efee6d0fe6405e94245e4a9e35f467985d309d570df3c5e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f2717bc730ba873706ac585ee915b4228d346513f4c8b739c17f4da75d11d0289c4477292a74e8efc93cab1bed1bc5c88edce75c9a7a0edcc0908e3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf51df69e7e3dd447c4de0cd8b0cae254cda4132a5a36c3b49afe69964869227e85ed081cd9a41b0c91ce2e6d665731b6cb2a3ca17e93ba981f3ef682d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b9d4c35406880be2d639095fc26f76b786205b78905fd665cb18a3303859a27f0d98b06d9eda8fd9f18d34e250a11523a9af4494975a0947102d7801;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36012db794985a2653a0da60a717417e334951d599bdf70655fc00a7ae141148ecc2b89fd22a2901d559b6d6d101f66e874cc8634644881ef8f6c14a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e5b8fe3f92b9a88129f039e59c61009a8f1eb8cc2834805d5f212a75ac9203b54b0a53958978aa9b92012479ebf12ac83cf7df799d796a99c7f594d4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99080b3a5915fe15420c630fa255a5d0bdce807e31a6bdf8deb382ddd453ce31e17dae275beed8237f93b7af8c71da8ccf1ce5ca3aeb76fede594b7ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74637e66909f40147ad17ea4a913cf361a7f20f708d6d3f8c2fe948011402bcc44a607f6ce85f3ebd7f3317e1216503f09cb3ec7eaf06ba7f5ed91253;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb29d90049b685814a5f755e0675030297544a9d271452771d6b32b81ca938a2ad8148fda8212437326a732c2fe2d2e30bd5f1ff35f5a7166ac08563fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4488b769543329204848d19279ae596ed223f379e0a4b1f2b472777d3790b0342defc402ecd886e842d687dfc20dad6e8a9e425445e3d8365a90904ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2184cf2cd7ffe0c20dc4043d456996d4f0d6319405299d4382bb82a091344314d7d8d00c9fcc4700c137ff3dbad68b41d4175db2f16421933cf7763bc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1dcf8aa6f0102b78fbfb4185d2fea631b0f5a1897e978ba88952c1532380182bcf97c2273cfb3f31fc8b09a13a269a1063d6e9e0e4cce3fac81492ac2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h74240f5bdc9bc2f77f695496290d782ce89ca9f3e5cab7ef8c24258b592c876a20a9c1f11591b4c7fdffb005fc1d285d87dea303badb008d9748df8b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf0c9b66034ad27a215e418c93c08575e584289b2dc7acdd752a34f3cf1aac6517ab9ed3be47c727d063cd43e73ec3a3e3a6775e20c3c5800572e5c855;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13cd0502fae16dfe53b39ecf29bcb6b54501e72313deae7fd466a8c7b7ec01c874318c06e97ff132176f53f489b433c6586ee9cf5d1f8a06121a1f8b7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15899d700365fbbb9877208aaa3dc4551b69bc0d878d17479f93e83e337f8f009db7ef4a668ad0ed07ea1e32dc0d540530917c0d3e096e7f86c8edf6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h48a2323d91aef39e292c702e5165479fdc46194508a8ec5ccec372bd16b1180c351b7057714f6fc0ef780d1f0a05071a40e1dc512c4b0fdb764e74a71;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4664f3be9eddd3e3a037456dd50e3f6135b363d096c41dd8a5809b2d504cdc6d3ffc194296d009941348706e2d7a61f39a24930afd51671bdbae84467;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb3b6b5c10827b0a1bde1d03551ec9ae64eb62e1546e1ccd7cbc81b8942f1ec18677dbbfd7d1e2e61401a3efa2ddf503e55225706f8dd9afe70a7383dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95e5b2125e7ffde0e7ecee6d17bdff092ddd5a35002f0e6902ba56eeb06e2c5722ded7b28645911283f387812f4f83fb00bbc25993a1e6163ed335b43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95f1b0886bcc846855176425fbbc4c0a943d9ec7bfa2d4179653d42d81314af77d5833df3f6b2f79e81e44b0a1819ffae928e9610fa7f97028462c2e0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf083db3682624450ed3cb9974b5c32cd75d24919f5ff4cc95971d118b02eff32cd224631c1faae30d03f5c5a2372bafc8ee1f2fd7d4528eb64d65c112;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h57f19f537e33344b3e6606756c4fcc1e67e2afa7de189a1fd65d900dc26982a11aa342dbf8cc1a5bea1c1c65d07eac671dc87525833c0338f73b5fc28;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habca43b18480ec91fd63028cf6e0fcb8a8ddae572ef08d8af9cffe9f40c323990ca7b4ff0213708187ba1ae1166e93e8123ba3953f91da4704f8193ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb58a2cbde16d01662e27cab52cbd069b8fac73164f65033c1f1d10360754db31514911d6313b711a6026cdc09483eaa6448dca01208a3ed42480c6e6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hceb1e16464747d8e834795f10ef1c04e9150687ab0413df9d8934d62c0240cc7cd2bce96367abeaef71a0385dd7fc887f6732ab46fef65b90ede86850;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb87981883c42cd92660969f114a08a1d94313c9a296e9e9f062eeacca7ddf654ff990ececf166065c61cabe85ba142001345d033ad2b395b32b2af9a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4327150f42bc32bdcce316999e2947194a81c691e7a0f0a0772473bf5f41b4b3605324b69b61c4f8fc39dd3487ff403674abe1c42757d1d592eb3b7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he57837d27e87f3aef7cbdbda63f21e3fcf74a7a798833f2a40a57c586f26a7dffa95672d0c1475037831d665d681ad12f597393d5e800f32685ccb876;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61e84c2bdb34d1e119ef2718f83173b88e48a19d97cf19d3480422ca8bc026fbc48a2fd50ff1ad3c8b9bb0a34ef65425532e1861a77aa79ddfbc592fe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44fc356b4de3dd241b3735dbeb772286c6dc33f945dc709373d83f2658ea1659f3f7d22cbf2c4c0280ab1ced22f6251e7e40e3a1259e352953940a84d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h540cc0d07b9dc4c5c0605f978d9df1efe3fd95471337900f48fcc60a2b139ba9571dc371e675b1f9dd7c9d85af9e309d08bcf5455b5100bb891db6a74;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h968ea56e515ea899bd2333cdcfb6c6ba884ca601903d57815fbcb9c1be46a474bafa4db21b7ade4a004c1074a944ab4eeaf58f09bc1bc71e8165567ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62ffb24033381cc78b287ac05486de0c3c48a1547c149d4a70dab407b62c54ab22875b7df926f8b8000dfddb11d6b0b26d9026d724e001bca750b2fa2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf5d873b100850688f0d1e7fefd920f1d36c3d4d61d1dad7db433e84222613866af8ec669be250d70af47a89f7ab173a91f61b0b3cbbf97b94b181898b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h27d540d7e92533c5dfb6a666103419e2f7d4afc7abee8dd7732f7defc2ab06c507ab20081952edc94f24b8b26a72c80bc9d61c0c439ff0a33354fe611;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15628fd5fcb86f2b4f4cd97e4fd82a287b018737cfb6294f43db29eb0e27ee8d89a3dc522a6f4376ce7e75876cb4026a488dda58c8f5566a8963d03e4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h486ef5d8f9b7b7c108e61a582d75df1fc5c4e0c12b82f7093a26f54e8c7dc17644c39190fdf6b5e3756264aecb3eac05999cc8fabf13f2fe2c880c71d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83212cb89a918713bdd2f348521b798f5435e071bc9a42671348772619948e79f9b2e1ad76836fa00faa20527adcc99ac40c70303a87f78906a938ab1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e58f0fb297854906069fcc4dbacbad6b6474a1f2a6b77575d16093ae8ca6379d25f8724aebb6dd6740825a126ceb410ab82ee7b6941fb981acd111b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf692f7451075c538764c01dbb186b691caf992911b8600c7aa9050429412eccbbfc87687e2a4b6c3cd82858a1bfbad256498e5c1bf71fa7c5eec05749;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b36f7b10046559185475891fce98dbe74e25b2fc976ecf969faa249c3c7d5c6c4005169718b4f8070b6905c47f39ae717fb4720faf4eaf1ba96a046b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d190e3bfdd986d0aa0fc037ae3b0f77e668f2ee48eb2a24e1890c88cd8d6572c2081efef14d634cc3268f45db7b36e3d78942ed630fc0bd53ebfce54;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf868db6f8e53105c324f9fe472fda705c2dc4d104e9903cd84ea46e09e82e9a7b52d1200077b44ac02adebbd4959156f45ab35ff109696802cbe32d45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h609b269ca952d926cff887b52b330612ee92013e7ebf1518eff1493fe0a53bf9fe3b392cb4028be269a59137a01680967bcfbabfa14b4df51592bcce3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccca2b0457df626bf7a79645d17a4215f75f25a858b2efa3ed482f14769c19b171d5d039e445cc947734e4636525e2603008b7711a01ab0e7b98ac6ab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd235827024e9289ab09fecde4815fc2feb15255e56dd7f61613f9a507bcbef86f763cbff92ed1d1269b7f25d3aade29f04aab7b553cf1f890d9f186d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86bd6b72a4449813940d5272bc0443dc5a284e1c8d631988cfbbcc7279b66b8ab5d1fc019249cabd2e594e153398df87a42c0109e9027a0c644f03eca;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd82cdf880368933b3464e9379752dbb6c5091c655d4fa4bf85fde215196ad38b1204e18e116488f5153f325e99403784e152b9a8f8550b960eb7dedd5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4ffc49704ed2e2de691b0fe72809059883973768c0164c5cdeb0e02e7cdcbd0d100ac953593abe61b13e9015df8687b8c898946fe2b05d0a776358161;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdce08e747d970420ac851b4d14c8292267933c952baf862222b0383a9b5b46bf5997acaeb2fcee1ed44a61daddc319531155b9c788ca28121128ad286;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h434d1d1afcc76dba1d5ba044ad6f7ece8108948ef709527a694663a83b3472d87136729f77f0239b803f0785551488d7e96831c3813dbc58d1165904a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6d4c129ee9e7f6ca419555d21127fcc6b05e0dce1e6934f070b182cb8a32cf8c44be0d5ae88ee6297451dc5a03a8b8486b9b33e29a78a4f9992ec7a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h999941646a4c68e1a8f9ae4383c038bb35ebc806ed455a2bb26bc675b1dd55065f433392841c70cb67f46e234f53c0114ccf9b7581cfc7ee94c036a2c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haffa9e49b9da67fa6a9a46807a87a38aa417a8c8bf83655385a4b87235e078d3911ddf10b88eadf5b7ba19bb465c3573197794f5bee2799d598ce74c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8755b5f2fae984f2abdc6ca1ab6e8131e6a00a56922e7aa7861f5b60b4aa3d89f026a378c7f7675001489eabeccc79d04a4a7f99875db728f5d37d626;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6305f4aa202bf6f91c3d751bfbd02f4e46ad067a9f893615fc28ee2e78cb28ac5b35de40c9819698a045d96c7d1f83010bc50a97360989653c09aa100;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb73fd585e86db227b3227ca80becc52ea42699806b2d384804c8879ce74f4c8d30e83c1786d77e1434d4910dac43d1bdff2a75e46e7e1aaf5a9fad0fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e633e0a43fe16afca773f0533a2d64f58ecb64b45dd4c01f43eff7828bf3d6b12570ea642cbffaa42dab8c4100c75a471ac597f12b4522c2f65cc02f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h411d87cff4076a3a9e18fa8b8799923c6d933c6161e40eb2195e7f4b858ba2214df265888a100a856482769a235e6e9e4fa16aa85c1255e9654ab7f99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f2db8a695197be1c72bd05264e02c403c3dbd55b8a9115833a77bfea349fd0681e48b6e37974fa15f1b506358c531fb5b27d1486afc323ba4a85abd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d16249c6f33827ba16ae25f5cacd5c72c761b53956a5b297c57a499f8f9b8f77cc92be12927cbbc5d8d7e91e29bec6c83f04a519d7d270a26ecb947e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2659423419243bb3c7c39a8c0fc071683963b561291a0ac9aa649940a47fbf29a98cd4a580837a43802510d575a5060e90f9af924ccd0925968a8d00d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62f52441b9668ff5d216353cb006fc05468b388d5ed53c084cde10d22cc12c5a3ec1accb52f807a0d2e9fd5877d5d0a2491c5b9b987f79a8fca93ce67;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7e5a3d742ba0394f84fe84e93d1a315503ca0c445354298fbe9e92110cccf2dc6325d5e199c9d9eb6aa2fb95ed6ac98a4f193496e6ae31f22c77c175;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb693832a4012b453cbff3f66f879190834626ccc6976c7e32698e60bffd0fac2dc8154b07e45719d9cbf34153cd58fb6730e5d70ade756ba20e9fc2ae;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55828255337eba59eb146936a005a9bc6c60e2e85f9dbe9d9c160808771443afdd9c4753c2a1e48e994624446c878db57c9702d1f713635faab701805;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49e7650ebde3f594493694106d3e4271d5417ce6677e9001bca5e6618c9ec629390061a0d8f4b14516e1b90391a86e9dae915110a8518e9343fed8d69;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5854a490530d0e14df6b577c91b3a43f65f161e563c615df59bf9e31dd75f2f22d1fefb8c866790e3b286f29cd616dff7e6d9ffc8d2b57b07551f3a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ceaef8d4dffb2bd3798ede1b95019550f0a1e26712a914790a19625e75b800e3d1943a76f3af8f9ec0f5ccb756b17a96affdb852d5b99ae06709014e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3fdadd60afecf31c00b4fa8ea68177b05832d6ed0f19a75cdd45b4468d50e472e70e4e76a2fcc5ebaa7710ef131c67d73c47a49c667eb3eca76965629;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb822b3460a000f97a9cd40b6ae3b16ea339bb2b8d56c9fc20d94360fffb98b2a6249c0e65bda0e9e6d559a714d12f01085b4590b6d5857d4b3ef59b09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd50d82a26bd460c4b2c38b1d5a4f5e68c7afd09604226657d61c63eee9acaefb03f3773b7d83061d7403cf9e0d9d9bdac46c7e00769daaa1018fd2fd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3d17d5c70a28f71461bb42f98ee3b571aa6034838434d9eae1c0408b49d42575529a6a3ae535fb6f70cb507c8f56c0296e6ac77fca21aec6e4e4293d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1cdcbcc1591f4add5256b65f634cefd4592d251e540d6a6382b9fa1f5591cea62bdefac7722e0a742603472776fba347a05a6381a6a406bc7c1f5cc26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4035711146ae3b213044ef697f1765cf6f0e95c0f306ffcdd3d7c435d8c8d273630b8732300474709e7e3f98ad5c808dd029bcc0e8e39f59eb610f5b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1becaf81a13e6e505113cfaab255726fe3348b3e2f9be717252f2aa10a8e43a7ae380c2e2872aa116d14f3191da617356d020c7989e7f5383fb04c34;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf982e1d630f11cc2c44aec6bb35c9e5412dcfddfbe1cc2cfe3be0a84af78dca2ad18ac09439191cd4560ae76776985cdf184a739b1332c70ad9c07d88;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd3b45922a6b96dda72def0a99d44d915e83d704553fe994cb238729e5fb60891c36033fef77137b2da94664ca4146231f2cdb9ae042075157ba068834;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7614218b0569cb541ca85195a1cb1ed54e08e17768be8a24fbf135902459f1bd0b3f5f57d66f6578f9d95f88fa8ee473f6dc1cffe0eac7f72809692c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3d7fc4da32e99f7c1739719d5e0f95fa5f0e00f0512bd37dcc843e68bb21540ea7730c8837184b506083f25f53344cce3f8e26757215ae297724f8905;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h911279b5889bd508865416f677fb721a93603f22db03c8f16347f6275860a126bf8b21f99711d3bcbc239c24546954b00881577d63f61161080e2ed9b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7f4ac06ac5dd729bfeed060f630dfe763bbd1a0ec51d6b9677bdca47319f79d5cb78164a5e8da1da913633110ff2cb5291b512d0e7facaaf4e03e139c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h854d70bcc14de17632ce9cd2b22e2a658ffa92a4d0c6f9fd4cb81b65a6a44ad5bb4bf6f734dc1a6cc0eefd859185c6b59fa4dd38faa02aab9d6b5400e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92d23f9fc630bb0d786e6243417cc3fd4cb5758d008d34b4b7bfc99e8c7d27cd3fa02b1bb92121745cffa53d2fcfb20839021401f30371b6a74232a72;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had6d43384a15873f4f7bf310d9fb46871bd6761d947b9902256a3d31fd69f677110ebeb6ef848e5b3cfbca2def7a9e1bde8b591157884dea08e69f83a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heaf72ccb860738f455c60127f7eb27a0b4f5f305f8fda9a48ec32c6130c99464eaee78b9cf5f0f2ee6e5dc8ccdb68046bb75cf6b8a33f477158d22cc0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c6ffaf7a2d991cb532e96ba8ca32eb1071741fd5cba5cf982c9f614c95afb80b4b432e522ff125c9600bf0d7b582b0b944e63c8b6eff4fb450fd98d5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51d31231be88568a62986edf386c8e9bff1b65a4e9ddec0244aab28e25ff8d2c8af9e6a3a3202aa4f34f62d5d8164b4b5ff1deb0fc54961973a044050;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6629250108f3d39037b047da12be1f908e7466e77cfb518302960e9126baf0e4a79e42a3540d53287d7a064a504245c08b96cdd9b359cf6c17ba0e48a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9db85b59112edd7e34e7c4fbd5a50d1f71f2c4018a44a17c0c191625cf551c7f116f3cf2e28d276af4df3abd2a675c1600f73b9ebc2bf17abd2653631;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18afae2708c6d913937ce6f44353ff86a999bda9c0713100998e6e7b36ff70b64945d82a639a8207d6ec8c8ae14ffef1df6302d90305a392f335ef262;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b4751fad16cf7a3d04a3df6ae52d9d9890a5a812de9fa499dba2f2b7c773a6a167129ff3a7a75a568b0302a5b562bb274d94b58a96ebe7cea4314472;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he954caaab85a3c79d17f52232df729cde0a41bf37eeda3740f4b2b7b13a955eff7e62d51a36aab59d4fd15e779c8aea8e0a689c701ad3c5686338004b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd921281c3034c4b4d1e03b223a4db097c601c8c74e1cb4ab4750277277ca6caa3d8e7504b6691dd07a649ab7e53429f70e6fbc99a8150ea4df3e2a813;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2e12b0c2fe0bb9a62112f817b8b396702d2018b21ed00149f96974735923c2c23b9fa202b4406739fcc3e7594c761f50a9ed587f3abeaf45e6f8a30b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43c5633a2502c58a5d1459fc893a55b47cdc38c4954602a32b8fc9e3e9339b6456ebb62ae8bb6a6d9f4f8b9b5047a03023f0cc06c7b73239af5e62d85;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6a8060a89eb5cda2c49070f69740ddff46b0b247d423ea9545255eacecb20c90d2d6604555b6e972b5da120c9df87af89fa4ddad5dde558eac23c0f24;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he13349f778fb869d49bf9c4b93a3f4675ed852c18a08a7fea212cbd33911fba681bb99c106b2cfe3a5a97036417ff2ea7d040f9d346bd6994a7a45b5c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73c94778a3416010769de0f95107d827dc2422dd4534508e6384703e19760b1767c0f75bd9d81de0ff8bc8855862a06df688d5368b89de7b2b82bee17;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h420bbc1078c75e9e39e77aca81192a6ba9138bc1a05b68f834efab8218977e3d3021c41b59763a0b5b52b0486227e53045dcaf49ad825fc591a2d55f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha923ec7dc1f4b2a888358b3d40bf652e1918879a87c0d1ec5fcf259445e7d25c5c75457dd1cff0b67eabc81f3caac4a1c8cde28554e61597638d6c6c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e3cf3cd9d96fd607e55ac8a70013d5dbc8a85c14f05166d196a96018fb11d648e19d787c39f95ed08693fa4267f2cc6edbb2e7caa9f418eeb5dacba1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3d23c6b74cf5ae6065e4ac4ce94d9eac0b31f5025b82044c300cf8906d2ba262990b22159895182f5be1f1923f96a13a8cfdb6a29f6af9ff31864fc3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e050f282e806f92a1b968ea562eae9c6842abc72059c1a69575def4d410b2f69d89391a9615abb0b84b8311a5975b9984d5f1b825bd28a644aea8a2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he54e1c60ee1ee2c8a93cfbb6a801906dc14f6ccdde7b62332010b64f3cb1d597970d75f9d3bf09cc9835b3a1f55a2ec318c9fda360c55c959ebaeb10a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8093088cc13a9b31fd1b8f719ce6fb0e1b3f0779362a8d4aa0d6390a192cbba18d959dea7988e1787fafad26b6835cf4268fd8d8174b649cc8609eba3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6daefc188e78fb79bb830fb58ee17f13dff1c1150f1b295c11275225536bf8041d15038646a47e7f4b16052137f099fe718f0f107c32518fd619aeb49;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha4a2bff55867aad3fbf1e412295cf6c589da441983e0a59ce3f7093674f112416e0f64d2c97dae2d61ad13d4ff7cdf86ea377085194561f387b4335e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ad8ac40bba74ad7594adfbc4374549e9dfeb0c6e9bd621390f038d602d313de514463e5f981a46ec3e192a7bf7dbc167bd1f82c7d4a953133fc24fcb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c169a6fb7ef20320436ae29c5339937c04c179b33819808552f2437b19d385ff10ec2bfb20c0acb8e13c487b86be1a011fd00d571f2febb55f4156e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f0a7fba35b105984a6d1a25409f5565fac05faa5cfb6134e7125dcc4467b740cc74a75291e19d338766739069fb3088b0289a861642a483f8341180f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h37700b4856201dc21e9f3b50615346ad63e609d0c22191bd8020611fd8730f065e028889202f1e27542c2bdf43c24523cb28693c22af4d485c0575238;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b9d37377e97e0aab4ea54cd5c3f6b17bf23b44112b0e1652ad0979fc840609cacd481757b34806ee4497e587fb5609d666f561227ad348147676ae45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcaf5635c6914590979a0c7dc2d13c51ef871e24a348dd8e2fcad458041f985d2eee62ef1ee1fef4c4f05ee609dd2d5c21a8992ca7f36b23438bdb9fe9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99f1a022de9950690ee7832912518c48b96ae7f6f633451be509cb760dcbaef983d295f4ad63f3dc9a40db4276790470d11bfa7312974b10a41584557;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ced6c43f7929fa53d4b4e35335dd936497f37f43e8cb5a392c2a7ecdf05784a95da24a77e05a279b94839b140333ac8813154aadea77cb9fd6a10616;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1e86a052f488cdf9d518886a8b8c23281160b66c757ab8d14f816d60c575b3cd811d727e86e2fccfba5b9a5c625ffb1327568454a595c7cf9a2b6db07;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h204f136eadabc71a5b611a2eb91f2a17bcf26f504375e423acc9a00d69bd873cef3e1c70b9cede5d66f8d049b2f61de6d21790fe36a371ec73b95d137;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcaa0b55bd1a1b29cdf634745e315bb637700fd9523f2145928aeb3e5db73a36720314064d8d521e540e3cec821fdc8ffda79ee8b7b0ed10ef1562853b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd899a2cd1c201801a720b5e12727a064d0cbb93d5c630aff9581c54ef816c9068d6a99f1dbbc9e44899e794d5e1221e657003612a6f26aa2a1f68bb8d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h11b8089ce36995c343d20c71d9b298abce2761fb590580be8edc5584db478db63f46f70b3352abfaab003ad3c343bc6078aedc2036dfbf1004e7e7ccd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f0885aacc916375db1a9557e683a48b875667ac0fdbd80b93524b92d37aa8bde561b9e29cfa2c132a2e9123aabdaeb846e0270aaf8dee02b618a58e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2cd62bd1fc559dc3332afcb30a7f49e883ac4860aa9f6aef6396ad0e85c7f05e91f64e93bb9287a8bdc2f097017804faf7611e9ea3316b4edec2ce77c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9e5624a9d0fa1f55711a3de561f9fc556a248bcfb53bad12a246edfb5f82ca23ceffdd3f8c09a386c20edae9e444a9b8f58c003b96af9bc428854da1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7792dec9a029db4a4bce5a612208a9f49d8dd5f2f097acd6f99f9d69800055114153d551a295502d1fb20664658650b5e4ce0a54aa3c230bf2f8f585a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdbfa282911931f3f73be91635303287d62628f1cd1d852ce86738603d8e45d1c8940a31b34bb187fee24f2deb3782d29d18fcc301c60c83013c396bbe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h42b69f4689f77ca95444204155aa114b1bee3d4f4599ce060817d4dcc6c1713778970e7283e8df8cfd6f3a95edcff3f4edbfeaf23cd941831fae1aded;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h63dba9d01033084d1f4e89fc892234ec561b3d642ecb3090f57044feba6c8c1a0e9e42e484a95ffd44d1cdc7cfc50ebbdd49c7b03415e7ebff534c8f3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a9311de7d50e6c4c255717f4b7699a0a62a7d27f50e9ac642ab2430eacfc03cc763d49eac84e97f92289963cbea01d6e44453de8a04773036c26d8ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h16a93640cf4417bba926257287981dbeaaf5effa71a15803418854bd8de1fdb531b3bc31b9a91801b131c70f3e4b702d1e058a1ff84f3a84f1d9e2128;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfead0ad8fe263771ef252c757865bc5948c9cf61e90962329159a299e9150c7f6dba49a542674b8056adc47c465d3e6bd7be424b3953960173690b2eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66733599fa794caaa688f14d045e24f7c0e6fd081997f5e28760f57d0cb3176221ef4092c2049fe6ec1a79af5ad2d48630ac1dcf9a80d4c165928e794;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47495097cd835c4bba4c6d97cf77907310aba8626ed56ee1f1f369a3f3406428c6616350eb6570acbc2e4dbcfce00524150ad50fb832c729cb92dfcd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b4e5e58783af95c2a4403bd38eaf9128a6745e2f70e7dd6c41068e756911c0f1355dea04ad9e3e829fbdd5019e4b52dc69c82f45f7fe5a6b496e86bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h505eca2555f9a51354b776bfa6ac4a68b4bf4defb090526616fcc72da3146ddadc254e23bbf9cb15adea596b930cb955ca2c13315035b7a4b85253123;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hedba36f13f818eb6db3941dc3232b245f94cff3a170e2a896b13051f8fbf09ae4317bfce04e8216cb95d80518ca45c07c18ec1f37124f6872b47a3d4c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28092f9855192792157e0a6f9e5b1dc62b73b072571265d873f4c5bc68728eb102bceed3298940b1b2ae4e613aee00649cac197ec4418ab610c624e9b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9518fbe199d8e2d54f49a259648f553597ecfbd053f6830e7dc230fe2877d885eaf915cdc616880ec01ecdd8b463a94317e27b23524fe05867cb99d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8825fddc92ce18bf94c449260e7990db4be2c1c3611b3533c43755e4449755cfd8d71dd307276c85cf0f8a10f060b702fa42d69c0b56b327dc622b7b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heea4ea7f9e52933a1d2551a1d96a45950a38bd2e94435690dca5bf174b06dbd5578199516f1680bc2a00c71ce32f243a5eddbf125f51ef7ccb9d4853b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49920aa245c01e1125e4a2229f8dcfdd913bea4d07916d23c8d7edc7ea2f07ee55cf4bf9307fc9a61a87ebc6576e9055093c3eed775a2560f966982a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h99c651e11b2bcf3b5c92c190d800a8d33b609104eb2890974ccc8edec1d6008fb1cc03eeb60b3bcacb9e9999afaaf5db4141f7e5d5c1330af8e1d11b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h971a4a002b98b48596dbefbf16c77502944f980869ca9e6675e59b1117324b98f9c06b9f9eee2a697fd14fc6d60378f4c835bcb59e2f25714b2c7c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89728e0716900bad25a96aa6199d7cc5f07a5cd04263097a17e863f7669f475fcff0cde8c88531e3c3ca22cb97f2260dfedeb5c06c02b08389f2cd35a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h614a4b6a7c64e3a1b0b02606c3698484cbf292fa47ccc6f58f7150913c11ed2652dbbdc1a8398621d9fd9c5cfe3fc409c0160b6ed102db17600b05a60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffb2fda84727322e3750ae29c4554822c029a71558a7ef5ebadb56183efd1ffa9993ddaee697bf2831f310c7236581ded85ebf4ff49281f3d14b6f7a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ffdbaf976d7b789edf7356b0d97b2c0624243689a4ed743c7bdd61d740e0af308c02c48094e05b69425f25b08423ae76b01b7e9320683f0c0299fc97;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36bf2c82ac3c9dd3659839839b697b12f5a14fa8e7fd4ddfc00fb77af67a93de572fdc312057a3258b4e1d8179445a7edc5ccd1717fccb50c4a319467;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3720777298bd830f23e9876cd691b9a7b459c3a865fe8e81590b8a1fb799bb9a9dffd37661d7cafa45b9ac268e02e15660dcc087de139a3796179444c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h92dacd338e81e53545a0a3aa806a64c87f06ed7fce3b9e27f8c457ba138eddd76e13037d20a0543a59547979b4acced7f1463d9ec89bb7fc9892b7391;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he2b635e59b01c9dd441b74df1452f19f5281741659af0f031fe31af12b852eac89e3c72616e588bd117c917d6740e7ebdf417a599742c528cddfd7ee4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc00d5a094afd7932cf068e6a2cf88ffbd0b949a972964e211ba5a1917016731f9f0c69d602bd6af242e9375392604639912beed6b2f27fc0a9c1bcebd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haad6fe3dcbb79c879273e556e9e2038be88ceb162f9b961be757d3a9a04da257d59d8c567e0e35a17992df5a3c42df49cadf481a4524dc548adcbacbb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c5e97fc321fdc5f14275058a6763b563cb4ce04a11353ea8975eb84717e6edea79b6ff7c0ec4e2ad7f148310275a7b9c95596760d754c575955d6776;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff79c4340c568d0d9a35a3b0ba82953af6d13d9fb2aa0f099059d999e9363f1b3de8ed1a62d3552bdf7372b39e9435a9ad4e5ebab905daffbdb38adbb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb7d3d36bf9a126100e8721a66aeca811d8d2daa6ccda0bc339871c1983e86e42abd176a14a4adc02fb3395102b563a6ce42430ed7c1b6b5ff4b64e77;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9ace33de9b6d5f2c6c326341b913e5600dffbeb24f3557ad713f4215e8911b3eb716dd3bc9509a050954143be293fb81797dca62424cbfa910caae38;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ad316c9509d6cce6de422a3dbcce26908e40b69eb893ee73fba50c1aa6f8c8ae928f582a151b0c6dbfbddd74ec11b6217c8140e9bcfd00880acc791c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce0c88c3f8dc159f4f4f4443ce2949475d60503a42c5237c5776727c0216dd16a2bb8ffaaa03fd748d791dd1a15c3f8ae10f2607b5efe2e84808af3b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdd32d923fbd67a1ac109e78cee2ad6671a8dfc219fbec751178c6abba86abb301ffee0894461e37454e7730aabc869168922d21ca386a9c6d3eb3a458;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdceeb46643360543ea341edbcab003404d7c9c596040b48852fe9b09aa99674297b2e73ed8aefc813496a1ffc2311c811f2f27e9fe82646fa232a4c64;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4dfa8bd713d2cbaee05f877ee9bee7b834f00f3406bfa86f893bd167117a26e6a23d4698460e34a07d5ce8e70277849c8211dbb2701e37f2aa31ff592;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5b5256259a58601e6dde22c5e8970a172c3797832104658a7d040b364817ba5d5f7960a517540db4eab8c1e6297c993ae7c946f193d1b3ad400b7d8d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hacab6d2cec5e5cc946665eada71c98c45d3f44a0effc95d266352c4f24de10a5da6b4c9fc7e0bee50a7dd496348d363becdcd3718100b9f0fd9ed1449;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb0092811f2d3c27ce403828c2c38da508d5eeca547d09a4cb7049ef8d04066e9b29cd31836fd0c9fee31194b478876b74c27e3d04243dd8c5ced68bf6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbbcef8850e9f86a90905e6bc1abc88a6f0fa9c14bda244b0abc126eeed304b043e2aea4c3ff26ccd49149c0fa0a1e2cff92c057819f4f3b5a4118057;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5cb05da77fa55a769d658de8e7382be6cbbd5777522dc9240386e8229097e1acbe2ad7dfc73ea65c171aa0db1bc99535a5cc16d230721ae538c1adf26;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h36376b081ac675a7e70932f5d2cc85e28caa457d25701c2a1735805998154790df76d607f57bdd792e72891ea1fd713d8adc788005deac76c0fc113a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf49507a601da13a3c8080616d3abb78459a0d75168fafda63fd444b59a19f84cea87ce82e7050fe31481325eb31844fba5354a89e6e245d156a1ffc19;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4ffcb0db1d4cbd672d3dd3b2ed88c2b73d1ca9192662803aa00cc191c0f8aaa79b788a1c97ba80d8496c4db4bcefd24b6737574aa7a75c61e824b90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2c7730a0baef191e3f0c5f5c113c48f5b0130050a39837ab55be6c3e7b5612d2146de4296774efdf164e49e2e7cdb45d15e191025431b820f3045c18;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he15762d88fc51ca05b37b8f96e85c286ccdf7beeab71f48be1665cceb42b4432f50fb221258c86470baa53b5c2372f7866200d631507740c3572babba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h934a005a2e4bdec03127f70c7194cb5a2e4184c88bfec27fba32c6ccbcf02087a4049d24357ed01fb70428ed4d19bd3314a98e2761990035d31fb0ca8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec253ea3cf0f7866780af5f943cf10ae94cc62b7ed1f19db4fd9c1704d0f5209358c8f83b96b8d8b67f9d608416a39abbffa72e52bb65e62f1535e9fc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ccc291fd9d338e5607e6bd04894133d21eb9dad225444ce0579af6f9de5c9544dcc9aafc712cee232410d999a5196f36fb09a49eef57ee7b7b79349c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12e803746442fb498ebafd74a8e92c85b89a2d61a9ec33edab1f10c1f19488d4814ca3ee8d5a2fd362773e3a5b8fea5f107531d0071cbb31807e127b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he5e4485ec4db7a2796b20b1a7ad7a849b9647e855434b77046c9e6b3e982eed3c4cf9486f88912aeddd1475e3cc39763f52333938de1aeb59c1c50dc9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h30458914cb275bb1dbeeb31a197dcc20fcd1a02a95d894b9b1f09d5eb52789b58e6e8ffe49f4faff0eb8ab3bedc6cad3687c7e5a2d7bdad2802e1e8b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb895c80eb486a83dad29c6e8e0232bf5dc0dbc62a810fb538d84110dc3f489da21c88284331bc709be5bc8cd132bced6d41d81c6289415d9035e45ee8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4ebaf4bee9111461ed79955d7f9d8b1dcd5367e92f26c3599ce0537cda8d46f7b43e04349682d0ceb65477d62806b90a6de870c7cdef3c07f899bfcc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha890aa598efe141909ea464a609f8eff03e046212504fd0bd20f7f46d5323a075e20be5cd8fc440d86862cb98b54e700b96ebabedf7b76e24d9199ab4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d5aa774c3abcfeacc7b4de860b11de0450c9373154c8f5ec8974f23476fc41c0e7d676fd19315f4ec9173bb9fac643eb7a0f403d13bfb1e15b925dab;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f33835bcf42857ad11234c03b3666b4f090bf1b1186e26cc957c1fa5a3aaaa76c60e8ad4bcba0b55196e3cde5bad485fda598113712b314b1e43c07;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6d9a625555fad76b6189a2c1910c56feff9ef8f64ddf6999dba8682d06a277152d765111015d454e71dc6a8d016f3179697dd04bca7618bfe7fe44ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h362fd277ccfb3a9a87b116a462df7c8280f2e657a73abaceaf95ee7a4edc07912f347b079b82d97cc51380ba75841ad93ccdf49d4673d3eb1b47f9eaa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7358d03996e6cf6461bec451e15a92533f82f9bc483ac1ff260aec744bc6f2f0e7c0c79285fecb9fcc69197246a13e493295dc348eaf7222ba49cc03a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a5203f5000db41c79068634303fec796f6b9c59b207f7fcdfceda36a04ba0c5608cce13c9b9ffe64641c33b5bd2f5564018f166b982b67ccdb22fff7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h13d1141021be3582661bc7ecf71d9c7bf8fffa96b0b17ef5c66222255752b4d1b87dec5dd1972246e87ecadae23f91e175876f35e637016c6c18af839;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62f3b7c796e5e4e79a4a13f54d8deffc5352cf87f478ab35f8dc31e68221b3eb7173ccc29c69beb98be3c0d97669bc8db7a56cf795490f427088f9f47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h845cdb29861721cdde3a59e9a8145bd20dcf7060e1c5b39c4a573cb3a3ba689cdf2de55bb752c056c8e5b4056c56e78903c37fd886cd6a8ce099908a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b0573d11f6d55f98633a3963ac3ecbd37953f96f485fc62bb40e32b8367fac4dd37a3128490d5e6698d39a0d1bbbc4f84b4192752a5520b7397eccf5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ea28a8dee090f169b9421381da873916a2b0021602dc9ea6a4ec933c128ad18495a80c4cad38455cad811ab0d3b7091b04190577552309c8a0335917;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7815fd20d98c2223a822af65a840781a57ec4c4c1544c6730216a216b66f9004d3f3f0d07ef4bb4d4d8c1cec230194584c64b63c1fbfce8c0c0639201;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf958f9c4e94f76d20c27287521843280a56836872768dcd2c96db79d43c663598d13fff0ae18891f81ebf4a955fe0dcea1d15a3606a05c7a7d52ce576;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb329f5ea5d491cad7e33aa51dc07b8483a86bcfe20a23b1e207e5b54af80469bb002973844a6c9b9678120b3c4651b11d8fdbc9bd2679c28ea6c126b9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha106924ce54bbc01a0715c7eee42c7f9331bad587eb01b29f9978bdb64b8612e464b20b10cbbd835cd846fa890a77b7c1d949d96f274a09d7b5c3df2a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f830b31d6a6f0863cba7f412b44f15479f17620844d75d3cd7adadc64fcd5027de93961ab0bb276fb95d7a410dc6742c5ab5acac0d2d096456a9ae6e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h55a9560990167a3077cfe2aeed3d0f0772b60d00284cc4922f55534328fba0623eb47e40d4487b6b6f0e1192087ce940f90381f752446409eedac60a2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h932c72d54a6736d47405548f1724fdaf1c9507e3ed4c5f851de0005e3679906ae404a8ee6618bda3ee7f58a2c6ea68b8d4fc1934cdbc3a7aee98de987;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff90f1a18e92c8107af82be933d859987bcf8a795dc71e00ac6783a9f064113dd343c26bbd79fdfee0ce1cc923eeb1d1fe266e0642c1522de23d52b54;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5efa7a23bd021614e3aeeffce4e68506a6d9f24bb0dc89bf17a54138880430db46058f1dcba5ffdd12168b6e06d2ab6da23297a1026f6947d39ebb92;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h656ebc9b34fdb98b61191654742c8412db02df9c794b56cb479d1143cfe8f63d751d296b302b6f674d67d8d1d8bc920b3b6c99a835ba597fac5f83ddb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39aff97fd750e3567762c9c2c9172d1105c95b608cc604dc0eed2c8821fcac8a4fc803148a91fff54cf20b1d2956a83969adae0bd8de0bafbc8730592;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5003d24250797b3166460c0fc5ba405030138ae251914f218d0f545a7dec64ab29dcf009959bb89567cc79a7dbd057d81cd1d78c12ecdf71b04a0ef28;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94d657d2d9242df80836e470ff9c70c176d811441ae67051d5979ac407696e0c6d3369c42f7ad45e3ca0c8cf746b08ab85a8f605c76823c0c2d2884af;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb4b85fff62533eb3eb5e3978d0c462050b3bfcbea364bc64e039548a8474e8ec53402aac6b350f1023cfca0c73ff0118b15bbea619b224d9334dda6a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd0aefd0c8bc1259e49d15e2a03716277a8dce08d9e15eb4b2a8298a741d8b7b8d9813323c4b5940549859fa213036b0485f8098ec7a5a7ed84889eac1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ea206f222a382abffc4e227f4fc96720b0186caf7bf52b24cb576c055db55f6de2424391e2a7d2997cd047e06a5ee40203e46eb5314cc214c7328f09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5df3359cb1ae8813b7e526d55d9944804c807476ad7a25f2d7ce9acaeb8c19c2178a8be6134cec798beaa63a5e2137611e4efa77fac8df77a871c4aff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb2fbc3592670ddb7058bbdf19614300ad3466730067dca51a255eb1d4a6dc1e6ca2a40650e05f071ac93acd9915b4bd75ce0055bcc7c44037326aa85f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h546271e2e9e300caa2293fcf0e69acb73b95561ecadde7553f8262b644df05ca53d2ea70cdcf34af53a40e187728720e230c8379f7b1ad505a9ae7ba5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb7240f53cef7393b00cae86764c1fc3b043ce2765a7b6f096877a150ab407bbab1aed0e9304f0fe5f57c4d18caede0d6f2ccdc990545c1824d44448d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9de5ed45dd33755f46fc4b969fa1e93f5bbae94065743ef663bc03dec23ca55983c077bff72d2f17975cacab4789577c83e38e4682659d473ec37d2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h219d5f2c176d9d9796db5f5b1023548456ef85dfd38ae127c6e23f3855a53429502e178592e12bb9425912b7c0b7afebddcdc473efb2d963123192d2d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h86a1911d4b5023e0e46604ab1d9271c16fa8e6e57494737d16a3f59dc8ded52ddea2456f5e438d22f3e1ce9ca8938cf1d03049e10dd59d86edbc8560a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf107aba5fe885b3ce04bc5b256c8e3ab909511e5c7fdda6933ca53e69af64d0951a2788c4ec2055dd4e0ea8690183cb18b43d2f72257af577643a483c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hede17e03617140767c39c01577d4c4f61ac812af48310b3ac39d942b5b8b8f3dcc2529d32afdde4ee1a9de71447e4a230c021d8264b2e0555fcf19e37;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28b9a5a4c6a566777d051c033394737d3bb5ea58d1427a46e66f3fb0e9971f373cdac00345f2c4fe44d514d06004db5e9424652e85bacfe63732b56d7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h61f7ae7e1f06b056932d6a562f3e512e64f9def4f229a50f27ebd70314c2cd17d3be1e9fdb4499ca3bc2540cbbee0cb09888871b7a7490f8d1d0a3cf0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h98519449030d043327212f1900d58c20e8a10f9182a4cc9c48e78997f0e2090ba6073d9749fa97bc6056537c5a9c078e6739a7ce6ac538c1c7f164f6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4f589ddb883d641cc493ef29c7029411e7e5ba96f97623220bb0f0f569458aabd028126c8710c5f0d9df62bdc87ef2c6e1f93269ba3b6ebe5f041da5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had00f6ed9dca1cfacc672197dddc32bc60b60628d3be311a535d6a22d524f8a75e5d08db2260de143ea4b14dd66918f36dce8c7f15044cbcb493ab41f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h97606622a5c264afc71df0583664afa1996620f05a8abc8da9a6f71ac36f2c5423395f593c5cc5132e664aad7968a7337f35675fb8968f83a411aec53;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h817a755e41be7e5ac57265186252a5240cc748833293a63b4337da0b3869b5c62a2d064c790c62dbcef1d723712a22ed6486209619035bf2a2b05ee83;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5ad462ee9ec340eea178cc05b2d89005fa35f5b6c1cd733419ec8ece00f209159574351d53cf507ee8f405e6e2dbc749837a5b55a7341a7d206c056c7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha9faeb60875715709765f2a62455a2a5df1ade2197cf77bac5ac90ebc2bde960ad50c662f358ce1dbbdf22fcde9ba802a14c0c1aae4438ff9c46c9b57;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4b6af7b4dcecefca003667d164b8c1cf62198674982c019c79fdc40a997b478e9d348efdc979675a207ba4c35fab1744b1ba00119affdb3b893fa7a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8126dc34c73000d0f042865d4135f26def6444c82494a4ef8bd1ced4f1d47854e3f7b312c2c51a218a948940f4f761f2f9b3c89a55afa054ee1ef39c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h111d9b53df6d146a4776e606b38015ed77922fb6203a9ed7b8252336a80c2725cdfb2859016f32792b1c1d5f5af6c2437114be402d02e154b42197ebe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h619d70c0e5a57c176a3fc47b292ce6ffd1656f26d6e62ec46769694eb6095924b2026754ca9d5603f226e6b96934363121481b9d833e674ceaddde04c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb8cc3e387130049bd101ba1881a0f348587a74c5c8f6ca16c0f2d795cd17c8d5218bda8052347fa24ddfb370a7c9790824d9980e29f695cafdc416d19;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h20caffcde49b0f6cb3d48d2371b649a3d3ea013d04e777f8cdbbc25d988d211abe9eb34c4d79105dea433be5f1f189c922d1127bed74e43f8b7b54d12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd72bfae56e8a47bda14bc0f24c54814de863a769bc18d22a8e1e4bd8d664234b1d3c2633cd08f3640abc285077540caffe6e49adc439acb7c655cf6dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h462a74cf2c93da3d8545d3837064957b9864f31c9b5decb30fe9b6fa1105fc3e54d19bac88f29d2616920f5c35e101fd8c93e71c000abdd231d945b29;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9b90f6b612346ea87135e631d833a567fdf7bf1e35a5809dfca9e10409a0f2efa436a7195193dc435a50f4c9879c9e461f5414017f284ca8a0c5c2667;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84ba6247fd21d06283d2c4f02b9e644e166651103e336400c360fa0e732e6922d7eeb5a3e0e44117ada8d2eaddaa72a7da4d0cb1b0bcbd83888a82b07;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5aa1e15ce8cbd596cf94748646f4b1f2a1d158f7cbb16eac3b5535e0b3ce6ee561bb46ecb8622376569446b8b8ebccd0c0ea9d7b4906181a749c394ff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haa3bab3ac22c656c5d96ede22e6a5cb95f62baee739e7ba347e71c99d18ba5670d68890edf7b284e273417507307dedf94dbd166f950df0a44de8a4e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he636007544d2f6d10f6f12b51792b4aafde9d1f629819539bcdd019a2c816a4d6ffa99cf5f3f8d1d7a52c8a5ef967ad66fe6b83ece31cd170e6ce6600;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadf159f6fb71549a4246bb0a060511e406c65f72cc2f441fc717bc615c9f591fd44e8679f606b112f9762d393ff90d7faccce57047eef58b0ac35f17f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4420bc373bca08a9385aaa2b77280d6a25c06bf67ac3e4ddf8a583cfa2b849469bcbae11ec9bbf9faa6659657e0441462e86086dc7487101eea499d25;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b1c37015dc55983b6be096e8ac282345f2135523f817414e366eb1e41cadb17ae3911bd9bc8a79ec14b260ef2a41265cb9d7e9c8f60330eb451e168f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35a609d97d8ddad56718872af87c1e75665f555d0d2caee728393dd89af2a07c047bbdaee0119c426fcca77b83d200e94a2485c94bc9a968928823a29;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h938832704aaf087522ef67c3cbeb0eb9ea9f739d49941dd0da7976eb6b3214eb56c2dd45c5188c7f510f2efc2391efb20119d83f5575ece47bf4e9316;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb16361ec3c3c0de252023bd3419d4ab7c3260de29918135d4d7bdbd4803cece50e76bf49729c38d26ddf2551de33ea4e34ae4e4c31233a25d685850ee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h12db70b539b79915ffc5123662eb32bcbdfa21f8b0749181905eea5168a7bc30693a083c548c402e25483575255391548afcf858f5dd8da331287b579;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcef8328fba100e477ee70c187a93f5808d51d69b6f411563019a173d9b9b0deedeec2baa2760b6a9b17fc07875bc58dd177de2d143e0ac79304f25777;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf37054eba7e2f9fb650816fe01224635f21690524bf19a8e34614c4f5ae1bdd4a9010eac2a1e2d4b92d48d695732b8b7cc62741b106e12c49b84cc194;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd51cea453cd914b91e01bee4dcd62cd425969a6e31964fedb773cd912b71666f8624875872130ce8b99cc944c53fc850a88228d0b3a5108baca20ac2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hff2d9f24e80a229c2fa66b631e36f2591cf45ad454f15c69e528c299d87b2850547e50acecae3630565098b5ce3d2bf82bb9a843fddb7ffd7836b5032;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4de1cfd092b694dca6a7b17b0d4a6745515c66a2cb870568d41d167a3e74fb5a6bd60ce159ac00fd2e71f94d8c73414c9d12b18d9eaa40144c20524e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d220d6358808bd35f101d4657312e9403e90fe27037002b7961d91ef0af7392d242528eb557dcc3c29c1472a8b67d787d8d64549b9d3807c788cd775;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45ade9a5ae88d9ebb8138df2d7298e152486f2e24427467cbc9ee7c80634cb853c6ac3ea5bcbd91d8045ded878674b4105d890660f2dd0506e9935ed3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8255cfc00b4c674e83f36b5dfd2674db2cb3567325777dee25703d1ce335055483dbe707d01f03f804ef82a59eec3051793b286497faae37e7aea98db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1200fac0159cb044620ff11fcf49ab230d4405b4720f41f300e6c8a68d7e3c1bea650d3538df9a102caaae65ec631e00e1c251883bdfaafbb56000882;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93e4f5a92a6590c8d3a4c50255a426cd1319e1bbc84176a59a9da84457a01793c9e1dff5817acce3436f60e9ac657a0fe4e265efffbce224a9d9fd0ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha24675b8a9bfc4100038b42756281d211edcbe3fc21b417bb868bb6d64122ed109c8d8eeb3d7f8677ab0b8f5200098e123dc9c44b90fc970f18f571f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h127eade96935c345a4a9b1770d9751e6273159640930b8e0926220d57ba35ff006857e17858bdcec4a24a765e9598b4ce38ad35c1040643b2c15d6606;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bc871ca7245d7939cc3a769c4477e09bced6f1d487e18d02f2ed623242a9562aa67cf61e544a2206da4205b294ac11127b8783cad76a031c33114303;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc5b332f9f405c5dacca8338ee541cb3d85afb0094b596e369bbf44062b5672dd12a8a5763b7ef43c27f8899ed4335b0d285c9ac2a38dfb8613a67a86e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b661ef728ad44a6c46728e87a5d19ee3650ecc63ef12c403d6c829b9a7210ed7f3c33fb86248a60166cd1df05e4fa5aebc0de34b22cfb4653497a1ea;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h830d55b2f20a0fbf452e0df78ebc0de38c5f1ed28416a15553efd0180182e6442915be936ebd3a93c9f0ba441f84a37a81d6c220a06be1a322ad79332;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf8b9cc4541b00eef7bf27db2e73cdbce5b8f9759e5d8664755cda10735d6b1a44f99eed960157c1b29df19ed104d3526632391c4692718e1ce72d810c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h106e36bd5fe61c4f3840292dedbcbb73050eae1ea257bc2a9b28d05d3f444188bb6adce6b05a1488f707e7373da461c2ee923ce9c02983723694df75d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc6b0a7be8353652c88291f33f4ad9129c4b4c095fb915f8f432f5c65bd25670ea84d6ebd0a63b8683b040657fe5d58153dd7feb3fdbcd11382ec78841;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a95213d59a5a9287917a41c16033c76a3e5b75e0f8854aac226f96eb534d004d10ef727d91b7c77edd8bdf15fd6b0b8002fe02149cb9e168987c3767;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e032af0839dab98f68aa4ccaee2788a1a2b037d082e05034e18ecc913087213587f4ae0159102ee9943535c84d221b5685d811482f71a1d8b1320b2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1555db0296b81c63f22ab9a49bffd4d6daab8256213ddb641106a1246da1c653477e7cc73395f9287399e455da2a6d97bea4f12c642f81a660a4bd7d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8e27aa9df9b97946492e4c5a967e391a345fc9d5874708100613ded7740a6b87d8358c97e87b7cb473e1047b2ee38a5aa4a70740a61a2c93385e02ae3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3c805d13f96238c1917c5ece4703a6e693db2046b28b83283770057b00771b2b84c0fec0c9bbd97fecd23cd52b8e9756e623440f0ef7238bfa526fb1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1ff5b4d1c9787efb484dcb5dab987bd085249c130888f269d55685dd5827425077cbf34393accc57bd0096ce458ee66df5711d2e7030986e6bd82c248;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2335472df41653f3115153685067c4d6f65e86bd5fd6fc01f64b43333b8d5eb1016890d06e81bb166964708712ba6683e7ca52bae6d51ca36e75b2795;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb771d23d85a5610fdddfe61a981cc6351bad2f4a1a5ff67380f5fd931d4a51f6a2e3913d59d0b18d126f28ec222c2ebe5fbd6e72edb63e605317584dc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cf6ed3f56a895b41bff31560caeb8c70b24a9222d64bb285a4b81bdafb6ef5344a3a1c74057672b5a194d666b4d7d96f47e4faddaeb674a8a8924d45;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had02d9110b7b96adbf08de3c9f03bb265b71a3d8862dd72e43d6a43d996ba6789f538020ebfe7eb7cf34e9f63b511588225987b76d5caab3cf587983c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heef9b1017cbc9a81d70274a9ba80af28705a6a79885ba2f0637ee993dad33d198fb47e05378e34b4c957b8d31ae1976823e01d96b8571e01562cc18a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4bf99aa3a218235d5556c2739e92a3c3be1135ae0b272a06fd78895996a2c1ceb89e2f157cb5ccea96a7b228ba453a877fe4d010352ac419abc5c33a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he98d3a9a44a15d06fc381461c5f63e018503e04f7f27d2260076f63ef55b40f98c8389d20abf61c925a2a56252fe60c87187a951f5e22013208d021fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0ba98499b84c0a0bfea5bbc83503b4e425d266d860ecf545190d90b8529b7bb0d06a1eba347af93f59c262f3c38e2bee8d69a24b32359ae8d736c6e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f4614e395dafc7efdfa48887396ebf0b5cf570320d865593fe4369794f05d5be1cf844819e87f5176115a4387c3b7de9a9cc412947362955d33e181a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc28f0377e1780c831626570ce9063c6ed278eb6ca069776e5ce0e3b7cfa4a4d9de7daeb5c00fffe34a0c3a6dcc04c1cb89bbc10c01c31dc66dda11c99;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habb57d1a6283f374b403d1e82810cffc08f48f8b69df3414c46deea869f022b7428f229f342bc4d3ffbf52b705af937bb1fe30e13575f53ac45cd7a73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c1659b714de95de256ea71cf20f3dd14d37888a5bf6da7850904e47a13fe9e1f3012f1443c61721aef9fb4bb60eeafa183e9e9cd2ee73c0e86ac7d7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb9a039b656973f19f9bff9376d82b9fd715c44c6e7ff6dfb78924b0c689c251e4feec0a8396d23ea405bbf48719dbeaf25e2af66b453c3a1ac77bd01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc184994fc02227f9f19459e58ef29157c9a6b4c5ebd91abf66f71e53c5db97456081715561d77f174a251a40858bec1ce2df187e75788882f144b36aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf61d186d1221c6bfc0e6a673bb5bab36278ca2057e0efc16c1a1e134329fe53b23f29ac2997036e80f138d8ea7da1c566620e8db4873d77b89fe54739;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7773a951a9ed9149af77daee956da210b61e614154e9099bf02014fa7d45392af2c55bfd7fe58c16d7f95c980aa14105afc9ad89a4f41d645577485b7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd83c0e30b194305e4345ce596e75d4541441373f4048ce7c2e97e6eb08aa9721f3749609ce2cdc78779300e01e7cc572ecbfca6306e975d00f6dfcdad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5eedab2833a749dee59d77bcea7de80feafc33790d97d2612d857939eac86bbf8c7bb20de2a18d690166859500f7482cabffcf340ca8525a973a199eb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h18ab30f65e5056bc04c97a57ff02e4145d1e65c70739ebd796e993ca0073a31c47dbf5827f3ec30524fac953da6a2d75bce492b1660438e9a66207836;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88b4970c31d767dd27caeeee7c709ef942b0923ee5cf9d66b54bc4b7db325bcf845b7f54595510b4a14fb11295e0d5cb9efc2e8f428e23d3304200bd7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h375a74c8daf0b5b121dbd416981ab5c618741a5c01a9bdc446d443605971bfadefd285c252067e6d710dbba921ba154896064778d62e46c59edf0c9a9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c1c8321b77fed3b56e86c7e9850a875d61b10fb21d4a13644f9391c9f0509d4fb96622b84a089f13c12762aad988850e10b832dbc32f9e063d0dbd93;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hadf0d6e739bef710fae839004683453addf0feac3b2eae840c8cd1ef953ac8ef827b265ae521f42eb0a4dad934483fbc519b3cddbd9aeba197fb077e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha8b6d9b3f913792ee47a4558ff71b6c0a0b7a193d4e0c3a429cfb9a6f186ed1c4801cbf3961d0472584bdeafac77f6ac38d881ea625ecaff32ca74035;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h29c7a173172af68848de1496395e234a7405fad242ec1f2ad68525762b5aa98d5fc38eb916fc21e85718c5c680ef962d84a0c9672ec2edeecdae39949;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c6965730408e0eab224ba5b072eb688b9e0b9c68338baa9f43bd8ef93d11e0c1acc810b278a9cdf06569ad27cec47b98f9d4ae015257b460380e6fe4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd30732fdc5dbe4c2a8c3859c4c97dac6d0ce4b518b74c88fc982d1efbe421ea8aeb4d3dcef22676a485ff861eef515c5d49822f7f324fae380b459c60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h939ccb6d28f4bcf81fd6e29632122a89b656b9086450db91c7630246ff7464a0208576551be21a092e640545b593a1dd5fa9621c4f67d63e51dcad1ad;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8d601e53bdcf02a93033da13a05bd3bda8d5029d5b92286b56bd38b360536ccc0372e8cec729e23e6cd09e5eb6bc8a55c0831231f047e6d22f4a64a54;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31451c3ae4539018281773e7e03de294d5455ae9ec650221cb45080852cb0ddc517943e10f1cfb16ea0cf525eacc4c8f95249d9e989df90f4af21e995;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h613c97e649e40b8dd16d34f5946d4c7869d9ddb2054e4bbab5c999d676434e58a19320d62805d9397abaaf1ff26a5f1957937075ce1269c7ed2308353;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7ed81e485493509b8e713735eaf5e2e4254f72e533ddbbc6dc216caa4824cc51dcdca5d4e9323134f7ef0227ed618122dfbbce0d8d7c3666095fc2a73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h816d00d65b70f72cfc9a0858e996dd852bea4d1d07160372d489eba722f7839210280140371ad2e26abf06b4783f0eea5dd5faef5f0342711fcb4b154;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfddb31ffedd87d5cd474438f148f53edfe2ba25119c5becf9e482c4a7d34c473d33404e91ee27d062a245436e48efe24d485d0549168aa24a46841513;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h342a23976e854bce505542473eb6f303de6074756b5fa1e81337e85c0f45ae1d933b4612582ab212c4fa70756f346023f2222808d8b127e83438935ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb32e379e9cfed160acb880919ea78445d77dad33a97d9b46e44dba634090d544a3c0c84a06317ebc01279c9bd44b7c96d7019c7c081a09980e42f6c04;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h891f3b266e08d6439a51d606af19f9ceeb78113144f2998fbba86df38365b70baf1fa95c5a3b6982c6d578f2b5308a91ceb0fe18f12d3b8a1be9c64da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2510eaa5ef74e128c94839106a8acb057fbadd29d681f9f5c3be6af9868b6c8805ceb46b01e8c69e6012b6b24941f82288edd1be57e77ea8dbea0f7db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a735e63d4484b9e1a0af017dd91f23487ddefbc0e3d0b5687b7471259e8a9b8bb28a5e3fffb4d7073b26408cae34e004efde83e9867a73e97d7124a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a0874ebcfd1200919665cfa39f997f449e5b5cdd22d975cbd5a4d71f3e5571fdd5bc6c018ef660b4e8ac7a15e89516321e307760e743c4c5ba1ab3bb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2021b73d6710c22e2453aecc1a64c35143d40717f232267a2f71c5177b27b1e892850ad84a1cb423887aa88c083b8391779a0a1408cdac591a70591a6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6427ef9c6817cfbaa4f87aa6566c9c441ec89df6eb25b2eeeeb6a3e005e42054a1189639f8bd60f585c5a57601331e6b7c48e8bdf25276e7a2fe127b0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7656002a6e321d28bafbd5a74ff55d7aebde5d1f8eb8b6053dd28700d50093985f8994a8ef2af24f03b1370cdb72b9daa88a5ed0b4e4fce35fe6b6659;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h62fbb56c43676e7a05b652762849e3b5246cbb4d99cf274e3af37b4d36ad7dbfbbcdaa5de4fea847e47bfc513711f6adf24709e475697c5d8ecad5e73;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h65672d09cb7e362f828fb7f5f8157edce29d95edf91f22ea403734dddd6595a12545e3ce65b63f152c06613a49390d44431939c425b8c8f449282cc05;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5d2caa34aa1d536933d037a3ca82f428ae8458fd38ac8c5cc52a3e0559aa5f5e4ceb0550b0827f362723f6958150897819f4d768f0e60b55bc44cdefe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h88a50a5d59b3b1fbec869e09a007d8d62de958a4f19962eeb988e4d2044f570b27211c60491a12536d48b0fcf6a30020eba0e483259a37e13b4b30363;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4e78e9f070d953970134b384bd10852bd90f267f4997795cfa213a5b10ce0632874b3a63608604edb13e4ee1fd95221bcd3cd52db1ee4b82e76c9c82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc21d47c0d0fb08084a78fb70ba0fcc680dbf46fb9c5b35c0e3747fa803a6c585d23f6545259f6f91d0963d6eb86ec47b786033a590855a485e7e24b1e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hccce5190cab018051d35779c4098c9771d2545dbb18241606155efce34bf6fd8cc3e33af8d788cd2b8daea889bd3110aa16fdc58693a7ba40f31c548f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h84db2d2c79a88b10fd0509b97ca8ba818a8e2af066f7d9b2e049ab3a2db0c6f201b054d16dfd3a0c6d3ec6485fd358d1b9f46bdea2c61d2905dbfcc59;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ce6ff575cd8f474ea95eb5ce45df500dee24a2189ad1f57ef30ed756a876a27b9229b2e7186f3e2368e84e9224450aaaa119ebac744e98cb48cef8f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf1f700da40411505bc4db915f20387149fecba9accd3250ebbaa643b56d06d6f708976229dbb49bab97b5fcce61d0148d12450ecdc2a9d4aac4c4b026;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4dc1d573d6bf3920a64e1566c32bbe45b3a2a04ad15c4fb36871a3745e6b8be1e1dc01e27a1825951eacfd3e0c6f8ecf49cd4e3eabdd16b700b10c8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79a95d6a9311b51f8061b81106bf3a21930c849ea9de6f32b3a35b4c19048b3dc3f4bb8665df9684298d8f80f4516bcd60daa7bb7bdaa38099886844d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72656f45fcaa0c494f49b5c5e31baaa875e3f812706ac6f29770e308d815df9ce2c39a3686f2819485422f5caf74006b3487469eda3c990472f94898c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'haf20c0843dc593063bd5abbf4de4fd91744c8f53aed7034e7e3d8a3526100d324789317f95f6e5be01fc3d7503c6523f0c7ea412a2bf6e1eebecc077;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfdd75c2b64f54cdf5afbe9bddf0329222e281916020ee155d3499849d6edb5b3ac4e9eafd9f526307053a5ad89d96936baa1e7010d82d33ccd73e059d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcf341afa4c4c11196371dfca6f142e8834dfb4e36bd499f1864dc0d02eb8db69ae978a609636ec355803ad97fc99f9d9106dc47332e332fbfd582265d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7ab4de0d2e9caba6e697595b98dbe13baf7505f172c8ee0c6842bfaa9a314446f0fb9712dc4c41ee29862a6cdaffeb498df294d5055bf09dbfadeaed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71f662a518cf386e7f9e0a69327372a8f830d3a745849ddb52fb26c82c3b4007874c0d548f9e094b93219954f90baa3a513ef7932c4d1883fc3bafae8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd49f7cf574ca9db9f10f6c0f0aa8496476cc19988595978a0822b99921fc286e3b844d8e3dba8fef64ce14bd26982139bc2e45dbe03e2b65953af1330;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2ea942bfab41ddfcfe14d510d26487224d8eb7804452da9e9ea0c4bf8dd61769a83154f38f772245bef7929a659051d3cd02ea07e941854cf3b59a2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h570cdfbe9550be3b56389df894caf8f35faeb56fb2b83af634cb30a336688b201dc3944806e757d084d476a86050536535837d6411da03aab9d7a1efe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h78b551b5e8656e1776332995100983486e2d0c6255a8d350b13742250d7600021f476e7786878a8ec1c3cb856f97952e4ed6f2b52bead28e02bca9ba5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ecf736d0d151a97dc0931c24db4f3799ba3784578b69183891fdb9e565dc484d37a7267cbcbd84dc77b7b91bb9f0fa4560bf0892614574f3c33a2ef0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h853a2323d6bd4cc301d997fa5800d53cdae64c2bf823f95fa425fa59ce57db67b4c4f6d8ba4d4505527317e4c2cd26cad872e7fb8f77e8ef01cf9df12;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hecb1e1c1ae1aab681a0ea2fba07e6a2ba39324b5f10252ed0d93ea73beba38db7467bd2687b4c59a5cc06fc758f773dc1ede7e80cc3c9e34069f8d401;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8806b4f538174950e7a6f7202de4debedc60116a0a4f0ce1ed3d6cd21a41a918c406b488c3e6693c176b5391599128a7a137c103b24489f8aaf78d8b5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79cb80f6953ef8b07dc37e7f0de07fdded7ad5ec732b5d92bcacbce6b7792a95829e960af6daa6a8685685dd00c54a93221229b2ff84f3a4a5a27e21;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ba1823229c6cf7fb6862273cea0b68ad387d7bf2336bb19f52261af7b71944c4d751719d8a084b469be362590eb005fdde4114994e315c88b98d00c5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d20bdda6460c2321e604f0b0aed05bdbf62fecc32fcb19dcbbc58d41d2520056edd91d85ce856b0aa34bc389588e3cd34efb6cf230ce10d76f3a173f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2ac9a3d02de308a530580c2cc2975013e6c81625f7a267bb0c717484e26ac124bb7d46e19d1d05c35da675bef4c0d31919376024d1fda4af237c53744;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf28213318f3a611987f2629c53c0d99ba0888991f4f0109b44bd1660b54694e9f3ee173fdfb91c09570c2e6a2686898622cdcc08dfddb3c4ceaad43a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h53d27e537af3d2a0be35efe54897ce67f3dc2dfc42664276d37b42ac5b83ac3a8207d4dbc0b3f54619b433b35bfdf52fa88de970911d98cfccaefd493;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75aa0a13a990bb2393e1422465f430e096fa4b2f39712b3ed7e5f88cade14bc0647014692f077d575f43d88deba7955c26064423392f0fe3273995c8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b0f2a1d9fca61a94a0e07d8e9ea5ed989a355840b36ec0a32144ad62bae7038e8ec9e784c08f38d0a1d6dbb63f840b1e1d2ae2dd9846557a09e02595;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h792c020b48d9c70f975c5921846948e57a5bca6866c63fc5d8ec38b1d1c195ef1b9f705956ad0d95fdf206b65ae3ed27dd7bb64d000cbaef5ca7e9700;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h849869f9ca0e8b29fe60ef4eb50289c25526802c9df96e852d8675b4e532c32b9552eb04bda82605d55a1fbdcbbf742f8218cf56611d78a5d6ff05546;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h849f65bd8e39da7470f7135144859d9079471434b97ffdbe5ee2b6e5f1886a4011068fbe5a39cf4a99399e7225279150650c7e9c6b527882aa1c2290b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9add22e222097a4e33343ac1484a63f6937aad6e4a355898f5d1ab9f70d31260f543e42b75e66a7f33ce1d5ea67c5237508c564c0417d430d97fc69f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h511e38a038d314d490a75c8f2f1f21f34c1194aed9012e16c80f264af6252577764b1c06152a95f9641b46b19fafc3108bc880ee8eba10c6071911156;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fb0c96fab687344c5ee155cac9deab9be584d207a42a809fc5bb10cb8ddeb17e0b632c2bb929dfcb56edf7f30643d5dda8cd6123104013acb84afcf5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h248cfb598632727f75b7f4374777ded5524058fd680a61abb31d4196ac6ade5320574ffdec87e792ae6a593ccbc530801d6f4f490e5e52c42c8cac8e5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1170db3d1f0e66a8f52d149be196b1eae7654913ddae0f134e2720bb5d1ea9e2fb963a10be7883353fbd33c8fcf8931c927f9384ef752488d1c19552a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a39ae3c4a7cad2d431a505cda93282c30c74932f90720c9302a5ec5c85b3fcb655ae0548f2bab5f092d2c4aff80cf8b9ab2c19e39dabb8bce736ac8e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd4415dd75e528d65d0caa1712a99415766a8b3ef9f5a540a33a05f21fdbb9f80c22da05fed346a35f998ea4a9d8fd487c3f59a48db5b38a6d0110f6e8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb6949334472ab61b1bc81b229336704078c2861ba274ab3369f3ac816adc5bc665ad00879c7a310e0c209d7971771086d84bb09d5155a7fe48c49203b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h93710e349d0f40bc07ff28db6deef39a81bf80c4c2c21ce2a395dca28283f5dc8b7e72ea10ce5d5f9c238dec3c35cb6290017e85e5a9042ab05397a66;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c3639e9e8456c5b3870651a7e14b3cf8e6a0f428d412b08dd64bf72f3955389b5d26fe67ebab69638f56aa1d896c96cc46d5e7a8a42be70c06bea1fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd48c70a88a1e92eca841d08393166a299749d1d83b58fa44a049620ba34e80c99fee893526709edadb59553a493883a9e222c7664cc4e9f3c0c2fd2f4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h124a2dda41fb729d0615c242cf925bfc544cbd82b73c035f2f9215f0e224c53ab10372e2c6330b25dc067145426a31ffab3b6181ad6284ae53a24a035;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf2f930aedd1613f7381519adb2b2965fb01e91a9eb8caa12001894468f04500e80a812f804438ffc63ffc0619de3da2b8f73a736ca2c613b5fd615fd5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h25d542ebd71bdabcc833f0135b55acf38ca21afcf2a8f0b60e789c7ff598c0cbeaf65da97383f6da97ed862e0fd3787cc3e146cf781fe7fa529edac8b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc8ba49915e043c7f0854c59accf1788a29de8af3ec13e1693202bfbff08912dc9a64dce61cd8c922fbb84f4d586e8cba0bd1600d58135679b987a4363;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h631d3480b04aa4daaf74ca481b929da0c8d90ec71217dbdb3e9fdf82f6970254e732c4869314efdf8ed1ced9a8ac48039fd399134e47c1c9bcf892aff;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbb4e73ad8b77af7872765107618b5ecd1e6195d61e0a030d6b78c7777c40e41845ea0ba22500faa523cdc1ef21fcd50cda3c356aaf46358f5add0c2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h551cfb1f0d871316fb56482830c47dd68e23da85417942663defda40c8e3abf351c536d6822fbbace30769b6a1e09f02a1bf33fbbd611ad5d94fc860a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd543fbbbdd4b9543b5a1486bda439161e9356a60682385e8736ef7ccc8df02459854a4359394f4b92cb7ec80b3b6bab5da6d12413682edb7d2e6ed82;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcdb8ce78b661fd528a6fe3fab7ace3004ad5924d65fc2f02d92a04882f616e97587d990b3b2ec5aa49669f2e2ac5db9c57f56bd37fea20e3b9811ce9a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3317b3079b4695a9183d9a0e0cdf9c4c3dad24866d370e740196a50adbc284576d62b6c1db567fb71d2af03e8a1c3f1d85dab7f8eaa01282d23490b03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7542e589fff8638a1af42ac526661cbe3971d5830c9aea405e66941e0a3fe4f56653fe2a8f25f5b9902a18d56141ef6e77d49fa3d702bc82e271df203;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he64892cdb0e3e59b9940cb2707975a698b9c4ba860794b139aee38107e3cbfc546c0ca590f67c0f2f3bc2f16c58b786dc6714cb76292a37c1e3419739;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha760cd4923597a79c327dbbff1278d82c574b91c4a409b2fbc08c1a542ca00a9cbad137f73edc2739502d2da4659a9f185d80b14c6b8427740bf2cd86;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdad2b7dddee15ffd770cef8f42d16b7e93b352e3f80157a3ac4396469126200fa07741e562675e6783fc378a82af2881ab25cbfdc7d96d7417f01a0da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h21b8a17f1b51a1454801d9deaf6b34d3300271d7454c75f188e53d6680b86571739803b8164f809fce10fd2b759bc13e827c7aa63f7279de24c4e8625;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h49ae1f61a0b08defe844277089ce9d0cbce4ff142f4d7d3de509523c9faa9637a06c2bd68347b13c052a0a6897863b5afbde76f729c10e0391de54335;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h300b1202eca81f8795400eb5624aa3973cd81591ef367e0a18bcb661c737169f881a00f4aec429893e3969d7fa4fc75cacb9c16bbe292b2d9f41755c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbb2423e583a63616ac1a92af6ff6ec3cc653cd358346c95adcf75a069dab1371697b8cf0810f0b13517b0ba67d8ddec2e3a5a67deab6aea722f1cb244;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96422f24003c1595632a4f3279bb91ec591fc65b34b806bfe3f8464a81c69a0d645ca74d304ebca7303425d5e9e008c88392a7d5aebb826ee4e8cae88;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7550cad9622119377d47cd1c991cba419997b1c41bc75149e09978faaba1e322f3d338efd3aa782b72d25998c74308cf5d0e32850ead6ba627ea975c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3962c1e90d519bd6088a855bd8e76e4fe802e0d1788b6e85458b845efa9a9d1f3cf5b76aa51e8f609794961c13b2caf47176891ad1688ad2527d1378b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1182320ed7a4f39caeb5ce3901e0aa1192d967c518ac4c7629ebca53006eee7ebdc7c4b42c6689753f2feda4abccda62f6ffc4c082297e8b373ee6485;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6149637f43229c0a81980c52f7a274d30e8bb6de2d5ccae3334f121d8fdb4251e117a1afb15989ed1cd98dcc72198be2625f05bf3a5f537bf1ef2622c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf242f805ed50b2cb51b6453eb88af0ef9cf19858f62d00013318954471586712abe75dd6d5c55f01371cc47733c159802151415bed1cba3603b475500;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfad64c1afd2c07fc86ef5fd21efefcfe2eeaccdc0dab7236ef1fe722068e18013e9c1449e4a4b479ae247f038be5793dcd903010e89f410e7d72a6512;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2750a05a3bc07c6ba4b164b4444893d3709c6ed343121b4b61c256625e6630d50c16ad51a56ab54e3d5d3bf94aad99746ff9a2c71747e140aebd6f04c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he6028d60ba33149feb4b4068aac5561e39b11257b901d14844e562bfb33c2f5c452f4a44a1d40fb396b5f0771bbee268302b4198a372c06e00697a0f9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha251b0514ca73128c27f5c28aaa0cce7fa362e7280dc64ebbfe541874a50d1eee063751c12e7f6a674a78bdb05aa1c99dc392112c6247ed2d1ac62cd5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h721b79632f4566336ab8e6f086cf2dff91c9d5629619550f70904e3b53ae757be6f3687c501bc783de011b03117009a315f103df0256f8664684d0103;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3f1e1757d3f4568a9598fb7fd8e94d402ca3432651a732ab0b37b448e200d0c7e6b802f91122dffe676ce1dbec66536fcc0711457124bc87168ddc54c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56f12c511b2e0f86b7b03282bda9f7e40f0f02ba0f86d124b44e8faf25b13ae364e8179d0676935637557bc1a0d5f66ae2ca4e2457fe8a05934004934;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67ee7d7bcaf86b7d24f79bbfcceb4b7c6dc664b78fc0ac9f7ff75157dd61ad634768d6230429208e6bf0543bcc4c681fa6580f02465737882f5f617b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h371adc7188eae0a5258765b3101c8836e58d2efde28526da6ffe3c6964e6d41e48ffd55dca94db704c27c0cd2302f09354a099288a3015c891465c3c2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbdb4b7de9fcdfe57ce9b1659785ca319a8041c18817e5288ee63fcff1e953960e229669279dca494906641b40837ac98bea4a7957109913941a139688;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha3f8af0cb79e7bfcae0a7b0b4989ae086b50898cac4f35fd562789ad1a9e3c2b41c0b1c1cb2722c6c436bb2c06e581400150946e43a1fa176cfa25de7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb74b8b7c3ae6d67da1fa5e470c9ec52fbe8936cc682d9cd135db70c06174f1b5a3001de077f9c1ccfb664bd91b5c1cfccfc5a0c1fb509098c6115428a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcefcb7cd38fe20bf9b010af789379397e785ca19a73805792183111bc64fa51ff90d6607748d9faa9efe4ffa56ebee401cf132c1ad96ef1c6411d822e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9cdc99987c224a0e00fba0ba7329bdb140f53fe8c63805067a02021596eca8048ad530aead17c9a4c3235042619553a2ade8d2521c1cce74bb7bc7bd1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbb2432784d01f1af9226f22e7607b7d987db8f44246e74837e782796fbd9996abc8628947cf11a93848691e6a880c74e4ee3afe4a09a51ec1f1c859;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha7c73a25c200990d7429525088816aa700188b7493599ea234437264a060062f9472f945b58ed7f097a0944c9d9c15d7547a3f69239fa12acf3514f00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf52d59de904362332b2fe1e71f14efdad99a1b0e50b77d023de620526a4432aeab423e23a55075921a744d18167ac67966effd025fff85f34e2eb4936;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd973301ae2f080a721e26794cd7b57a43f18318eaa96971e1eebcef80c7f52e83c641de3b1c030d8e59b7d72616e6372d52914cb676d4b2ab3652fff5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb39c253b010e88d1cc989b5688b349c78fa6c7ad5268c94324019048c838237db27a90fa8182215e2ade7d21be31a2e18cfdcd849da420a93f2cea4ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb42f3996698a46bedb5e718a4f9087330567fd08db93042db2a41e36b61199abedcee443449056e7695edc44902669a17674b37e7d03633ebfa4f9e0e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec38c5bff18d7398c839f34e588b0fc797f5e2dbed6abe483c9651db0abb3acfe9505769844003f70e964fdb4dae0d88b2a8672a78b32942a73c6bcb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h28ac88f7756497c119250a990d96392512c18d41d9835ac42d4eb96d9eddf28d2d09a3207172ee0109dcbb8c475fff57fba7740a0579d2c6fbb31d0d0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h322163490221cb1fc9fc8c56115fccaeae8c5d8388413e4804377f9c9eeeb5b68b69a7c9a43a954cae27e3dda9ec771152b8e2ffc77b63ddbbcbb05d9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1515ddfedae15a0b397f0575e22257d243ba2b17b34f8850d8b104e120069be5f908c33de10a218b94b46d98b6725b0acf2f78d0123ed86fdf8bd91ed;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h516fcf7f95c20eabda6e86e15414a4979d5336be75a4edb11f3a65897dacf9a67df3417348113048b084b1a9feb9b286d110485cbfff148749d74c4cf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15e2bf210c36f23d81791422ee3febdf1268874020a10515adc5c434ea62cbaa243b6c75b59632714431e29fdf1ada72e4557f723159c050ed4127768;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebc620c93b0c418b03c54367750621ca61440b5d2126f3809a69b451212a8adf8e9b8c0eab936581fa6c04f46fcdf4628278135372fb97259016ae70a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87ec47dbeb1ffb5e5798eeab4d2ce33002b3c0102e9733d3c119ba4c70128609fbcf81bab9f45c8a86d84f405aa91f8057deb8577ef1b10d442e0bdfc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'habc8a6bf894eb5d05d81ce099f015c46d4c860791f55128c93014ff7fc4f68da565d98729808dcd215007ce0df0007657064101f748c1ea1b564faea5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4c852570158ae3511e9c94144275446df2fd1801fa162d707d25fec8ef330fc3daf21b8b0cbc128003268439e649319085b90767cd14f074c233cf60;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e17227fbb6963404e555eb40cad5fdda5d5e7ba028180f28592af4a1c0822c14eb6793d91afc20cea1da71484e5237c6ea953d8c03262d21f848f867;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1194ee914b805557763b89e43a2b17434d13544df74ac0aafbbd6d5472177f86d10cadd921b703e49a87043be8b3e957590c4a30e0975d65ce1232765;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3b804896ca8c75e7294044c3b7e3d6fe79478a8c285a928116aa3aa490bf5fb36cae2affd0ddb55229bd6597cfbed335e03297ac93960c82200a94a96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc4bdc9f7e74d88ba70df36bc3bae17ea299d1d8b03c2b855f0b3fd6ca374565b44ab7e4122a507641f1a6ed61ed9b8128e9bf2fab11fcb34dd0584df5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8971da2a817fb8240e18915894e46e6f8a553af77004705d60539299f232bd52535e704ff899ef3277b4089b620a0a47ec65f8a430306d592b1a98f4f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h707f2c86142655d008a3d29418fbe9ef4d49a2b7b88ceefb8fc3a7772d964df49307a7f0423ec86a942c057c8ac3fb7105f5524dbfd625f29e7e9417e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h64d7384c4b72f9b55c77eccf387ec6417108a5dba086abc6813e94a8cf96894b750f885e4c879232e48bc107d8238de7336c680f1978e9382ceac83a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf75519e5701159a55c0c529cfa97f0ab3c842f7f234f2757f16ffbf162b5aeff0f89becc46ad569530ee1038af7011b1378555192a8e9e7081c6b7120;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h44836e7088aba99e3cca6692c4bc43b605b0adfa87f13a3fc5bb21d8975ff80715692d383207c689980ee7a5dccea8d7b582cd05d6f88cc8385bba53e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h76e8b8e5210887057230c3b07b800016efff499cfd519a4754a928f6cea067d1771267438b0cd86e20b061134baf41272dab55edaba85f40c28c26c7c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed9602d3d1d357c544dd90d75be5d7d7134dcede00f77c4f4c473a3363ab576b2a7dcf2d04b90be3e4f2dc239f2335fe68a93881ee39f431d05e95914;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96d93780348b60551c021f812cc053a1e5d6b20d6ce188d9847cc01e8773df1be21c8509adfda725541dff3a64c8afcdd3ebb494e5385e9b2d5254354;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7bb5ad2b7b96de093ab4562e8e3b9340944fe7e75f6f0f0d6e515ad24b0c42a2f273ba2548e6e1bd4c4c3c07cd416c6476e0ec4126f165bb54c38ecec;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd19bce857c3e5da90e1d0ca8775706511a758fb1236e368484e7ca916e18ce7d9114cfaa14982f919a62fbb819abbc12edd06b62606e6a87c9b40c62d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf345013b31a310fc717a649bdb7b33298fcae24262ff243a83be209300cc5401b70422ba31093fd3653bc248d2598b96e882fe7f3cbe67378d47c9ea1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4d45e05aaf7d05dc2f7ea9f6370d7ade252271043a984a472386f5e7de441cf18763cfe1043c7b7fd44ccda2ad930399f10af9f3aa5ac76e1dbd3a29c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d57da5fdd53bace7cff25cccd82882dbfcc88683953065b40847ec9e504038eb1668c163d3c0540b6d06e806de8a194b99a005f92eee19b43e279de9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43e397fa1c74d3d961db9371534225466df09d4f39a5603c84bae4e3c7b6929869a2fefb20165156ac5bce69cae60532383390e451b489c2a278d9132;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd00e17e2c5c6de0d8efda16c3933463fd73503301cdfb1c84fab61b3b92e69b094b6f4ad8cd3b86123d89e8059d75d6fb9a62e6db6cecfef0318adfda;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h79671b6c7c7f377162c16b900a4f05e0f7d031845a942e1de6330504b51f9a4ca82b12928c6e142e59790e1571c3d0c2a91b40972d547151d5bdcce58;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb4e1f3966ba4233196d05c95461e4a62e6a7e2071d53e19d7473118b4bd1d012e82aec898a7a11a8f0ff169575a1795bfa0e05c022e4dcb00cce81b03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h434fababa99b67922ca61a3804ba3dd059dceb8925f80d743574fce26d94da4d10f5ae9b0ba0dc04d2fd53f90b44f38edd6d753d40f7f60db18c9c459;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77a611c6d591cccb178237382a9a5a0b13d4f370a6f54332cc30007c32b7000e41241934e4856216dc8165d195df2d6b77311bae3d2992627a0863af9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h443ab5132c529fe7193317432843da650cd1c1829f91255768859457c647150e806a20ae53b626fd47b4e974d488253784b9ba293a0dc5d230295a536;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5bf45eb5b47ee9581767767f082a1744c7cea8f573c871bb7b1905d924710be91142e58bfacc2e4666f0d1775f431ad9c55d610620d44208bbc977016;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h377a4df3f9ded504130d6602b789ffceadb844a92bd8002e5d87851b0ef4cb466519eb5891a9fbaaca1b12ba0748bbbf1290db5abc4732ca8f7d9b6e2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb16491abf33d7c5097ce2619376d048fb13d6a2cb3e1897f7fdf48e608dd4cee147fb3c9b2a145aa9fb0e374ca2cadbbe20e3a84503d92ab5ad70dcba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1a48d33ca046bf044fac8a6a0d0d495a800790195c9ede9ef72aaee3d2f6c17fd543faa2bb7893db90c9cac42d68e5e06554018458d06ee42e29d128f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1f9a07859f716c6bc3a375128707eb36442905a5479ce5fc5939d4103c91f397477dc27ecd4be4f4809851f6f58d0ed806b91d28bb0fb52c6d2b82f89;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h83e9333bab6f213e66814036a5a6eb7e6dd0a35337ef645395b1673df269b291ff05ab02759c5a10a3ce10ed12c8c8878131dcc3d5380c7dcae63f76c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2a0944ec9a709dee7e06a2719cce4c07649190182b22f69fd7691cc6f30f38f296ad47a04a619386460230657df3aa33958534bd4bf10f3bb7fa5d9da;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1c4d8696519070150994ee8d65bc26de70b309fa660527857064afd2eed9134072230acb52b7dad99c58ff126eb8efae40d1ae186ac121d95506fa96;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h590b8e848a0a1e44e604a87a44db6a0be314b28e265a5df42daabe172294f772d135a03026d5582e1c721027c982b296c1e9086a16ac91553d88d7371;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26979b8cd52c5037154b18d21c9934619c9cf6dd953bc9084b50a0aba2554153e6e4c23eca40dc0da8d128691c6f0075c5b3bcbdf8c5e7521482b63e7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4e2c9fde5b3a11d66ca734d8997132a8a5a532bc0ff3d01e6be73b88bcd5f3b4482b45f3bd1aa003c62e91c80c0b299bb3edd384c9be259440d0512e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd49db604299ade20e29e6dd5d64e3a67381001c50c1532bf35fdd3edada121915ff71152b9fb3e30809e4b582ea63e35856ee33733dc29169dbbe536a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h15f9a27420b5329ed09097fc587701c1f97db8dfb8b082525b469e236463d4fc3392cc822ff6e6b33e3a662bb5f41fe3deb071caa7dc7191aec76b185;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hac8d6feede8a6efa8ab2ffc1df8820dae4de063ec395f7fb884038cbd7129a0b46d3fc102179a8fc58d1c5fe1e8d101663d678fb40a75cdb910b5bc4d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h66a2faeb1b38c581c3fd47301c89e0b71fef3dd8aa949b0c268d91dd9dd8768195a01c40ee68a045fe5427e481668daa30b4f6bf50f1113d2ff3886e6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab75ea152770d06f7549ef367001d564bfd018355057b71b0dbbbb8d958ad5d1cb2d601b225825cad3fb0bf8387a1673c26090de6c752b9e4c44becb7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7927f2ea086c337b777210b39966f15872defde04f5811ba79737b7af14b380455f44420e8dda27118fbdfede5d548840e34090cd6ca8e9586c74fbb1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfea2fce874f286be8a82a7734a8b8051b18a07584e4b47bb3d8bbe98522741d4da87f28bec7471f94963ed32a626dce4059248787c23634b86039e2cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2042e61b9d546fd2736f15485ce26f0d52933a348f5da9a5c60e2a9ccd36b019cf119ada8b07b840d9c931c37e6ff57c92916e6d78ad3613a0654df09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbba104f59a1f45db28d8d24f3559ab1cd144684bc2a2c8b089af2d5a82368b6a8def801868fafdb9d1939e4f6b4f1fcf862766dbd76ef1ef45337ac53;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5af69ab402c9f488bb070b17a36df35c522cf6b904478b7598a339f85f727907fd79fb00ae85c9db100a022e9d952cadb83ec4bb7bf6a937cbd4cf452;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha5046778e4e8266c3659252380b26fda1d1deea8a8cdf74e56d37d795f8a327db2fd5db29b293b40351f21a90babdecedb1b836f8034838a3a9917735;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7c954e18be9c7b167407f427eb1099cba4e054e10ea8ac165818d854674fca1a6ab9bfc34b2ef58af1eb7a8496befa133614098e3bf8a11b4b262b04b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he4630f009b5190db5eacd2bd72cf65dedea6923d93fcdac0b97ab6295e570ee7692d7d966a5ff0383f68f1f9e1ac1144386944ed755e0beebcc7883f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7caecf16b92af0425935128a56b8ef47e70b141bdf882e73e98e35982f8736d403639ad70c90f609c66f97e953079cd101c788e318dbb30a0cc9d714b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6fb8074c805763ecc81df6819ad059809b92f5b8ade866534cdf0dac8d382c21a4e5e45723313b0738940678221301d6a01e1f7a55ae11f3ef6e8cd41;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf7e7f8e9618ba2e04ae2b28cb17cef451e65b977b3dec862ef6421e5c3d994bfa9e7a64f3d1ba917dcd55584bc3b50aea6a604787d2a1b8c889153f6d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd67183f6cacba47e71a7e341e991f0f849e77166f3020666a6fb27a9e08a0618b21d1ea636c4b7a8194a1455323e1b93bc230f95e2e4ec967536ebf6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'had380c98e792a1f88dfe527b0d247424178b00fb80dfffe089059438a85e297b1d0715294e779ca1910a319615157f3ebdbc1019306fc4c1632b5a18f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h264a105613393791361766b0652e8d2ec8775d8c26142cc2e6b6f8493a22e153f119fe4acfa2d3a73dd475a25975e26733c84340c280dbf8a716f5985;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha0d51ec98a1e0f09ff06c89dc12bea9b923dd7d79c71e213409b1058cce62e38e42656dc5f81652049aadf1217a15518b878f0e3effb3c1b81c35c492;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfc0379164dd19b1be05d763894af962cecba3dee86f2dc109c653f871dad3caf317ea5f9d4c29fa3567f97223ee1e0c04c9fe71bda39b88e78b856469;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4f42dcfba04d920239df606068b786028f555bb7a05b9f6b23d1352f3e21117a7e6191d97059ae90cd04a876c3b2b42fdccd247f793b89683ec72ad33;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7d8078dc271422d4ba6e36b8c1ce47e49161173db32984577c3baf562a667171b721e7b5ff402155e3943018f51222eaa4cbef31ab4c944dd217614aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd50c5a6170f1f4e345c0ce47f95d0f8965a77f50475a99c0b5020fcd36bef9c3a33b4ed60fa0c408800f32e3269dd308a3abadb77780dc37afc590e5d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h95cb093ca460f6fb97681e35ecbaaa7005b01867aaf42d6516eec2b3d995605f6bb95cebe13b8e3a56632c1d4398a5c6f167f7088392dff5ada2399d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h626c56bef8ca609a1c052a2cf17db2c4aa007b56b87a3c78b96a39702212cbae78b4c2d271973b31c3ac02a7fa10ee1158a9f46659d82dfcf0a5e27ac;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8ab3c401ee212014366b34bed909b330a3a1ddfe90cfc489416d3579e7c2370885fe71d707c8c98390cc960d6b7f307b13aaef98a79be8a56137d00b2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8388c211454b9a930a54240180e5011e153c4f049c1c00de70184a23cc849c062d9f66719facd7550c4efeaefbfaa153cd5106b976f7a701d3d1b316b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19b2bb1fff5d3e4ed7f8bded63d655b0ea7f7282db29bcfc03e1a018e2fc23f6a6d9e05d2428091ffa4f10e71093d6bc3ca06b42ce2dafd7977e83998;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha38c2a5e754f0c85fdbe58d3c1179b7bead3468b8282cd833bd62959f13c06dd1c3428c6c413650ac1c0ee8bec7b72dc690ed46b36e358ad0b55761fa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6c1853b41591c312e6caf7bcf8fd2dba4ecafe6f5576943f53c193805ed575a47460b58c587358860a1a58adef0a741392e638afad7a8effe138d0c0a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he9e1d76519b820566f45493ef9c95789b539a0b3a2b8eb0a5fc6d0eb9ae2ebd8c6c4c6f96c5353b5644d9f298519b8c7d861c8f328a0271198619d519;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h696743cc4c36832df42b56c8ccd1d2bc1d3bb483c631d29ed991bffc690b0591cc27e1394c821fecaab7fa3bf1b6fcadbe6f766dedabccf0c9fa36deb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h307dc5f20b6fa2457673d03781e9c89fe2e98eec2a527a28483eabb3e08d4bca491aa91b6872a46461de4cdd676dfe938027fc948a9bf33d67a3a040c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf36b098e062d6bf00a3667b93b10f0a5c6513f5d55f53c75f3a77db3183af5e255c58a485f65af21343039dfa74c03e9c3902acdd601f45513592eb98;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf01ed543b58435a6cbbc8dab98296a651b86ecc3aaa58b5c4a29b87e61a7fbdad1adc6e6633a40accd1ccbcb0b0eee2196bd21242c4d4c5e23eff3d01;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef9ed078f67300ee0da672f99c1ec5cae990dd29763a0d212a6fa9c3258cc46fc8b218d90a287ca159a194f4c2f940744fe5ecb6cdd8a0d5b4085da58;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae7da27591097a3e17c89e05996275b72df310c672f41f62ee304d69b19c50baaa93df414dfbb678ba350a2f264c044fab3e9a725ec24af2c384c4279;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc71d8cd053f745f3441503de8be839e400ee723ea69e17f7eec5713934394727de0683931a9447d23d57858218cab2cb8ef922dd98f02838ddca5eeba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e42019c1bbbb299c8a1767fe7adeb375ee7096adf29254abda5fee6c2ef4fd5110f80efc5215247d99e0da387cd347f470c93f6bf4a67f8f1f90fd6c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7203c49a2c080537df71a6dfdf98c0991d5f04a0719a6d0bf61336155aaaa6165f1e816794f308e22a37bcd23ea6994db0ee94edaecef7e286bf40c00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he77bb6cefe044ae408fa6f3cbc09a096e8d297f072393002c48340b3ed16e194e3003481bb0eda56df61d7bbe0238180c86365824c61d5cf7ab0f238f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6f3ef24a288def7652bad6c842b2b73812012b51352b0882dc8e4b7a93cead383494e12b9640de207c91740a0deb5b2c302048c711a8b081c17913882;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h949d4a83912a49c70ee209a7095ac32d1132bcb2ad75ea3427cf6a550c15e474ae6cad79778de165a71c49c977df1e5501e0a7fac38cf427d338d358b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3195bfd4ab3be2261128e911d75d221a3a1a752a26440799d6988793b666c46221d6793bf6b5697e68f3678c18f848e7ea98a75b7493989ca39a61677;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbeb23902d25885a8ac27f80ccfc60401b0701ef57c8049dc3b02438b42d2005941c983e29cc302c242429eea0221bca0c376790abcbeb9952a831d34f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdadad8b68b95382e8a6d59f028b81ee3f34a83d5dabfbde00ec6a7c4f66d2a6f108ca641bdd6251065bd3f82bf6c325e67a152845ac0d6251d208ba09;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69af9ff0fe64050436f5b71a7475a977483fccae74ac7d483da58e5d9ca16f748b48793457f0a867d44006c6beed17617f7c4b2b58a6fcd9746a5d76e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1bfac5011a4ced33231fd6730189db43dd918025e679ba263700725fba0b3c1835a6fd0db6dd0fbb4536462efe061af1e18340c311132447d5bf0057;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5c0ecb4377f268496fc4861453df1656e8c5ef8a17c78c54ba438599e69b81b0115f99603ab0d3954b6ff8465602a08825f2e7d4f5eefe33f12a66288;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69fcd225ad56796c30db875f11790055c0679a4a900d45841e82bda2c45039b1ba47a5954bdd9139a0959f6da7044474224722621f181df60299391aa;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h73a4c4d033a58000bc64fd2013241fd6df5675a01329e65d860969b734f6dd2ba9e792cc01fe7e52a2c6911e00d62c34b8eb0cbc6d8184167033ea763;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb50d05b16cdce2a0402dff0cada322a14f6f8a64f36ce093bbba33fa85427e60eaa833442a5a4cc7f3a519ccac281006d981d92fc5c6c8b0dcb358aee;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4eb5e46e51e8c49c56c9dff37a0156ae8fa7b16becbbab8a775690f0633a3d6712ba628381cbd00587f1b1ddd767796440fbd02b2bd3bd6c62b03de8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd67be93e9120bc3ce881cb0407ed7fe8161dff0b43ca0519e2d82ab6ff57ffe9d4432a413b9f106779b9fd568f1f64cb822d0f87115109116d83a26b1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7dfe29571b3cfd948fa42855212d8f0c4a8e1acde97f5ac3118ade11aef0c023a2241b6339ba3bd12aa02e3c54bdb7d27f0b9dc425884efdf43f891af;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2d4656a218ce120775caa12d696092108257a633da610c634fdf70508f1d61ddb71d814e85351d105563bbe4bb408584ba592ae0a3e5effcda68f5714;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7b16503249a015c6059c5b5c46671f6670cc0fd79e2c0d0ec2b74e2f2d24c233cd3f110fa7823e7caa21a8b3262a1ef615f72b044164652f66200bdc1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h19f5ca0adbf56d99bfa0d2ffc7d4d57d52f7f6d2bc108922220c595ce2ceac29845f3f2b6eba972fb0de5e00e25ae2cb3a25291c98e1d95e375caaebf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71f3f1757ee5403c0e45c68e3ad89d2830fff7ee51bb01a2bb6d9d2020a9d1c295abab172af95f36e89c9caed4d2d0597f39181f4c8b5179b413d2e2b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf499feb7aa994ee06c1071c626f3a06a0b8ff88b430ced4152cecc192affb7504a3b2ec2dfa279aae59eca8be4a67b533c3c8698d04e834c468483986;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h45e859fca6b69bb800111587866c55d23125f84fc0dfe362f742bb9f32ca070dd4aed797e99ca682ecac729281294d011e4787a51c7acc35025b61225;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h89065463912a68303d81ed38f310ee6a9533e7c3ed1a5d82697bb16ccd3e7959f842fc0d7fb88ee0f714c771abe966bbb2526d35804340a5c9c484d16;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf6c565ca93dc6f7afe585a696e15e5305e0365956ba9c0afd275ba6227a790bce852504add48249551d85143d64cbf0e022eac7bda1dee7604155a501;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h291e917729ec33f22a144084a0007ac4b06f0e5dc5047f07f91e3353bcc3d96a64ea2eef8b285e15845bd4298f351b7e6682fb305eb85450becc45a4d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha829392bc9ab388d775885f2d4090aa3008b90c23d29d4442a686bb2bdd35b5ad8a2b1a99c22e8ed2f4ff060bd5928150b0bbc00d5fcd6f096fba9c4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc1367b07573879d477d9eb4c40327e3491abdcc390d2556d9803ba8375ee9dc782be8c3a3c91af0abca41484f5f55182dba0b8fe6b9b858f99bbc7ed8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h32627873c20584e40652a9c84597e3892053ad1dd6a6f51ac2c232ea7affc255d61f9eff8cccdcb4f6bca0a2e7ba76ff73b405110e2e289b6074068a7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h424f51adc503377047a1a3b6a572fd8108f62df88b18496292614836199a5b04b8cbd5c122470bd0a9122c2176ee8c2d5e8e5d4d7540d7f2ece4ba02e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbb2527d9adedaf951a1e6dce33c6183b51ef7934df0d0471e0904c2d981602312eaf371b20040a8f52908d5a692b22f048fc1fef00ad9dfd5170b611;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab9e53ef6a196e4282735b1f848b04f60689dd3c6eaf2ce890f77d6c25f90bd429cbead552421c15c18c71cb59205463a18633c5da923c33c3ff76d1c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b2e9827503c04b1ee6de795952dc171ee59ab08717008d8476f785c2a69a655e79bf0e50a395cf52c37de6e1a0040c43e75dd0e12bf22c9807089c94;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e857ecd6a8ca0480219cfb62c24ba0b603d1c5bd3ad32a933771aee075ddd770eacc9250d4402f9c14de7ecfa1fca5e9d2a8c06df6f69c90cff11eb4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1d84fa9c85a99bea01982f9f5769ec89ae60fcd53f6aa2d3baf4d036cd3a8489f50b020a7fe0b21bcdca8e42ae1ce76ad6f29c201ba6d66935c091adf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebf998accb6065a90731ea7738c584fc4869fce622214b3dfe23bf8566a5056da6d5aa4e42a631585005bbd75983658c9cfc06acd989fa5bb9483a9c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf949a1ab3fbdbab8c25b3152c9576582ccd75638cc24b8d3dd51b7d8a9fb85b31e30f7c568877dc0fc65fcabcbf5ee3a2bf0103d571affb0823ea823e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf996365296dc7933e899060e63cc32fc1f186f106c8c967f97d130fb3194f1be3896c1df139e07d28d5ea452b42c973fe2798d3aacd8d9e29b50b3f0f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h94678f2749a106d7850a0cb566591cdba03eaf43cb33f5c74dc22f4d1c36eae813bdd7b3ac36f56f9d8cf66d19ccc397e48ce8f74cd3fa468a55ca733;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hba70e216c7bf908fcc6bd60808ba71ffb44336a5a205d1db2268e26271998be6b3e01a24963f0fd79bbba4a204de8985cba73ae418ebf6953a4acb9d0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e7d1a9031d9d0965b2c5dafc2a4b913eb555fdd3e61ef6b61f66e6ab39dede638c52131cb0786c8b9b44846cbb77d7907b2bfd8da23a3967e13ad555;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h167f820f98b71e283349e3466b4a5abe2ecdfa7b41b9f5613d31f2babda7ccba0f16b44c950178ac2922a5856ce250cf441346e7c589ddd74d45b1fb8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hffe3abb8aeb69b4204c220a258a3746e697d6bb514d2d069dec94b4d2a1d255331cfaba3ff4211d9119217b415812d754f0bd474cbfd445adc8b94759;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b1529da068a28f7caf5648a0ee104c92dfb5f45ca30a2f3ab0d00593f9155bb8b41f197cca7817e5d11202ed8dd84751113bb80a88f434d0dd89f1c0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a02977e4f9e7f6871ba3bb163939dcc6fadee88e3ccfcf93c32f9b269daa57460a08ab41ec50397e41120a49bcd1ac0ea8a6b3806ad01574295fa0c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h75aa4df7106ad711cd2a3479bea6d82a31d3ba493189be65f4f8a64ca874a1cb233a4b50a14cf745ca367317ba070e2a49c7316b60eceadef4c1948b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce3bfbe6dc7f2c44976a22d7140dcf671f30fc5b07cde32ea8ae7a263cb99fced2108e23c30ad0087a42503c47c79889db0dc0d1e97945ef75284c16e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3e3a1f39d1ed7861842bb1f1d41332fdca555f780d352857ee729a2d231d4081e676d482db2830d897add2fe2a27177bf1e9eb1b3e54a239caa26990d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd7cf18bd97f4829d6ff3315a82eb46eaf2b77d4f72144a6ccbb0aae2d85bc32ecd1385329cc3e8b64ef5e171dd94400d6a8d9a737f2da65feae82f7f2;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h68801195f342741501e1e9400af916c9dde2f451c181b763ef9b07a545a4a64fe7e1eaebf7665ea7150b8b0a0f1e15ec23aa11456d7daed5df39393f1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h87b490e5422c6903c323b7474662db5a667fb581250c79ff97f9772d6598d40e9ea564943665ba5ffe96d7f946c28624c76dde3f6409741d563c85bf0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h788edc9e860a018804edca0aed558209b77e838328cd5b479b55e65a67f2e90bdc7cd0b3a490a8f3f7a01f55bb01acd931699b466c1943f52486dc87c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h946bc423a9530337e38a3029a449d94db0fa7ee5631c51a80bf74faa37040700cb1f37b7eb34e70414e24321fb2d0438d0e90af528eaf4ffe0322cf6b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb866d487b0b81d669587912bb6cf50dd3b53334f9634afe6d741b565f6a2ac8c6c434d788c387521c5a8bcf5eeef73ad508d766cc1aa7803ce237db97;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7e8b06ad3869751054e1783389997137e820497751c373186b68ab4bc5cafaa711bfe5fdb515b80ce31ec45bfd34680c259a17f0da396156ce208c1fd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfffb9027279e949093e3f05c8a9b4c57df107080cb28f288a1bb5b76802e881234e290407d13b60b1cd31a02293df6ad2ca8a8916f02db81f30e98508;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h26794ce20c04cef6039cbb8654d5a996ae8072e2eb945b1cc0b46bc6df87d92c104b89e0dc4afb53b8c5264ed9b37f2d892f89df5010a45e34db76e39;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2b31062a72a69abf1742295a9a2f0ed68665596ead70235fb124b61c67813dde025670013779e75161236979b91f02d88745fdafeccf1bd7d1da8571f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfd535114523fc7af8b76309ebf34008e2558824a2ba4193b950d68d76e2dfb36ad5757f2fde7330a6b6885a8f64bc209ec98436c6b3ec2efd902cf6d8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52db439c610e3dbc07334064ecad15f16819016e7c11cd09fda9ce8ee72dd26468763e5ac1d126ab7a83952cb149f17e48ab73c9ae6d686cdcc43ba2b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc60911890718e1904a26d3335dea0de1cef7918e4484c66aaed6f2af20cd91953f5db1e59ad2fa40b1df5e8e2dc5ffeabd64116f8e388466e24a70356;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdb904e07bc2e47d69430ab64fcb34e37f08aaa10e85b2ff2e028ec038128c7eb2c4fc65f117ac0194ccb95b757862c2dd9bad085ca38f95e5a9a8af2f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h700972e495b3db4be7ed716cba895f5618c98dbc3e63bc69a59b4531651249666d502d9963ab05843fe209bc2a0c8e94354a09a18472cc64a99b44c65;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfb10dd30af5563f06276f95a0eebf7b5861c527644aefd87c473f57721ea785b2ccf67b8ebbc3f65087ae3f8e5ff3e1074cf33a159457610dd78d527d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9c99265855e5eb33560c3e59947e64ca9d720fbbe8f535d297549f91e703eb3b0db510e19da7f1f923eacd02fbeab5b7574d5b03c529e10c6e105fbd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdee604ecbd7ccc4922a53fbe821a1f01f26e1aa2a6988b6b2adc6ed745a06dcd4efcd9478fe8156e08ac3eef7f91a9f5236c0e925004e865222a39b21;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd23e5919cd4217610913f125c391442cb9e82146f56c13b2a9c66feebb0203a253b1991ce3d6371d170487305341199b8dc3ec8963fa0622d4dd19aa5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb7957609865cfc79fc4814394605ace5ca28e18e76781611fcc83eacf45fd47a600b4e7919d1c2decede407f505d92ec3d3494d9a781a394be3ee1faf;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hebcfdc2359877adaf2d1921bce83eb764dd5ed00835015b6bbd9273a62ce30271a9d9ee10f7b84e009710310e7f75a9bf57fcb94aa867029b219bd62f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c740503b39c9a7550b400ad20471f9b6ac21e44c64e2cab5e3724d67350c66a9b64943f520ca1f03e06e9ab269a812557732f58ec2e3c4c35aaa57f5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h51c55a8b79343862c078778853cee41aed2f2f1b40bc2546bb32e47b731f4318fcc9474f4b06bbf5b6748c23307f5626e57009dfa0de921d3ec9aa3df;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h59d92f9732f6ab1f12f584d027f44878f600d60a1786ca5436a66d80f08481fb915bedc5d19cb90e5a1380231a3612aafffd22b4667d235600088628a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h72dc6bbf9c4eaf9dc555df339cec3e800ef137e7c1e99862324bf7a8cc1f495ebd3ee684bca26a3724dcff46a30176d58d5a5aa3de9065558ee87b70d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h39965005868f2a887b03c980a3f7e6c48fd3420073289647716cd2ecc3cad4c31c9cef720ad7c0d5f14adbfb73c1017d9920bc05b3f94bd6b7b697900;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ba9945a418dcd9e03de90ec7f82bde91ce9466de3948a1d8e15dae527b3ba31bc83afe4b2d2a7508b94cc6fa4915d98b8b69ae53ace895241faa402;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6551b9b7bbca51d23f30d4119c3d7be753ca71eda60fb972ef276cf0315fac7f395ff0447bbe7ad0528a91d78e5bea1a0d4821fe50587980b6ac70ed7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'heb6c935bff82e97156d585ffcf13ebfc5ee4768083ede9985ce7261795ebf5d4b594c06684a37aad190bedaf5965571bb05c920221e850a84578c91b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3eb9dd17daaaaff595c1c1184bc545bfd28014e7757981b272d4c0cf31b0ab9da9e7172d9bfdc62968c2a0047c4101b6b70e2093df66364d9d68b571b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9413bc9cc695ec76a42a8085a5cf5e8f129a4217b0f3a4b547bef94c4a21704706ed62edd2dd2feedfda0a2af67922205fe2cb2367320a8dd13b5de38;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd90eea25da776555bfef3cf35d3688ad65ed0f6977b3eb6871ba32c44ea1f18e4cc387366894f2b46edf0d7886a2ddd12d822ccbfcb4267ca5622c94;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1b3c5b7fe3c8795f408cee3347be137310a4825c8df38934f26ff56ba8dc1f26bcdab2b3a250004baa3b0b54b625f6cfa8df057303bb16a6c141fa5de;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1c9180c27dc10e609faea7819974018c641f34b808affc280eb21792da668ab539e4ac10c3553ca77a696a83e458bf7449b30668d7fa79774f15686f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc18284286ea6feec3bfa64d8c00a228c603c31570e8e8d44d73b3b40a9bc0a933eba0c87aeb4d4306c4278c6c91fa9d50ddb4877f7447790666c88136;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9d506076a5dd3035fedc9c3ba3dc9ea8e26fee98a615a8a59b510c2ca6f1f9a770cc0d164d0da0c0aa6dcb60a078a12a48607ca89a5f093cca41a34d;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70e0f099bdb2fcfed3a0ee95db4d733072fce6c0071c40cd744cad05b6cab60927d38b840c42fb9e53c24269ae18d3bee3c5acd6806d1cd2f8763c806;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31c5c437389456240201ffa9157d1715b67457ca8eda467a24f9b4b5cbc7fb55e4f820ac8c4876ec0ff9d76d02f57e32069bf4211b909725605e0605a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h77c7b78f2852da4d11b8684bb21ea03d7401414477ec8b4165cf23720db91e32791f16c2f28cf86b20339143c81b24c77a86cf733321a58ce57f5f8b8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcd882ae0d8147a21795566391e13870c19421f58aba6336be7d3092aa223d552107b0ee2898a5988a0e429b1457f26bf5b31828e1a042237fe562becc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd6039b1151f58ab64354cfb9382f67c86a2e56d1eeccc9a463653148c89bf493f91d5238b67b86002ab0bddd319e84542378c9ab71ed50b114ce4560f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5e56960993bc15dd491330e12adb18bd13d86c7ea110e22e30f274dfb840841f4617e4f4ea1bb49ab065059c96141553495fc37f439037d108ef4fb90;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hdf19335a983f4ad5065de90545e221c8c774d5462d887451681fc2b19bdd21aa80676b75f36bec604f7b74d88797328abd00e55d51c259140f46b6524;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8c9bd55461f3d8a8104cd88a75fda5628cbead89591af3506a0c15f858bd076bacfbe2b1033ccb9d8ff9671d67b9dfff109851d83e96f47bacc9f6836;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h972516fef4b107279c16ed0124e25583dd3cb77add7b68211deadb7619348500ee8298c6e5d5ca00cc0776e316f89363cde5875115c9f0662902c2578;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3e873b9c8362d2593bec216be625b41677817948f77b99e194db974aedbf6324778d66dd4d476452f9fafc4132f397c936cb5de62aa4dd2f5858f8ba;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h1593aa15837a38117935ab73fb18c89712f0dc58ad7a29a41eed03dbc6a769e767a266a5a8582d12a1a9c1f9324d9e4766d1c3dda9229e1fb234558f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9ff08e76ef89e77f33a50b18c45db93f0898596293a2da360d95d1e8cc4e321b452edfa8d6786e473fd33f2e1068d26d7eb06d579155239ad9769d8a8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3c60af805d99f6ef27213e017459a23a88e113a4a9c71ed0dc17b1ca1d80470ff2cb1050c3b2fc5eedc22c3f81e289090272dc28a804bdf22ef5787a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb66c62b0acf3195a33ba25ff64bb1629789804588bd0473ab6c886b3e3b32080359eac7b00fba88e22f532c8a84ab993dccc42f2aa3d6b4e31f76b1a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb855dbb5751c69db596924f478500252f91ccfd4e38f338885809ec3cba3fc48715518412022a904244179d73ff30df23c4c09dbd57d0d81593923b47;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h202866a5ab4236edb9d33335f2d01089bfa50de305df5f37c80f82a737fa8022904f5cd336fd097fc86bfabf70b31070858d033fee98c2bae35ce1935;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31612b0e9302e98673b09323b3f34768fdc5752c2b495706880da9d691c88878f170085118bd6df888f651c7b5812bcce3fddeefa53c3963f7abbb507;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hed4f7d6ee01b4b9a2300c9db896226d5d36d89534a30e9e28a188e11b029288e0709ff9319c51c484a9a49186499c478b15fa8b74742ac6a94e441709;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7149ddb2f008ce61e32be179d770099c28f5984cc6bb72c76d7d8a96ebd7facdc074a4d340a1e5f4510684a79dfe022842751c415d397ffa328c69e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h3ab32655f21c8f4947746d2caab2e123c97d594f96618802b1348304029abaf829cfcf56c347c42e064846757380955d4b591102195e117e8c487802;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf80f97f25987e8189b6dd3b87d00428385b973ef4dc66f2f8cf057074eb23b20d883c79d8e85a9085db8d50d2f2aaf9ab77584491b0eb01aca0e25ea1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae0bde8a471962fc8d0ff088fabdd89cd339789b3036e6b61f6219757e096078f1e506e5fdd393952dc1256e5819513599e71b82a69457a20c8a18830;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cbf4f250f8203a978a85e4f0198c637a4dc90b902e280f35ad4f1fbc150ad5230daab1860e1f147bebc12a09a004dde9863a3b6d3c77cac888b4771;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4854ba25b47f81f211e5b67df61a51ba671a66f74535b162468ef7ddfe19c32e2332b2127a5049d5659ea254e7c47c20c9d28a58f12c2fa46a4cadeb5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd40e49c8ebfb22958b9af4fd3b7a9fe3da54d0759cdd7d5bf3d823d138a40c4d33849d76d25b89a991f7054ebe76dacc3be0a2985cf606e59a9f7328;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8b5f9b21f11f4032c76d34b3c4ba5d0fc88f7efa4299cc2ae34fdc4d94f206f5be534dfd2109b92d1ba5a6717f9984e49eb473afa9e66a4fa63407593;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc642f5a169e6231db866ef8c6046ec8e7bad5cf019bcc1c5edc9654cd813236884dd37d86a90c3c8b3d13b308376e86f2bd7cb7e27f3ccbbc129b3a1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6b6a2eef878cd03c0ef8d062e4546ab3f7a1fd0157339341785e55adb57e17afbfcb3e2ee310ec683185fdc022b6fd934b9586e96e05f668e63c8834f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hec59d2d99279f016a518ccd92b14034c78a548c979d423151b27997c0efdb5ec63aad170cd13e0c353b702c004649e3356d19d19a160b3af864654244;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h43e1ba7ca0808bd88640927b2c1df7b73aea4957832a70024003b260113d2fb7b88ce48f0dac9329888b4f3068d8ca9b11f8d79adb4bbd7cf327038c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc434bccf2d11fef1a6c0c19093a9aea8f3eb862643553f62b421cc98229ef85103956b3092bcef75848a140f799fe37ee42ff91d9a6b8536047a92016;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he3648d293308434bc293c09ee1211b6309f1924bb45ac37e33c334675a227dd2a6d4ce5ae46ed1bc6fdf35d0587fad0377229d93096e3a3f532035b57;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4027e1c56cd6ab6e3a19f4c4bcaa3616f949b8b4797c8a4a17428120460af25f93ec153621e92f3f3ed57a3789864c83a3d31f40b738cd3daa2cba109;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0da36c704302291f0605b6a11c75b327f99d558b7ac6813358243e8de6e330420f7f20249dd7c25842c1fbe3f37fc54a74923d106817763beb10dd8;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2551fcbb06c0445ef6ce677478699beceece59052959a93968fc51e6cbdd774ce25d2e335136cfbc649ea273c74d0d09803b50a06ff612b70a37fefbe;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h462aa05dc2d8312643b09dda424245d996f1e6d706bd41ca0cdc1b2fd3fe3d8f9e2ee9d53643bc71ca3fe9967a6147a5525f6a71cc0cd90d9fd881b92;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h822d277fa0e87d033901de238ec47360aba82443aad981a9d7b5742ff26ad9667fcf4c0ee17a82b684f5ff811f49ec4b72bf16ef009ab75d69e7e3f00;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h67381663f03988b2227d170c7e0e3581677dd92377a590970e7c5a84d719746dd0ea779005a59accd3f5a4b060555e037e686e08f5e4fc87e21e93322;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5745a77dbb9a883746b25de08ea108e8e61e4c6a660213be9fc26d457e1f057ad9d862457d7caacf1b9598557d95214ce2cf9c3d673b04b240904f640;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hae4f736ff899dec1afb4bf8f18e17920411611f453a1224eed021882ff7177a6a7bc0cf743e778e4d30f1275c627841bb5dcea8132d28806cc1edd596;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35b74a3e88c6d25e855beef6d1d566cec110092db10be03193e4a0de93bf3f4e7cfa9024c0ff31efed098c00fe456dd144f16aa648353a321e89714a3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7892005c12ec98e8d36d004ceb7761802e30f719f8e8099ceff1728c0eb18187298a405757f862ea16243a1a16a666828d95b818937b980e193dda4a0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hda2914cf724243bf28d2cb501be90e5746384b66bb1eab97703aaffe4d2016fcd4809bb90e68170178be4a032c75662bc961006b2ad60576088619bc6;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h279c9ac5b58a9acf4faaaa33c5dc85de7a457c9e9445e52a0ce921e43aace0cfa0d4270a226fbb4b676adfea0e1bfcb6573f6533b08ad837f70bf91f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hab53bab182991b1706a32350b3e1e68939c7ff4e282bfd02f1f91e6b3cad733d15864ecb392e0ee5c7f0b7c6ababefde3f4c60795719e4516734f6fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h52ee11e492bbae4a9bb2fbc266715ed180751d8f5a9a07af8c471e3b303d7fc8029dc60f20f9dd6613b0ff48e32458cdba8cf0573058db9b389bfe5db;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h40454a36e84b5f398cd99d9aed64986163a8aa55442079ba081a8fd35c6fa528a7c68639e53c8460ed3aed9f0602b8c2865fca604e98efa81b5ee1d43;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hade48643674ceb4c96173d296f99b342253e8576b180385b4381de4e45063a0606b711758b730672da90673ccba5c6864c391a8a2eac55e8f17f0862c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he7f0d4f1682dc3c92545fb4f8d9bd7415c1f248b43429fc26df74fc335b308c65f2f79bb80bfd387e91cafce58251d190bf651792b637d557fcba5264;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h681e232c42ea667a140ee4675cb1c766c6ec4e68d17babdbfcb61cab61465f901b0cfc2e4a0cdc4b71e30106a5684f549759e8eab346a52fa6dac42a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h70952e3c4869646bfde21f3604e1ce773808e377ebc288e6af94742cac10ecdc67ad2fbd387be3386fb0b426c51b2805d6411a7a7feb80237b742fde0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4cbd5e53a24f72ea703c4a0a263c96fc54e20cd223af62c45877ddb4ce20a3e4667e49291fc06624678d107db30a40ae415f1fc2c814f4719c2df131e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha55be31d4da4a89f56853a8ae24c0dbe62eccdd63028b1b8c2b2fd479b14b08f76a230c0ac9dc1a23e0f52955d4ed20efba7f9435e66dfefe23b12151;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9a1229790c48e7b33bb0afc7b6d0794279be47e9350eb368f0540ad0f488bbe4d166c6a2f458388862263a1117defffe28b4cc84d4eb474c63f55e5e1;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc0763d1b566ecb7df44a6d3546980a5133b8eaba320e7045887ca4abe45dfcb25b7dc48c33925741b9970814855dd466eaf79c7ca47f09750589b3e2b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbd371688b280580155870a5c4924f8cfa1aabdf88c26f89394cff441b00c6f783ca79c3c5ad5da8ebd3fe318fe75c0e89c978f0981921d8c56586d0cd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h71f6925eeac30eff14cbe3d77ac7538593c06421a0e8e374fe8fc05207275fe3ac8fd3226c1b51ce6b71c8dc1bcbd3dbf47ee5842bf834dd46f9edc4e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbe6cdb81915145c28a6b7a0d3274c0e20d16da86e2669049d2c997652645ce86df4656aa7bf11a6a3d14ccf147b1c4467f798204ca9a39be8731838cb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9bd287003164b49467c4ed4cbbc18c806691de9f528d7490c58ff916c5c7adbeabd42e01a0200a65b970a978280f6baeeca2345bf3a5388bcf9bb633c;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8569f319e77be6cf1e8d9ca7968812a4cb669c7c71ed03ee17e4c6771f0af11b39744dba9eb54e8dc26c51b0685cfb197587f6dade2f52909315febc0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'he0d24d444461ffcabd3759464fa532ab17fa8cb492fe515e7f4034ccc0eca811245bddb8caac61c5b60c1514b57c1107808f7310f543ba7bac1dfae91;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb1d6bfd12e330b24e86119d9bc6013d01948883f8e2e1be260419a97c1447eb2ff057d7add4224787f181debf12ab49eae1ac49e43991aff529cc24e9;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf08f3ce651fdabbb9b085f022a67e3dcbc9aef0c6ca53fff36af88f6719293c367b422f24f3ab302a5454e9a5143f86aa939c47962cfed442c5762ee3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4fc5dcccb0c60dd2c1fa8fcfad1ef8f60b6388f80d5e8e9ee2e75013857cd79a7006f094df4799f7daf942e466e845828b39316d15cda7dfecc91ebe3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h96f46f9104c0e557d934cf5b2ba20f11f2699944fd11865154272ea84adaedc6693f7faa361955efdb2dcb717b99708c17e4be971670781ae2c1796a4;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd514bf330d77b15021729d234e4fbc57aa6301e8735a43630e3e7be3a1c4dce77e28e32dafa837b701e5a810fa455e732719d2378bb5cca4235d1fd0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h950f2c13e2861f16ee44c3de20ec78587c142c0fc2c577885a5ce8fdb92a18366157e2a59158590745d50d7cf5ac70d2d3c5cb6908037897011dbc51a;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h56b22d4624a41f44daa4b2f35261fb57100cb77a68b32fbe786f1fc185adc9dcb637be2f445baaf4c3cd392aa6f6063632a9733db20fe8183b01783f7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h9efe38120ff23f4df61b5bf0aceb88dc0f09e4000e72e7911d6766f7f55b2cb08df443d253d93a60f36fa3b96428cdd052f9b03f7897d22589975a805;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hcbf6f849e8585e10a927a4d8d2e8c75525656050655f0743894f21b66059cf291214ae71113773c9ce3eb6e73b6b9249f94672c2b03422631cc5bcdcd;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hceabaf1228faaa96de0f250704eee7cc43c573bb1aed151655209ad7dba9be5646b8e209e7e1e975aeb7c09468715cc4c1e0cf352c5980b89c8992a2e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h80e7c06084fbca6636ee808f39b954636c87228a36b1565358eee6354523d6b211c7a1cb207072da937d3a4f65b046aca388730c1a481c5e585c507cc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf4db91c5d9b01c357ab3d804a143c7bcb1515bfa20fa739b026e0658613cde7ef410003800210b3e74fdb452cc24645b063cff6c9f1a901caaea8a721;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h6ffe2a7e2f7946074cfdb2e8091be1a89ca0aa63cdb87c351d593b8b5695a921300120d12327dd00f82dfd68eb1d25663c984bbe225cbe70a568e37a5;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hef1fce3c92a633a1cf7486f12ba726a67b65010b99c15f2e0bb1b5ccdef6b1fdb6fab352321898a9cc4f1455bee13858ff4d8f073edc4b512273b813e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hd8ddff2d5fb02298fc2300ec0f308f4b0216d30af689751b96f27ae8874cb8fdde70d7e01ff9aba3ce5a705dc992edbf3d4d290c9fbf307c2a86c2fb;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hbbebcfdc0eb61a629195829715222e10178ce5f81e998360860eea2ec76b818c46fd00709525b2618b563aac4bec3ee920ca38a6b1ec8621ee57a9d63;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h47b0953532ee44ee2c3080911f7d8b9bcb20160aefb2f6577b7e8cc4e665007ff1429f7324adc1b72b2c587d9cae05d25ab58a3ab0ff1cb62bfbcbb35;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h69f4d6c25f6f2b0e3809c6e026ae21a2a8c88e009cff0f39a23015ea8b01c833604b77e85478cbd00f56489b72da9277b8b3c2871c1b20abd136d4265;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h4049457d8737a5023841a216457c68f168a340b18fb065095c6a12155ed761cbe09274bd4a3ef804398017516f2127d7d1b6e2c7d779e77cdb428bfe7;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hc20858c36449e45b4eaf40e28afeecc4ddfad866076c42a2f1b66de804025b1ac940492171fe154a13759856dbb9e752760c23d4b2557b87ef89329c3;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h2aa1b4f82a24356031497ae98994e60ca46c5d15f7ff30308cfad1f8cc9a2710c6204291539f284feb3e5f4009859253471e28e4923ff03dc8d4e231e;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h7a862fd4ba192d48955b2de16c7be4acf44ca83a80c1075245906f555ed8fa14095d8c441f0f27ac3e67c50ad8283e5313a2f51866fcd4399aa1896af;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha943db66b972cbf235256b60fa59f7eed2f2390a1056c91a85f9b33b6caee149738fdba100e14083879d2faf9c3440a763280cf49db5bb3d110209f4b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h31fb152e9ae73ea40e72d9a311cacd1e0dd7b5a9e749626a546c67aee98de7d20834f1085a58002c7963ad67e16e3a85ff72cf216bab99830bf917471;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h35bda7546bdac0dff2dbf0ffb38a254d86c4c93481bf653b2e06fdeeba6421dc7743ec8d37f90ca28975f8ff3e1b4da34504638c9c07c46dff67bff0;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hfa838b20b36f1eeca11e1049ca897915a867a3542c4f32aa04afce4cce3e08f3b795a1e3a09b4e17f7b468a96a724c690a429276442a84622b3c7807b;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h8a423652f0c068a794a70d3ba7896ada08684f90cfa125baf8598331333029d54be03c9592ebf12011d194f579562511fb42cb6f8ac397b042a5546ce;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hce7a94f35cb35ce06b385b05e22915bf9d602e51a84800767bc1664237ea307e9d1a49430e8e84538dfc490a7b324ead931ddcae32612159e1b98f566;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf42148e7a13795e629ba344d36ea4c8b6880f3ee4267fc31829e11fe8aee7ed99e923c448025afa63db2967dcabe601b8ab365dcb14eea826dfd5971f;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h5236c40118fe2bdeaf51b3a3e8e25393c8806e9b5c3179a7dde2dd66400ba3ce5554990b5d1e2ffe9e774f6f4e99a88292960c3e7cecdbd8b8c223dcc;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf9543a3c8cfd243395365ac533bfe3165422134fc10e106fb209e38b3e2bacce712ca0d5341f77dc395ee0e8945fcf49ccdd4753b50d9b17940901161;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'h17cb8d1b9830ac851ad6a764cbdb1e29247e453332f48af7a53008f5540abb12cf9639c6a84758e2f8be4db9af40e826f86c779bf3931cc751e1adb87;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'ha021f9d004346130d226afac59b0cd1e7b0512d335715f56235bca55f1252e5a9a1570bb7e52be72ec3e827ae036e1f1f2cc73a7237a355a0fe89af32;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hf41a0465e15c1c564c8a527aff859b64e7037930d9975d9907986a5069ca5a1693fa63e2799fd9ca1072f1a317bfbcfa7666e86b48e5245b9d7f7bf03;
        #1
        {src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 484'hb973b30d8ad6577086590bd3950d6317d3dc49e41b3159e3f356cadd89096f78372a553dbbd78b772f30f754a3a0c7555765d88c5147df2b109ef6f61;
        #1
        $finish();
    end
endmodule
